module x_100_mod_47_(
    input [100:1] X,
    output [6:1] R
    );


assign R = X % 47;

endmodule
