module x_100_mod_53_(
    input [100:1] X,
    output [6:1] R
    );


assign R = X % 53;

endmodule
