// Benchmark "mult_3_8" written by ABC on Fri Dec 09 22:21:29 2022

module mult_3_8 ( 
    x0, x1, x2,
    z0, z1, z2, z3, z4, z5  );
  input  x0, x1, x2;
  output z0, z1, z2, z3, z4, z5;
  assign z3 = 1'b0;
  assign z0 = x0;
  assign z1 = x1;
  assign z2 = x2;
  assign z4 = 1'b0;
  assign z5 = 1'b0;
endmodule


