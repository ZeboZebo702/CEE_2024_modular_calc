// Benchmark "X_68" written by ABC on Mon Jun 05 07:05:00 2023

module X_68 ( 
    x0, x1, x2, x3, x4, x5,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10  );
  input  x0, x1, x2, x3, x4, x5;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10;
  assign z00 = 1'b0;
  assign z01 = 1'b0;
  assign z02 = 1'b0;
  assign z03 = 1'b0;
  assign z04 = 1'b0;
  assign z05 = x0;
  assign z06 = x1;
  assign z07 = x2;
  assign z08 = x3;
  assign z09 = x4;
  assign z10 = x5;
endmodule


