// Benchmark "X_10" written by ABC on Fri May 26 04:01:40 2023

module X_35 ( 
    x0, x1, x2, x3, x4, x5,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11  );
  input  x0, x1, x2, x3, x4, x5;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11;
  assign z00 = 1'b0;
  assign z01 = 1'b0;
  assign z02 = x0;
  assign z03 = x1;
  assign z04 = x2;
  assign z05 = x3;
  assign z06 = x4;
  assign z07 = x5;
  assign z08 = 1'b0;
  assign z09 = 1'b0;
  assign z10 = 1'b0;
  assign z11 = 1'b0;
endmodule


