// Benchmark "64_64_mod" written by ABC on Thu Dec 01 02:02:21 2022

module const_64_64_mod ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z000, z001, z002, z003, z004, z005, z006, z007, z008, z009, z010, z011,
    z012, z013, z014, z015, z016, z017, z018, z019, z020, z021, z022, z023,
    z024, z025, z026, z027, z028, z029, z030, z031, z032, z033, z034, z035,
    z036, z037, z038, z039, z040, z041, z042, z043, z044, z045, z046, z047,
    z048, z049, z050, z051, z052, z053, z054, z055, z056, z057, z058, z059,
    z060, z061, z062, z063, z064, z065, z066, z067, z068, z069, z070, z071,
    z072, z073, z074, z075, z076, z077, z078, z079, z080, z081, z082, z083,
    z084, z085, z086, z087, z088, z089, z090, z091, z092, z093, z094, z095,
    z096, z097, z098, z099, z100, z101, z102, z103, z104, z105, z106, z107,
    z108, z109, z110, z111, z112, z113, z114, z115, z116, z117, z118, z119,
    z120, z121, z122, z123, z124, z125, z126, z127, z128  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z000, z001, z002, z003, z004, z005, z006, z007, z008, z009, z010,
    z011, z012, z013, z014, z015, z016, z017, z018, z019, z020, z021, z022,
    z023, z024, z025, z026, z027, z028, z029, z030, z031, z032, z033, z034,
    z035, z036, z037, z038, z039, z040, z041, z042, z043, z044, z045, z046,
    z047, z048, z049, z050, z051, z052, z053, z054, z055, z056, z057, z058,
    z059, z060, z061, z062, z063, z064, z065, z066, z067, z068, z069, z070,
    z071, z072, z073, z074, z075, z076, z077, z078, z079, z080, z081, z082,
    z083, z084, z085, z086, z087, z088, z089, z090, z091, z092, z093, z094,
    z095, z096, z097, z098, z099, z100, z101, z102, z103, z104, z105, z106,
    z107, z108, z109, z110, z111, z112, z113, z114, z115, z116, z117, z118,
    z119, z120, z121, z122, z123, z124, z125, z126, z127, z128;
  wire n139, n140, n141, n142, n144, n145, n146, n147, n148, n149, n150,
    n151, n152, n153, n154, n155, n157, n158, n159, n160, n161, n162, n164,
    n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n176, n177,
    n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
    n190, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
    n203, n204, n205, n207, n208, n209, n210, n211, n212, n213, n214, n215,
    n216, n217, n218, n220, n221, n222, n223, n224, n225, n226, n228, n229,
    n230, n231, n232, n233, n234, n235, n236, n237, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n281,
    n282, n283, n284, n285, n286, n287, n288, n290, n291, n292, n293, n294,
    n295, n296, n297, n298, n299, n300, n302, n303, n304, n305, n306, n307,
    n308, n309, n310, n311, n313, n314, n315, n316, n317, n318, n319, n320,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n332, n333, n334,
    n335, n336, n337, n339, n340, n341, n342, n343, n344, n346, n347, n348,
    n350, n351, n352, n353, n354, n355, n356, n357, n358, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n375,
    n376, n377, n378, n379, n380, n381, n382, n383, n384, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395, n396, n397, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n411, n412, n413, n414,
    n415, n416, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
    n428, n429, n430, n431, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n448, n449, n451, n452, n453,
    n454, n455, n456, n458, n459, n460, n461, n462, n463, n464, n466, n467,
    n468, n469, n470, n471, n472, n473, n474, n475, n476, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n488, n489, n490, n491, n492, n493,
    n495, n496, n497, n498, n499, n500, n501, n502, n504, n505, n506, n507,
    n508, n509, n510, n511, n513, n514, n515, n516, n517, n518, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n534,
    n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n550, n551, n552, n553, n554, n555, n556, n557, n559, n560,
    n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n572, n573,
    n574, n575, n576, n577, n578, n579, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593, n594, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n620, n621, n622, n623, n624, n625,
    n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n638, n639,
    n640, n641, n642, n643, n645, n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n671, n672, n673, n674, n675, n676, n677, n679,
    n680, n681, n682, n683, n685, n686, n687, n688, n689, n690, n691, n692,
    n693, n695, n696, n697, n698, n699, n700, n702, n703, n704, n705, n706,
    n707, n708, n709, n710, n712, n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n740, n741, n742, n743, n744, n745,
    n747, n748, n749, n750, n751, n752, n753, n754, n756, n757, n758, n759,
    n760, n761, n762, n763, n764, n766, n767, n768, n769, n770, n771, n772,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n784, n785, n786,
    n787, n788, n790, n791, n792, n794, n795, n796, n798, n799, n800, n801,
    n803, n804, n805, n806, n807, n809, n810, n811, n812, n813, n814, n815,
    n816, n817, n819, n820, n821, n822, n823, n824, n825, n826, n827, n829,
    n830, n831, n832, n833, n834, n835, n836, n837, n839, n840, n841, n842,
    n843, n844, n845, n846, n847, n849, n850, n851, n852, n853, n854, n855,
    n856, n858, n859, n860, n861, n862, n863, n864, n866, n867, n868, n869,
    n870, n871, n872, n873, n875, n876, n877, n878, n879, n880, n882, n883,
    n884, n885, n886, n888, n889, n890, n891, n892, n893, n894, n896, n897,
    n898, n899, n900, n901, n902, n903, n905, n906, n907, n908, n909, n910,
    n911, n912, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
    n925, n926, n927, n928, n929, n930, n931, n933, n934, n935, n936, n937,
    n938, n939, n940, n942, n943, n944, n945, n946, n947, n948, n949, n951,
    n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
    n965, n966, n967, n968, n969, n970, n971, n972, n973, n975, n976, n977,
    n978, n979, n980, n981, n983, n984, n985, n986, n987, n988, n990, n991,
    n992, n993, n994, n995, n996, n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
    n1015, n1016, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1029, n1030, n1031, n1032, n1033, n1034, n1036, n1037,
    n1038, n1039, n1040, n1041, n1043, n1044, n1045, n1046, n1048, n1049,
    n1050, n1051, n1053, n1054, n1055, n1056, n1057, n1058, n1060, n1061,
    n1062, n1063, n1064, n1065, n1066, n1067, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1126, n1127,
    n1128, n1129, n1130, n1131, n1132, n1133, n1135, n1136, n1137, n1138,
    n1139, n1140, n1141, n1142, n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1172,
    n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1181, n1182, n1183,
    n1184, n1185, n1186, n1187, n1188, n1190, n1191, n1192, n1193, n1194,
    n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1204, n1205, n1206,
    n1207, n1208, n1209, n1211, n1212, n1213, n1214, n1215, n1216, n1218,
    n1219, n1220, n1221, n1222, n1223, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1235, n1236, n1237, n1238, n1239, n1240,
    n1241, n1243, n1244, n1245, n1246, n1247, n1249, n1250, n1251, n1252,
    n1253, n1254, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1286,
    n1287, n1288, n1289, n1290;
  assign z121 = 1'b0;
  assign z000 = n139 & n140 & n141 & n142;
  assign n139 = ~x4 & x5;
  assign n140 = ~x6 & ~x7;
  assign n141 = ~x0 & ~x1;
  assign n142 = x2 & x3;
  assign z001 = n144 | n148 | n150 | ~n151 | (~x0 & ~n149);
  assign n144 = ~x1 & ((~x3 & ~n145) | (~n146 & n147));
  assign n145 = x0 ? ((x2 | ~x4 | x5 | ~x6 | ~x7) & (~x2 | x4 | ~x5 | x6 | x7)) : (x5 | ((x2 | x6 | (~x4 ^ x7)) & (~x6 | ~x7 | ~x2 | x4)));
  assign n146 = (~x2 | ~x5 | x6 | (~x4 ^ x7)) & (x2 | ~x4 | x5 | ~x6 | x7);
  assign n147 = ~x0 & x3;
  assign n148 = ~x1 & (x5 ? (x0 ? (~x2 & x4) : (~x4 & (~x2 | ~x3))) : (x0 ? (~x4 & (x2 ^ x3)) : (x2 & x4)));
  assign n149 = (~x6 | (x1 ? ((x2 | x3 | x4 | ~x5) & (~x4 | x5 | ~x2 | ~x3)) : (x4 | (x2 ? (~x3 | ~x5) : x5)))) & (x2 | ~x4 | x6 | (x1 ? (x3 | ~x5) : (~x3 | x5)));
  assign n150 = ~x0 & x1 & x4 & (x5 ? (x2 | x3) : (~x2 | ~x3));
  assign n151 = x4 | (x3 ? (~n152 | n155) : (~n153 | ~n154));
  assign n152 = ~x0 & x1;
  assign n153 = ~x2 & x0 & ~x1;
  assign n154 = ~x5 & ~x6;
  assign n155 = (x6 | x7 | ~x2 | x5) & (x2 | ~x5 | ~x6 | ~x7);
  assign z002 = ~n159 | (~x1 & (x6 ? ~n157 : ~n158));
  assign n157 = (x4 | ((x3 | ((~x0 | (x2 ? ~x5 : (x5 | x7))) & (x0 | ~x2 | x5 | ~x7))) & (x0 | x2 | ~x3 | x5 | x7))) & (x0 | x2 | ~x3 | ~x4 | ~x5 | x7);
  assign n158 = (x0 | ~x4 | ((x2 | x3 | ~x5 | ~x7) & (x5 | x7 | ~x2 | ~x3))) & (x4 | ~x5 | ~x7 | ~x0 | ~x2 | x3);
  assign n159 = (x1 | n161) & (~n152 | (n160 & n162));
  assign n160 = (~x7 | ((~x3 | ((~x2 | x6 | (x4 ^ x5)) & (~x5 | ~x6 | x2 | x4))) & (x2 | x3 | ~x4 | x5 | x6))) & (~x5 | x6 | x7 | ~x2 | x3 | ~x4);
  assign n161 = (x2 | (x5 ? ((~x3 | (~x0 & x6)) & (~x0 | (x6 & x7))) : ((x0 | ((~x6 | ~x7) & (x3 | (~x6 & ~x7)))) & (x3 | ~x6 | ~x7)))) & (x3 | x6 | x7 | (x0 ? (~x2 | x5) : ~x5)) & (x0 | ~x2 | ~x5 | (~x6 & ~x7));
  assign n162 = (x2 | (x3 ? (x5 | x6) : (~x5 | ~x6))) & (x7 | (x3 ? ((x5 | ~x6) & (~x2 | ~x5 | x6)) : (x5 | x6))) & (~x2 | x5 | (x3 & ~x6));
  assign z003 = ~n169 | ~n170 | (~x2 & ~n166) | (~n164 & ~n165);
  assign n164 = ~x6 ^ x7;
  assign n165 = x0 ? (x1 | ((~x2 | x3 | (x4 & x5)) & (~x4 | ~x5 | x2 | ~x3))) : (x2 ? ((~x1 | (~x3 ^ x4)) & (~x3 | (x4 ? x1 : ~x5))) : (x3 | ((x4 | x5) & (x1 | (x4 & x5)))));
  assign n166 = (x0 | ((~x4 | n168) & (~x1 | ~x5 | n167))) & (~x0 | x1 | x5 | n167);
  assign n167 = (x3 | x4 | ~x6 | x7) & (~x3 | ~x4 | x6 | ~x7);
  assign n168 = (x1 | ~x5 | (x3 ? (x6 | x7) : ~x6)) & (~x1 | ~x3 | x5 | ~x6 | ~x7);
  assign n169 = (x2 | (((x3 ? (x6 | x7) : (~x6 | ~x7)) | (~x0 ^ x1)) & (x0 | x1 | ~x3 | ~x6 | ~x7))) & (x0 | x1 | ~x2 | x3 | x6 | x7);
  assign n170 = (~n171 | (n174 & (x5 | n172))) & (x2 | n173);
  assign n171 = ~x0 & x2;
  assign n172 = (x1 | x4 | (x3 ? x6 : (~x6 | ~x7))) & (~x1 | x3 | ~x4 | x6 | x7);
  assign n173 = ((x3 ? (x4 | ~x7) : (~x4 | x7)) | (x0 ? (x1 | x6) : (~x1 | ~x6))) & (x0 | x1 | ~x3 | x4 | ~x6 | x7);
  assign n174 = (~x1 | (x3 ? (~x4 | ~x6) : (x4 | x6))) & (x1 | x3 | ~x4 | x6 | ~x7);
  assign z004 = n181 | n183 | ~n185 | (~x0 & (~n176 | ~n180));
  assign n176 = (x3 | n178) & (~x3 | ~x4 | x5 | ~n177 | n179);
  assign n177 = ~x1 & ~x2;
  assign n178 = (~x5 | ((x1 | ((~x2 | x4 | x6 | ~x7) & (x2 | ~x4 | ~x6 | x7))) & (~x1 | x2 | ~x4 | ~x6 | ~x7))) & (~x1 | x5 | x6 | (x2 ? (~x4 | x7) : (x4 | ~x7)));
  assign n179 = x6 ^ x7;
  assign n180 = x7 ? ((~x1 | ((~x3 | x4 | x5) & (~x2 | (x3 ? x4 : (~x4 | x5))))) & (x1 | x3 | x4 | x5)) : (x1 ? (x2 ? (x3 ? ~x4 : (x4 | ~x5)) : (~x4 | ~x5)) : ((~x2 | x3 | ~x4) & (x4 | ~x5 | x2 | ~x3)));
  assign n181 = ~n182 & ((~x1 & ((x0 & ((~x3 & x7) | (~x2 & x3 & ~x7))) | (x7 & ((~x2 & ~x3) | (~x0 & x2 & x3))))) | (~x0 & x1 & ~x2 & (~x3 ^ x7)));
  assign n182 = ~x4 ^ x5;
  assign n183 = n184 & ((~x3 & ~x4 & x5 & ~x6 & ~x7) | (x3 & ((x4 & x5 & (~x6 ^ x7)) | (~x4 & ~x5 & x6 & ~x7))));
  assign n184 = ~x2 & x0 & ~x1;
  assign n185 = (n188 | n189) & (~n186 | ~n187 | ~n190);
  assign n186 = ~x3 & ~x4;
  assign n187 = ~x5 & x7;
  assign n188 = x4 ? (~x5 | ~x7) : (x5 | x7);
  assign n189 = (x2 | x3 | ~x0 | x1) & (x0 | (x1 ? (~x2 | x3) : ~x3));
  assign n190 = x2 & x0 & ~x1;
  assign z005 = n197 | ~n199 | ~n203 | (~x1 & (n192 | ~n194));
  assign n192 = ~x2 & ~n193;
  assign n193 = x0 ? (x5 | ((x3 | ~x4 | ~x6 | ~x7) & (~x3 | x4 | x6 | x7))) : (x3 | ~x5 | x6 | (~x4 ^ x7));
  assign n194 = (~x0 | (x2 ? (x3 | ~n196) : (x6 | n195))) & (x0 | ~x2 | ~x6 | n195);
  assign n195 = (x3 | x4 | ~x5 | x7) & (~x3 | ~x4 | x5 | ~x7);
  assign n196 = ~x7 & x4 & x5 & ~x6;
  assign n197 = ~n198 & ((~x0 & (x1 ? (x2 ? (x3 & ~x4) : (~x3 & x4)) : (~x4 & (x2 ^ x3)))) | (x0 & ~x1 & ~x2 & x3 & x4));
  assign n198 = ~x5 ^ x6;
  assign n199 = ~n201 & (~n190 | ~n202) & (~n152 | n200);
  assign n200 = (x2 | x3 | ~x4 | ~x5 | ~x6 | x7) & ((x3 ? (~x5 | ~x7) : (x5 | x7)) | (x2 ? (~x4 | x6) : (x4 | ~x6)));
  assign n201 = x0 & ~x1 & ~x3 & (x2 ? (x4 & ~x5) : (~x4 ^ x5));
  assign n202 = x6 & x5 & ~x3 & ~x4;
  assign n203 = x0 | (n204 & n205);
  assign n204 = x1 ? ((x4 | ~x5 | ~x2 | x3) & (x2 | ~x3 | ~x4 | x5)) : ((~x2 | ~x3 | (x4 ^ x5)) & (x2 | x3 | ~x4 | x5));
  assign n205 = (x3 | ((x1 | ~x2 | ~x4 | ~x5 | ~x6) & (x5 | x6 | ~x1 | x2))) & (~x3 | ((~x1 | ~x2 | ((~x5 | ~x6) & (x4 | x5 | x6))) & (x1 | x2 | ~x4 | x5 | x6))) & (x1 | x2 | x4 | ~x5 | ~x6);
  assign z006 = n208 | ~n213 | (n207 & ~n211) | (~x3 & ~n212);
  assign n207 = x0 & ~x1;
  assign n208 = ~x0 & (x5 ? ~n209 : ~n210);
  assign n209 = (x7 | ((x3 | ((x1 | (x2 ? (x4 | ~x6) : x6)) & (~x4 | ~x6 | ~x1 | x2))) & (~x1 | ~x3 | (x2 ? (~x4 | x6) : (x4 | ~x6))))) & (x4 | ~x6 | ~x7 | x1 | ~x2 | ~x3);
  assign n210 = (x2 | ((~x7 | (~x3 ^ x4) | (~x1 ^ ~x6)) & (x4 | ~x6 | x7 | ~x1 | x3))) & (x4 | ~x6 | ~x7 | x1 | ~x2 | x3);
  assign n211 = (x3 | ((x7 | ((x2 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (~x5 | x6 | ~x2 | ~x4))) & (x2 | x5 | x6 | ~x7))) & (x5 | x6 | x7 | x2 | ~x3 | ~x4);
  assign n212 = (x1 | ((~x6 | ((~x0 | ((x4 | x5) & (x2 | ~x4 | ~x5))) & (x5 | (x4 ? (x0 & ~x2) : x2)))) & (~x2 | ~x5 | x6 | (x0 & x4)))) & (x0 | ((x4 | x5 | ((~x2 | x6) & (~x1 | (~x2 & x6)))) & (~x1 | ~x2 | ~x4 | ~x5 | ~x6)));
  assign n213 = (n217 | n218) & (n215 | n216) & (~n147 | n214);
  assign n214 = (x2 | ((x1 | ~x5 | ~x6) & (~x4 | x5 | x6))) & (~x1 | (x4 ? (x5 | ~x6) : (~x5 | (~x2 & x6))));
  assign n215 = ~x4 ^ x6;
  assign n216 = (~x0 | x1 | x2 | ~x3 | ~x5) & (x0 | ((x3 | ~x5 | ~x1 | x2) & (x1 | ~x2 | ~x3 | x5)));
  assign n217 = x5 ^ x7;
  assign n218 = (x0 | ~x2 | ~x4 | (x1 ? (x3 | x6) : (~x3 | ~x6))) & (~x3 | x4 | x6 | ~x0 | x1 | x2);
  assign z007 = ~n222 | (~x0 & (x5 ? ~n220 : ~n221));
  assign n220 = x2 ? (x7 | ((x1 | ~x6 | (~x3 & x4)) & (x3 | ~x4 | (~x1 & x6)))) : ((~x7 | ((~x1 | (x3 ? ~x6 : (~x4 | x6))) & (x3 | x4 | ~x6) & (x1 | (x3 ? (~x4 | x6) : ~x6)))) & (x4 | x6 | x7 | x1 | ~x3));
  assign n221 = (x1 | ((~x4 | ((x2 | ~x7 | (~x3 ^ x6)) & (~x2 | ~x3 | ~x6 | x7))) & (~x2 | x6 | x7 | (x3 & x4)))) & (~x1 | x2 | ~x3 | ~x4 | ~x6 | ~x7);
  assign n222 = (~x3 | (x5 ? n223 : n224)) & (n225 | ~n226) & (x3 | (x5 ? n224 : n223));
  assign n223 = (x2 | ((x1 | ((~x4 | x6 | x7) & (~x0 | ((x4 | ~x6 | ~x7) & (x6 | x7))))) & (x0 | ((x4 | x6 | ~x7) & (~x1 | ~x6 | x7))))) & (x0 | ((~x1 | ((x4 | ~x6 | x7) & (~x2 | ((~x6 | ~x7) & (~x4 | x6 | x7))))) & (x1 | ~x2 | x6 | ~x7)));
  assign n224 = (x0 | ((~x7 | (x1 ? (x2 ? ~x6 : (x4 | x6)) : (~x2 | x6))) & (~x1 | ~x6 | x7 | (x2 & x4)))) & (x1 | x2 | ((x6 | x7) & (~x0 | ~x6 | ~x7)));
  assign n225 = (~x2 | x3 | (x4 & x5 & x7)) & (~x5 | ~x7 | x2 | ~x4);
  assign n226 = ~x6 & x0 & ~x1;
  assign z008 = n232 | ~n234 | (~x2 & (n229 | (~x3 & ~n228)));
  assign n228 = (~x4 | ((~x7 | ((~x0 | x1 | (~x5 ^ x6)) & (x0 | ~x1 | x5 | x6))) & (x0 | ~x1 | x5 | ~x6 | x7))) & (x0 | x4 | ~x5 | (x1 ? (x6 ^ x7) : (~x6 | x7)));
  assign n229 = n231 & (x1 ? (x5 & n230) : (~x5 & ~n179));
  assign n230 = x6 & x7;
  assign n231 = ~x4 & ~x0 & x3;
  assign n232 = n233 & ((~x1 & (x2 ? ((x5 & ~x7) | (x3 & ~x5 & x7)) : (x7 & (~x3 ^ x5)))) | (x1 & ~x2 & ~x3 & ~x5 & ~x7));
  assign n233 = ~x0 & ~x4;
  assign n234 = n237 & (~n171 | n235) & (~x4 | n236);
  assign n235 = (x3 | ((x1 | x4 | ~x7 | (x5 ^ x6)) & (~x5 | x6 | x7 | ~x1 | ~x4))) & (~x1 | ~x3 | ~x4 | x5 | (~x6 ^ x7));
  assign n236 = x5 ? ((x0 | ~x1 | (x2 ? (~x3 ^ x7) : (x3 | x7))) & (~x0 | x1 | x2 | ~x3 | ~x7)) : ((~x0 | x1 | (x2 ? (x3 | ~x7) : x7)) & (x0 | ~x1 | ~x2 | x3 | x7));
  assign n237 = (x1 | (x0 ? (x4 | (x2 ? (x3 | ~x7) : x7)) : (~x4 | (x2 ? (~x3 ^ x7) : (x3 | x7))))) & (x0 | ((~x4 | ~x7 | x2 | ~x3) & (~x1 | x4 | (x2 ? ~x7 : (~x3 | x7)))));
  assign z009 = n239 | n243 | n244 | ~n249 | (~x0 & ~n242);
  assign n239 = ~x1 & ((~x3 & ~n240) | (~x0 & n142 & n241));
  assign n240 = (~x5 | x7 | (x0 ? (~x4 | (~x2 ^ x6)) : (x4 | (~x2 ^ ~x6)))) & (x0 | x2 | x4 | x5 | x6 | ~x7);
  assign n241 = x7 & ~x6 & x4 & ~x5;
  assign n242 = (~x4 | ((~x1 | ((~x5 | ~x6 | ~x2 | ~x3) & (x2 | x3 | x5 | x6))) & (x1 | ~x2 | ~x3 | x5 | ~x6))) & (x1 | x4 | ((x2 | ~x6 | (x3 ^ x5)) & (~x2 | x3 | ~x5 | x6)));
  assign n243 = x4 & ((~x0 & ((x1 & (x2 ? (~x3 & ~x5) : (x3 & x5))) | (~x1 & x2 & x3 & x5))) | (x0 & ~x1 & ~x3 & ~x5));
  assign n244 = x4 & n152 & ((n246 & n248) | (n245 & n247));
  assign n245 = x7 & ~x5 & x6;
  assign n246 = ~x7 & x5 & ~x6;
  assign n247 = ~x2 & x3;
  assign n248 = x2 & ~x3;
  assign n249 = n251 & (~n153 | ~n253) & (~n250 | ~n252);
  assign n250 = x2 & ~x0 & ~x1;
  assign n251 = (~x0 | x1 | x3 | x4) & (x0 | ((~x1 | x3 | x4) & (x1 | x2 | ~x3 | ~x4)));
  assign n252 = ~x5 & ~x3 & ~x4;
  assign n253 = ~x6 & x5 & ~x3 & x4;
  assign z010 = n255 | ~n259 | ~n263 | (~x1 & ~n258);
  assign n255 = ~x0 & (x2 ? ~n256 : ~n257);
  assign n256 = (~x3 | ((x1 | ~x6 | (x4 ? (~x5 | ~x7) : (x5 | x7))) & (~x1 | ~x4 | x5 | x6 | ~x7))) & (x3 | x4 | ~x5 | ~x6 | x7);
  assign n257 = (~x4 | ((x1 | ~x7 | (x3 ? (~x5 | x6) : (x5 | ~x6))) & (~x1 | ~x3 | x5 | ~x6 | x7))) & (x1 | x3 | x4 | x6 | (~x5 ^ x7));
  assign n258 = (~x5 | ((x0 | ((~x2 | x3 | (x4 ^ x6)) & (x2 | ~x3 | x4 | x6))) & (x2 | ((~x3 | ~x4 | ~x6) & (~x0 | x3 | x4 | x6))))) & (x0 | x4 | x5 | (x2 ? (~x3 | x6) : (x3 | ~x6)));
  assign n259 = (~x6 | ((x7 | ~n260 | ~n261) & (x4 | ~x7 | n262))) & (~x4 | x6 | x7 | n262);
  assign n260 = x4 & x5;
  assign n261 = ~x3 & ~x2 & x0 & ~x1;
  assign n262 = x0 ? (x1 | ~x5 | (x2 & x3)) : ((~x2 | ~x3 | x5) & (~x1 | (~x2 & x5)));
  assign n263 = n266 & ~n267 & ((~x4 & ~n264) | n268 | (x4 & ~n265));
  assign n264 = x6 & ~x7;
  assign n265 = ~x6 & x7;
  assign n266 = (x1 | ((x5 | (x0 ? (~x4 | (x2 & x3)) : (x4 | (~x2 ^ x3)))) & (x0 | ~x5 | (x2 ? (~x3 | x4) : (x3 | ~x4))))) & (x0 | ~x1 | x2 | x4 | ~x5);
  assign n267 = ~x0 & x1 & ((x2 & (x4 ? (~x5 & x6) : (x5 & ~x6))) | (~x5 & ~x6 & ~x2 & ~x4));
  assign n268 = (x2 | (x0 ? (x1 | ~x5) : (~x1 | x5))) & (x0 | ~x1 | ((x3 | x5) & (~x2 | ~x3 | ~x5)));
  assign z011 = ~n276 | (~x1 & (~n270 | ~n275));
  assign n270 = ~n274 & (x0 | n273) & (~x0 | ~n271 | ~n272 | ~n265);
  assign n271 = ~x4 & ~x5;
  assign n272 = ~x2 & ~x3;
  assign n273 = x2 ? (~x4 | ((~x3 | x7 | (x5 ^ x6)) & (~x6 | ~x7 | x3 | x5))) : ((x3 | (x4 ? (~x6 | (x5 ^ x7)) : (x6 | (~x5 ^ x7)))) & (~x5 | x6 | x7 | ~x3 | ~x4));
  assign n274 = (x3 ? (~x6 & x7) : (x6 & ~x7)) & (x0 ? (~x2 & x4) : (x2 & ~x4));
  assign n275 = x6 ? (x2 ? ((x0 | ~x3 | x4) & (~x4 | x5 | ~x0 | x3)) : ((x5 | (x3 ^ x4)) & (~x0 | (x4 ? ~x3 : x5)))) : (x4 ? ((x0 | ~x2 | ~x5) & (x2 | x3 | (~x0 & x5))) : ((~x2 ^ x3) | (x0 & ~x5)));
  assign n276 = (n215 | n279) & (~n152 | (n277 & n278));
  assign n277 = ((~x4 ^ x5) | ((~x2 | x3 | x6 | ~x7) & (x2 | ~x3 | ~x6 | x7))) & (~x2 | ((~x3 | x5 | ~x6 | (~x4 ^ ~x7)) & (x3 | ~x4 | ~x5 | x6 | x7)));
  assign n278 = (x5 | (x2 ? ((x4 | x6) & (x3 | ~x4 | ~x6)) : ((~x4 | x6) & (x3 | x4 | ~x6)))) & (~x2 | ((x4 | ~x5 | ~x6) & (~x3 | ~x4 | x6))) & (x2 | ~x5 | (x4 ^ x6));
  assign n279 = (x0 | x2 | ~x7 | (x1 ? (x3 | ~x5) : (~x3 | x5))) & (~x0 | x1 | ~x2 | x3 | ~x5 | x7);
  assign z012 = n281 | ~n285 | (n152 & ~n284);
  assign n281 = ~x1 & (x3 ? ~n282 : ~n283);
  assign n282 = (x2 | ((~x0 | ~x7 | (x4 ? (x5 | ~x6) : ~x5)) & (x6 | x7 | ((~x4 | ~x5) & (x0 | x4 | x5))))) & (x0 | ~x2 | (x4 ? (x5 | x7) : (x5 ? (x6 | x7) : (~x6 | ~x7))));
  assign n283 = (x0 | ((~x5 | ((x2 | x4 | x6 | x7) & (~x6 | (x2 ? (~x4 | ~x7) : (~x4 ^ x7))))) & (~x2 | x4 | x5 | (~x6 ^ x7)))) & (~x0 | x2 | ~x4 | x5 | x6 | ~x7);
  assign n284 = (~x5 | x6 | x7 | ~x2 | x3 | ~x4) & (x4 | ((~x7 | (x2 ? (x5 | (~x3 ^ x6)) : (~x5 | (~x3 ^ ~x6)))) & (x2 | x3 | ~x5 | ~x6 | x7)));
  assign n285 = (x6 & (x5 ? (x7 & n288) : (~x7 & n286))) | (x5 & ((~x7 & n287) | (~x6 & x7 & n286))) | (~x5 & ((x7 & n287) | (~x6 & ~x7 & n288)));
  assign n286 = (x2 | ((x1 | x3 | ~x4) & (x0 | ~x3 | x4))) & (~x0 | x1 | ~x2 | x3 | x4) & (x0 | (x1 ? ~x3 : (x3 | ~x4)));
  assign n287 = (x0 | ((~x1 | ((~x2 | ~x4 | (~x3 ^ x6)) & (x3 | x4 | x6) & (x2 | (x3 ? (x4 | ~x6) : x6)))) & (~x4 | ~x6 | x1 | ~x3))) & (x1 | ((x2 | ((~x3 | x4 | x6) & (~x0 | x3 | ~x6))) & (x3 | ((x4 | ~x6) & (~x2 | ~x4 | x6)))));
  assign n288 = (x1 | ((x2 | ((~x3 | ~x4) & (~x0 | x3 | x4))) & (~x3 | x4 | x0 | ~x2))) & (x0 | ~x1 | ((x3 | ~x4) & (~x2 | (x3 & ~x4))));
  assign z013 = ~n296 | (x3 ? (x4 ? ~n290 : ~n291) : ~n292);
  assign n290 = (~x6 | ((x1 | ((~x0 | x2 | x5) & (~x5 | x7 | x0 | ~x2))) & (x0 | ~x1 | ((x2 | ~x5 | ~x7) & (x5 | (~x2 & x7)))))) & (x0 | ~x5 | x6 | (~x2 ^ ~x7));
  assign n291 = ((~x5 ^ x6) | ((x2 | ~x7 | ~x0 | x1) & (x0 | ~x1 | ~x2 | x7))) & (x2 | ((x0 | ((x1 | x5 | (~x6 ^ x7)) & (~x6 | x7 | ~x1 | ~x5))) & (~x0 | x1 | x5 | x6 | x7)));
  assign n292 = (x0 | n295) & (n293 | n294);
  assign n293 = ~x5 ^ x7;
  assign n294 = (~x0 | x1 | x2 | ~x4 | ~x6) & (x0 | ~x1 | x4 | (~x2 ^ x6));
  assign n295 = (~x2 | (((~x5 ^ x6) | (x1 ? (~x4 | x7) : ~x7)) & (~x5 | ~x6 | ~x7 | ~x1 | x4))) & (x2 | (((~x1 ^ x5) | (x4 ? (~x6 | ~x7) : (x6 | x7))) & (~x1 | x4 | ~x5 | x6 | ~x7) & (x1 | x5 | ~x6 | x7))) & (x1 | x4 | x5 | ~x6 | x7);
  assign n296 = (n297 | n299) & (x0 | n298) & (~x0 | x1 | n300);
  assign n297 = x4 ? (x5 | x6) : (~x5 | ~x6);
  assign n298 = x7 ? (x1 ? ((~x2 | x3 | ~x4 | ~x5) & (x2 | ~x3 | x4 | x5)) : (~x3 | (x2 ? (~x4 | x5) : ~x5))) : ((x2 | x3 | ~x4 | ~x5) & (x1 | x5 | (x2 ? (~x3 ^ x4) : (~x3 | ~x4))));
  assign n299 = (x7 | ((x1 | (x0 ? (~x2 ^ x3) : (~x2 | ~x3))) & (x0 | ~x1 | ~x2 | x3))) & (x0 | ~x7 | (x3 ? ~x1 : x2));
  assign n300 = (x2 | ((~x5 | x7 | ~x3 | ~x4) & (x3 | ((x5 | x7) & (x4 | ~x5 | ~x7))))) & (x5 | ~x7 | ~x2 | x3);
  assign z014 = ~n308 | (~x2 & ~n307) | (~x1 & ~n302) | (x2 & ~n306);
  assign n302 = (x3 | n305) & (~x3 | x5 | ~x7 | ~n303 | n304);
  assign n303 = ~x0 & ~x2;
  assign n304 = x4 ^ x6;
  assign n305 = (~x5 | x6 | x7 | ~x0 | ~x4) & (x0 | ((x4 | ((~x2 | x7 | (x5 ^ x6)) & (~x6 | ~x7 | x2 | x5))) & (x2 | ~x4 | ~x5 | ~x6 | x7)));
  assign n306 = (x0 | (x3 ? ((x6 | (x1 ? (~x4 ^ x5) : (~x4 | ~x5))) & (x1 | x4 | x5 | ~x6)) : ((x5 | ~x6 | ~x1 | ~x4) & (x1 | x4 | ~x5 | x6)))) & (~x0 | x1 | x3 | x4 | x5 | ~x6);
  assign n307 = (~x5 | ((~x0 | x1 | ~x3 | ~x4 | ~x6) & (x0 | x3 | x4 | x6))) & (x1 | (x0 ? (x3 ? (x4 | x6) : (~x6 | (x4 & x5))) : (x3 ? (x4 | ~x6) : (~x4 | x6)))) & (x0 | ~x1 | (x3 ? (~x4 | x6) : (x4 ^ x6)));
  assign n308 = (n164 | n311) & (~n152 | n309) & (n179 | n310);
  assign n309 = (x2 | x4 | ((~x3 | (x5 ? (x6 | x7) : (~x6 | ~x7))) & (~x6 | x7 | x3 | ~x5))) & (x5 | ~x6 | x7 | ~x2 | ~x3 | ~x4);
  assign n310 = (~x2 | ((x1 | (~x4 ^ x5) | (~x0 ^ x3)) & (x0 | ~x1 | (x3 ? (x4 | x5) : (~x4 | ~x5))))) & (~x3 | ~x4 | ~x5 | x0 | x1 | x2);
  assign n311 = (x0 | ~x2 | (x1 ? (x3 ? (~x4 | ~x5) : x4) : (x3 | ~x4))) & (~x3 | ~x4 | x5 | ~x0 | x1 | x2);
  assign z015 = n313 | n317 | n318 | (~x1 & ~n316);
  assign n313 = ~x2 & (x6 ? ~n315 : ~n314);
  assign n314 = (x1 | ((x5 | (x4 ^ x7) | (x0 ^ ~x3)) & (~x0 | ~x5 | (x3 ? (x4 | ~x7) : (~x4 | x7))))) & (x0 | ~x1 | ((~x7 | (x3 ? (x4 ^ x5) : (x4 | ~x5))) & (x5 | x7 | x3 | ~x4)));
  assign n315 = (x0 | ((x7 | (((~x3 ^ x5) | (x1 ^ ~x4)) & (x1 | x3 | x4 | x5))) & (~x3 | x4 | ~x7 | (~x1 ^ ~x5)))) & (~x4 | ~x5 | ~x7 | ~x0 | x1 | x3);
  assign n316 = (~x4 | (x2 ? ((x7 | ((x3 | x5) & (x0 | (x3 & x5)))) & (~x5 | ~x7 | x0 | ~x3)) : ((~x3 | (x0 ? (x5 ^ x7) : (~x5 | x7))) & (x5 | ~x7 | x0 | x3)))) & (x4 | ((x0 | (x2 ? (~x3 | (~x5 ^ x7)) : (~x5 | ~x7))) & (~x7 | ((x2 | x3 | ~x5) & (~x0 | x5 | (x2 & x3)))) & (~x0 | ~x2 | x3 | ~x5 | x7))) & (x0 | ~x2 | x3 | x5 | x7);
  assign n317 = n152 & ((x5 & ((x3 & ~x4 & (x2 ^ ~x7)) | (x2 & ~x7 & (~x3 | x4)))) | (~x2 & x7 & ((x4 & ~x5) | (~x3 & (x4 | ~x5)))) | (~x5 & ~x7 & x2 & ~x4));
  assign n318 = x2 & ((n196 & n319) | (~x0 & ~n320));
  assign n319 = ~x3 & x0 & ~x1;
  assign n320 = x1 ? ((~x3 | x7 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (~x4 | x5 | x6 | ~x7)) : (x3 | x4 | (x5 ? (~x6 ^ x7) : (~x6 | ~x7)));
  assign z016 = n323 | ~n326 | (~x0 & ~n322);
  assign n322 = x1 ? ((x2 | ((x5 | (x3 ? (~x4 ^ x6) : (~x4 | ~x6))) & (x3 | ~x4 | ~x5 | x6))) & (x4 | ~x5 | ~x6 | ~x2 | ~x3)) : ((x3 | ((~x5 | ~x6 | x2 | ~x4) & (~x2 | (x4 ? (x5 | x6) : (~x5 | ~x6))))) & (x2 | ~x3 | ~x4 | (~x5 ^ x6)));
  assign n323 = ~x1 & ((~x7 & ~n324) | (~x2 & x7 & ~n325));
  assign n324 = x0 ? ((~x2 | x3 | ~x4 | x5 | x6) & (x2 | ~x3 | ~x6 | (x4 ^ x5))) : ((~x2 | x3 | ~x4 | x5 | ~x6) & (x2 | ~x3 | x4 | ~x5 | x6));
  assign n325 = (~x0 | x4 | (x3 ? (~x5 | ~x6) : (x5 | x6))) & (x0 | x3 | ~x4 | ~x5 | x6);
  assign n326 = ~n327 & (~n184 | n330) & (~n152 | (n328 & n329));
  assign n327 = ~x1 & (x0 ? ((x2 & ~x3 & ~x4 & x5) | (~x2 & x3 & x4 & ~x5)) : ((x3 & (x5 ? x2 : ~x4)) | (~x2 & ~x3 & ~x4 & x5)));
  assign n328 = (x6 | (x2 ? (~x3 | ~x5 | (~x4 ^ x7)) : (x3 | x5 | (~x4 ^ ~x7)))) & (~x4 | ~x6 | ~x7 | (x2 ? (x3 | x5) : (~x3 | ~x5)));
  assign n329 = (~x3 | (x2 ? (~x4 | x5) : (x4 | ~x5))) & (~x2 | x3 | (x4 ^ x5));
  assign n330 = (x3 | x4 | ~x5 | x6) & ((~x3 ^ x6) | (~x4 ^ ~x5));
  assign z017 = n332 | (~n164 & ~n336) | (n207 & ~n337);
  assign n332 = ~x0 & ((~x1 & ~n333) | ~n335 | (x1 & ~n334));
  assign n333 = (x3 | ((x5 | x6 | x7 | x2 | ~x4) & (~x5 | (x2 ? (x4 ? (x6 | x7) : ~x6) : (x4 | x6))))) & (x2 | ~x3 | ~x4 | ~x6 | (~x5 & ~x7));
  assign n334 = x2 ? (x5 | ((x3 | ~x4 | ~x6 | ~x7) & (~x3 | x4 | x6 | x7))) : (~x5 | ((~x3 | x4 | x6 | x7) & (x3 | ~x4 | ~x6)));
  assign n335 = (~x1 | ((x2 | ~x3 | ~x6 | ~x7) & (~x2 | x3 | ~x5 | x6))) & (x2 | ~x3 | x5 | ~x6 | x7) & (~x2 | ((x6 | x7 | x3 | x5) & (x1 | ((~x3 | x6 | (x5 & x7)) & (~x6 | ~x7 | x3 | x5)))));
  assign n336 = (x1 | ((x3 | (x0 ? (x5 | (x2 ^ x4)) : (x2 | ~x4))) & (x0 | x2 | ~x3 | x4 | ~x5))) & (x0 | ((~x1 | (x2 ? (~x3 | x4) : (x3 | x5))) & (~x4 | ~x5 | ~x2 | ~x3)));
  assign n337 = (x2 | (x6 ? ((x3 | (~x5 & ~x7)) & (~x7 | (x4 & ~x5))) : ((~x4 | x5 | x7) & (~x3 | (x5 ? x7 : ~x4))))) & (~x2 | x3 | x4 | x6);
  assign z018 = ~n341 | (~x1 & (x6 ? ~n339 : ~n340));
  assign n339 = (x4 | ((~x0 | x3 | ((x5 | x7) & (~x2 | ~x5 | ~x7))) & (x0 | x2 | ~x3 | x5 | ~x7))) & (x0 | ~x3 | ~x4 | ((~x5 | ~x7) & (x2 | x5 | x7)));
  assign n340 = (x0 | ((~x2 | ~x5 | (x3 ? (~x4 ^ x7) : (~x4 | ~x7))) & (x3 | x5 | ((x4 | ~x7) & (x2 | ~x4 | x7))))) & (x2 | x5 | ((~x3 | x4 | x7) & (~x0 | x3 | ~x7)));
  assign n341 = (~n152 | n344) & (x3 | n343) & (~x3 | n342);
  assign n342 = (x0 | ((x7 | (x1 ? (x2 | x5) : (x2 ? x5 : (~x4 | ~x5)))) & (~x1 | ~x5 | ~x7 | (~x2 & ~x4)))) & (x1 | x2 | ((~x7 | ((x4 | ~x5) & (~x0 | (x4 & ~x5)))) & (x5 | x7 | ~x0 | ~x4)));
  assign n343 = (x0 | ((~x1 | (x2 ? (~x5 | x7) : (x5 | ~x7))) & (x4 | ~x5 | x7) & (~x4 | ~x7 | (x5 & (x1 | x2))))) & (x1 | ((~x5 | x7 | (x4 & (~x0 | x2))) & (~x2 | ~x4 | x5 | ~x7)));
  assign n344 = x2 ? (x5 | ((x4 | x6 | (x3 ^ ~x7)) & (~x3 | ~x6 | (~x4 & ~x7)))) : (~x5 | (~x4 ^ x7) | (~x3 ^ x6));
  assign z019 = x0 ? (~x1 & ~n346) : (x1 ? ~n348 : ~n347);
  assign n346 = (x3 | ((~x2 | ((~x5 | x6 | x7) & (~x4 | x5 | ~x6))) & (x4 | ((~x5 | (~x6 ^ x7)) & (x6 | (x7 ? x2 : x5)))))) & (x2 | ((~x5 | (~x6 & (~x3 | ~x7))) & (~x3 | (x4 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n347 = (~x4 & ((~x3 & ((~x5 & x6 & x7) | (~x6 & ~x7))) | (~x6 & (x5 ? ~x2 : ~x7)))) | (x6 & ((~x5 & ((x4 & ~x7) | (~x2 & (x3 | x7)))) | (x2 & ((x4 & x5 & x7) | (x3 & (x7 ? x5 : x4)))) | (x3 & x4 & x5 & x7))) | (~x6 & ((~x5 & (x2 | (x7 & (x3 | x4)))) | (~x2 & ~x3 & x5 & ~x7)));
  assign n348 = (~x6 & ((x2 & (x5 | (x3 & x4 & x7))) | (~x2 & ((~x5 & ~x7) | (~x3 & x4 & x7))) | (~x4 & x5) | (~x3 & x4 & ~x5 & ~x7))) | (x5 & ((x4 & x6 & ~x7) | (~x2 & (x7 | (x3 & x6))))) | (x2 & ~x5 & x6 & ((~x4 & x7) | (x3 & (~x4 | x7))));
  assign z020 = n350 | ~n355 | (~n293 & ~n354) | (n152 & ~n353);
  assign n350 = ~x1 & (x2 ? ~n352 : ~n351);
  assign n351 = x0 ? ((x3 | (x4 ? (~x5 | x6) : (~x6 | ~x7))) & (x5 | x7 | (x4 ^ x6)) & (~x6 | ~x7 | ~x3 | ~x5)) : (x3 | (x4 ? ((x6 | x7) & (~x5 | ~x6 | ~x7)) : ((x6 | ~x7) & (x5 | ~x6 | x7))));
  assign n352 = (x6 | ((~x0 | x3 | x4 | ~x5 | ~x7) & (x0 | ((~x3 | x4 | x5) & (~x4 | ~x5 | ~x7))))) & (x0 | ~x6 | ((~x4 | x5 | x7) & (x3 | (~x4 ^ x7))));
  assign n353 = (x7 | (x2 ? (~x6 | (x3 ? (~x4 | ~x5) : (x4 | x5))) : (x6 | (x3 ? ~x4 : x5)))) & (~x5 | ~x7 | ((x2 | ~x4 | ~x6) & (x6 | (x2 ? (~x3 ^ ~x4) : (~x3 | x4)))));
  assign n354 = x0 ? (x1 | ((x4 | x6 | x2 | x3) & ((~x2 ^ x3) | (~x4 ^ x6)))) : (((~x2 ^ ~x6) | (x1 ? (x3 | ~x4) : (~x3 | x4))) & ((~x1 ^ x4) | (x2 ? (~x3 | x6) : ~x6)) & (~x4 | ~x6 | x2 | ~x3) & (x1 | ~x2 | x3 | x4 | x6));
  assign n355 = (~n356 | n357) & (~n358 | (x1 ^ x2));
  assign n356 = ~x5 & ~x7;
  assign n357 = (~x0 | x1 | ~x2 | x3 | x4) & (x0 | ((x1 | x2 | ~x3 | ~x4) & (~x1 | (x2 ? ~x4 : (~x3 | x4)))));
  assign n358 = x7 & x5 & ~x4 & ~x0 & x3;
  assign z021 = n360 | n364 | n367 | ~n368 | (~n293 & ~n363);
  assign n360 = ~x7 & ((~x0 & ~n362) | (~n361 & (x3 ^ ~x4)));
  assign n361 = (~x0 | x1 | x2 | ~x5 | ~x6) & (x0 | x5 | (x1 ? (x2 | ~x6) : (~x2 | x6)));
  assign n362 = (x3 | (x1 ? ((~x5 | ~x6 | x2 | x4) & (x5 | x6 | ~x2 | ~x4)) : ((x2 | x5 | ~x6) & (~x5 | x6 | ~x2 | x4)))) & (~x4 | ~x5 | x6 | ~x1 | ~x2 | ~x3);
  assign n363 = (x3 | ((x1 | ((~x0 | x4 | (~x2 ^ ~x6)) & (~x4 | x6 | x0 | ~x2))) & (x0 | ~x1 | ((~x2 | x4 | x6) & (~x4 | (x2 & ~x6)))))) & (x0 | x1 | x2 | ~x3 | ~x6);
  assign n364 = ~n365 & n366;
  assign n365 = (~x3 | (x1 ? (~x6 | ((x4 | x5) & (x2 | ~x4 | ~x5))) : (x6 | ((x4 | ~x5) & (~x2 | (x4 & ~x5)))))) & (x1 | x2 | x3 | ~x5 | ~x6);
  assign n366 = ~x0 & x7;
  assign n367 = x3 & n152 & ((~x2 & ~x4 & ~x5 & ~x6) | (x5 & (x2 ? (x4 & x6) : (x4 ^ x6))));
  assign n368 = ~n372 & (n370 | n371) & (n369 | n373);
  assign n369 = x2 ^ x6;
  assign n370 = (~x0 | x1 | x2) & (x0 | ~x1 | ~x2 | x6);
  assign n371 = (x3 | ~x4 | ~x5 | ~x7) & (~x3 | ((x5 | x7) & (x4 | ~x5 | ~x7)));
  assign n372 = ~x1 & ~x3 & ((~x0 & x5 & (x2 ^ ~x6)) | (~x5 & ~x6 & x0 & x2));
  assign n373 = (x0 | (x1 ? (x3 | x4) : (~x3 | ~x4)) | (x5 ^ x7)) & (~x0 | x1 | x3 | ~x4 | x5 | ~x7);
  assign z022 = n375 | n378 | ~n379 | n384 | (~n179 & ~n383);
  assign n375 = ~x1 & (x3 ? (x7 & ~n377) : ~n376);
  assign n376 = (~x5 | ((~x0 | ((x2 | x4 | ~x6 | ~x7) & (x6 | x7 | ~x2 | ~x4))) & (x0 | ~x2 | x4 | ~x6 | x7))) & (x5 | ~x6 | ~x7 | x0 | x2 | x4);
  assign n377 = (x0 | x6 | (x2 ? (~x4 | x5) : (x4 | ~x5))) & (~x0 | x2 | ~x4 | x5 | ~x6);
  assign n378 = ~n164 & ((x0 & ~x1 & ~x2 & ~x3 & ~x4) | (~x0 & x2 & (x1 ? (x3 & x4) : (x3 ^ x4))));
  assign n379 = ~n381 & (x0 | (n382 & (~x1 | x7 | n380)));
  assign n380 = (x2 | x3 | ~x4 | x5 | ~x6) & (~x2 | ~x3 | x4 | (x5 ^ x6));
  assign n381 = ~x0 & x1 & ~x3 & (x2 ? ~x6 : (~x4 & x6));
  assign n382 = (x1 | x2 | ~x3 | x4 | x6 | x7) & (~x1 | ~x7 | ((x2 | x3 | ~x4 | ~x6) & (~x2 | ~x3 | x4 | x6)));
  assign n383 = (x1 | ((~x3 | ~x4 | ~x5 | ~x0 | x2) & (x3 | (x0 ? (~x2 | (x4 & x5)) : (x2 | (~x4 & ~x5)))))) & (x0 | ~x1 | x2 | ~x3);
  assign n384 = ~x1 & ((~x2 & ((x0 & x6 & (x3 ^ x4)) | (x4 & ~x6 & ~x0 & x3))) | (~x0 & x2 & (x3 ? (x4 & x6) : (~x4 & ~x6))));
  assign z023 = n394 | ~n395 | (~x1 & (~n386 | n387 | ~n391));
  assign n386 = ((x2 ? (x3 | x5) : (~x3 | ~x5)) | (x0 ? (~x4 | x7) : (x4 | ~x7))) & (x0 | ((~x2 | ~x3 | ~x4 | ~x5 | ~x7) & (x2 | x4 | x7 | (~x3 ^ x5))));
  assign n387 = ~n164 & ((n388 & n390) | (n171 & n389));
  assign n388 = x3 & x4 & ~x5;
  assign n389 = x5 & ~x3 & ~x4;
  assign n390 = x0 & ~x2;
  assign n391 = (x0 | x5 | ((~x3 | n392) & (~x6 | n393))) & (~x5 | n392 | ~x0 | x3);
  assign n392 = (~x2 | ~x4 | x6 | x7) & (x2 | x4 | ~x6 | ~x7);
  assign n393 = (~x2 | ~x3 | ~x4 | ~x7) & (x2 | x3 | x4 | x7);
  assign n394 = ~x1 & (x0 ? ((~x3 & ~x4 & ~x7) | (~x2 & x7 & (x3 ^ x4))) : (x3 ? (x2 ? (~x4 & ~x7) : (x4 & x7)) : (x4 & ~x7)));
  assign n395 = ~n397 & (~n152 | (n396 & (~n264 | ~n272 | ~n260)));
  assign n396 = (x2 | x3 | ~x4 | x5 | ~x7) & (~x2 | ~x3 | x4 | (~x5 ^ x7));
  assign n397 = ~x0 & x1 & (x3 ? (~x7 & (~x2 | x4)) : (x7 & (x2 | ~x4)));
  assign z024 = n399 | n402 | n403 | ~n407 | (n147 & ~n401);
  assign n399 = ~x1 & ~n400;
  assign n400 = (x4 | ~x5 | ~x6 | x0 | ~x2 | x3) & (x5 | (x0 ? ((x2 | ~x3 | ~x4 | ~x6) & (~x2 | x3 | x4 | x6)) : ((~x2 | ~x3 | ~x4 | ~x6) & (x2 | x3 | (~x4 ^ x6)))));
  assign n401 = (x5 | ~x6 | ~x7 | x1 | x2 | x4) & (~x5 | x7 | ((~x1 | (x2 ? (~x4 | x6) : (x4 | ~x6))) & (x1 | x2 | ~x4 | x6)));
  assign n402 = ~x0 & ((~x5 & ((~x1 & ~x2 & x3 & x4) | (x1 & (x2 ? (x3 & x4) : ~x4)))) | (~x1 & ~x2 & ~x4 & x5));
  assign n403 = ~x3 & ((~n405 & ~n406) | (n271 & n265 & n404));
  assign n404 = ~x2 & ~x0 & ~x1;
  assign n405 = x2 ? (x5 | x7) : (~x5 | ~x7);
  assign n406 = (x0 | ~x1 | ~x4 | x6) & (x4 | ~x6 | ~x0 | x1);
  assign n407 = ~n409 & (~n152 | ~n408 | (x3 ? (x4 | x6) : (~x4 | ~x6)));
  assign n408 = ~x2 & x5;
  assign n409 = (~x3 | x5) & ((~x0 & x2 & (x1 ^ x4)) | (~x2 & x4 & x0 & ~x1));
  assign z025 = ~n413 | (~x1 & (x2 ? ~n412 : ~n411));
  assign n411 = x3 ? ((x0 | ~x7 | (x4 ? (~x5 | x6) : (x5 | ~x6))) & (~x5 | x6 | x7 | ~x0 | x4)) : ((~x6 | ((~x5 | x7 | x0 | ~x4) & (~x0 | (x4 ? (x5 | x7) : (~x5 | ~x7))))) & (x0 | x4 | x6 | (~x5 ^ x7)));
  assign n412 = (x0 | x7 | ((x5 | ~x6 | x3 | ~x4) & (~x3 | ~x5 | (x4 ^ x6)))) & (x5 | ~x6 | ~x7 | ~x0 | x3 | x4);
  assign n413 = (~x4 | n416) & (x4 | n415) & (~n152 | n414);
  assign n414 = (~x5 | ((~x7 | ((x2 | (x3 ? (x4 | ~x6) : (~x4 | x6))) & (~x2 | ~x3 | ~x4 | x6))) & (~x2 | x3 | x7 | (x4 ^ x6)))) & (~x4 | x5 | ((x2 | ~x3 | ~x6 | x7) & (~x2 | x6 | (x3 ^ ~x7))));
  assign n415 = (x1 | ((x3 | ((x5 | ~x6 | x0 | x2) & (~x2 | ~x5 | (~x0 & ~x6)))) & (~x3 | x5 | x0 | ~x2) & (x2 | (x0 ? (x5 | (~x3 & x6)) : (~x3 | ~x5))))) & (x0 | ((~x1 | (x2 ? (x3 ^ x5) : (x3 ? (x5 | x6) : ~x5))) & (x5 | x6 | ~x2 | x3)));
  assign n416 = ((~x5 ^ x6) | ((x2 | ~x3 | ~x0 | x1) & (x0 | (x1 ? (~x2 | x3) : (x2 ^ x3))))) & (x0 | (x1 ? ((x2 | (x3 ? (x5 | x6) : (~x5 | ~x6))) & (~x5 | ~x6 | ~x2 | ~x3)) : ((~x5 | ~x6 | x2 | ~x3) & (x5 | x6 | ~x2 | x3)))) & (x3 | x5 | x6 | ~x0 | x1 | x2);
  assign z026 = ~n419 | n429 | (~x5 & ~n424) | (~x1 & ~n418);
  assign n418 = (x2 | (x3 ? ((~x4 | ~x5 | ~x6) & (x5 | x6 | ~x0 | x4)) : ((~x0 | (x4 ? (~x5 | x6) : (x5 | ~x6))) & (x5 | ~x6 | x0 | ~x4)))) & (x0 | ~x2 | (x3 ? (x5 | (x4 ^ x6)) : (x4 ? (~x5 | x6) : ~x6)));
  assign n419 = (~n152 | n423) & (n420 | n421) & (n182 | n422);
  assign n420 = x5 ? (x6 | ~x7) : (~x6 | x7);
  assign n421 = (x0 | ((~x1 | ~x2 | x3 | x4) & (x1 | ~x3 | (~x2 ^ x4)))) & (x2 | ~x3 | x4 | ~x0 | x1);
  assign n422 = (x1 | ((~x0 | (x2 ? (x3 | x6) : (~x3 | ~x6))) & (~x3 | x6 | x0 | x2))) & (x0 | ~x1 | x3 | (x2 ^ x6));
  assign n423 = (x4 | ((~x2 | x6 | (~x3 ^ ~x5)) & (x2 | ~x3 | x5 | ~x6))) & (x2 | ~x3 | ~x4 | ~x5 | x6);
  assign n424 = (~n425 | ~n428) & (n179 | n426) & (x3 | n427);
  assign n425 = ~x6 & (x4 ^ ~x7);
  assign n426 = (x1 | ((~x3 | x4 | x0 | x2) & (x3 | (x0 ? (~x2 ^ x4) : (~x2 | ~x4))))) & (x0 | ~x1 | x2 | ~x3 | ~x4);
  assign n427 = (x0 | x6 | ((~x1 | (x2 ? (~x4 | ~x7) : (x4 | x7))) & (x1 | x2 | x4 | ~x7))) & (~x4 | ~x6 | x7 | ~x0 | x1 | ~x2);
  assign n428 = x3 & x2 & ~x0 & x1;
  assign n429 = x5 & ((~x0 & ~n430) | (n153 & n431));
  assign n430 = ((~x2 ^ ~x3) | ((x1 | x4 | ~x6 | x7) & (~x4 | (x1 ? (~x6 ^ x7) : (~x6 | ~x7))))) & (~x7 | ((~x1 | ~x6 | (x2 ? (x3 | ~x4) : (~x3 | x4))) & (x1 | x2 | x3 | x4 | x6)));
  assign n431 = x7 & x6 & ~x3 & ~x4;
  assign z027 = ~n444 | n443 | n441 | n438 | n433 | n435;
  assign n433 = ~x0 & ~n434;
  assign n434 = x3 ? ((~x1 | ~x2 | x4 | ~x5 | x7) & (x2 | x5 | (x1 ? (x4 ^ x7) : (x4 | ~x7)))) : ((~x1 | ((x2 | x7 | (~x4 ^ x5)) & (x5 | ~x7 | ~x2 | x4))) & (~x5 | ~x7 | x2 | ~x4) & (x1 | (x2 ? (~x4 | (~x5 ^ x7)) : (~x5 | ~x7))));
  assign n435 = x2 & ((~x3 & ~n436) | (x3 & ~x5 & n152 & ~n437));
  assign n436 = (x1 | ((x0 | x4 | ~x5 | ~x6 | ~x7) & (x5 | x6 | x7 | ~x0 | ~x4))) & (x0 | ~x1 | ((~x4 | x5 | x6 | ~x7) & (x4 | ~x5 | (~x6 ^ x7))));
  assign n437 = x4 ? (~x6 | x7) : (x6 | ~x7);
  assign n438 = ~x2 & (x7 ? (n152 & ~n440) : ~n439);
  assign n439 = (x1 | ((x3 | ((x0 | x4 | x5 | ~x6) & (~x0 | (x4 ? ~x6 : (~x5 | x6))))) & (x0 | ~x3 | (x4 ? (x5 | x6) : (~x5 | ~x6))))) & (x0 | ~x1 | ~x3 | ~x5 | (x4 ^ x6));
  assign n440 = (x3 | x5 | (~x4 ^ ~x6)) & (~x5 | x6 | ~x3 | x4);
  assign n441 = ~n198 & ~n442;
  assign n442 = (~x0 | x1 | x2 | ~x3 | x4 | ~x7) & (x0 | ~x4 | ((x7 | (x1 ? (~x2 | x3) : (x2 ^ x3))) & (x1 | x2 | ~x3 | ~x7)));
  assign n443 = ~x3 & n207 & ((x2 & ((~x5 & x7) | (~x4 & x5 & ~x7))) | (x4 & ~x5 & x7) | (~x2 & ~x4 & (~x5 ^ x7)));
  assign n444 = ~n445 & ~n446 & (n449 | (~n447 & ~n448));
  assign n445 = x3 & ((~x0 & x2 & x7 & (x1 ^ ~x4)) | (x0 & ~x1 & ~x2 & x4 & ~x7));
  assign n446 = ~x7 & ~x4 & ~x3 & x2 & ~x0 & ~x1;
  assign n447 = x4 & x5 & x6 & x7;
  assign n448 = ~x7 & ~x6 & ~x4 & ~x5;
  assign n449 = (x2 | ~x3 | ~x0 | x1) & (x0 | ~x2 | (x1 ^ ~x3));
  assign z028 = n451 | (~n179 & ~n455) | (n152 & ~n456);
  assign n451 = ~x1 & ((x3 & ~n452) | ~n454 | (~x3 & ~n453));
  assign n452 = (x2 | ((~x0 | ((~x5 | ~x6 | x7) & (~x4 | x5 | x6 | ~x7))) & (~x5 | ((~x4 | ~x6 | x7) & (x0 | x6 | (~x4 ^ ~x7)))) & (x0 | x4 | x5 | x6 | ~x7))) & (~x5 | ~x6 | ~x7 | x0 | ~x2 | x4);
  assign n453 = (x0 | ((~x2 | ((~x6 | ~x7 | ~x4 | ~x5) & (x4 | ((~x6 | x7) & (~x5 | x6 | ~x7))))) & (x2 | x4 | x5 | x6 | ~x7))) & (x2 | ~x4 | ~x5 | x6 | x7) & (~x0 | ((x5 | ~x7 | (x2 ? (x4 | x6) : (~x4 ^ x6))) & (x6 | x7 | ~x4 | ~x5)));
  assign n454 = x3 ? ((x6 | ((x2 | (~x0 ^ (x4 & ~x5))) & (x0 | ~x2 | ~x4 | ~x5))) & (~x0 | x2 | ~x4 | x5 | ~x6)) : (~x6 | (x0 ? (~x2 | x4) : (x2 ? (~x4 | x5) : x4)));
  assign n455 = (x1 | ((x3 | ((x2 | ~x4 | x5) & (~x0 | ((~x4 | x5) & (x2 | x4 | ~x5))))) & (x0 | ~x3 | x5 | (~x2 & x4)))) & (x0 | ~x1 | x2 | ~x3 | ~x5);
  assign n456 = (~x3 & ((x2 & (x6 | (~x4 & ~x5 & x7))) | (x6 & (x5 ? ~x4 : x7)))) | (~x6 & ((~x2 & (x3 | (x5 & ~x7))) | (x3 & (x4 | x5 | ~x7)))) | (~x2 & x3 & x5) | (x6 & x7 & x2 & ~x5);
  assign z029 = ~n461 | (~x1 & (~n460 | (x2 ? ~n459 : ~n458)));
  assign n458 = (~x6 | ((x5 | ((x4 | ((x3 | x7) & (x0 | (x3 & x7)))) & (~x0 | ~x3 | ~x4 | ~x7))) & (~x0 | ~x5 | (x3 ? x7 : (~x4 | ~x7))))) & (x5 | x6 | ~x7 | (~x0 ^ x3));
  assign n459 = (~x5 | x6 | x7 | ~x0 | x3 | ~x4) & (x0 | ((~x5 | (~x6 ^ x7) | (~x3 ^ x4)) & (x3 | x5 | x6 | (x4 & x7))));
  assign n460 = x0 ? ((x3 | (x2 ? (x4 ? (x5 | x7) : (~x5 | ~x7)) : (~x5 | x7))) & (x2 | ~x3 | x5 | (~x4 ^ x7))) : (x3 ? ((~x5 | x7 | x2 | ~x4) & (~x2 | ((x5 | x7) & (~x4 | ~x5 | ~x7)))) : (x2 ? (x4 ? (x5 | ~x7) : (~x5 | x7)) : (x4 ? (x5 | x7) : (~x5 | ~x7))));
  assign n461 = (n179 | n464) & (~n152 | (n462 & n463));
  assign n462 = x3 ? ((x2 | x4 | ~x5 | ~x6 | ~x7) & (~x2 | ((~x4 | x5 | (~x6 ^ x7)) & (x6 | x7 | x4 | ~x5)))) : (x2 ? (x6 | ((~x5 | ~x7) & (~x4 | x5 | x7))) : (~x6 | ((x5 | x7) & (~x4 | ~x5 | ~x7))));
  assign n463 = (~x4 | ((x2 | ~x5 | x7) & (x5 | ~x7 | ~x2 | x3))) & (~x3 | (x2 ? ((~x5 | ~x7) & (x4 | x5 | x7)) : (~x5 ^ x7)));
  assign n464 = (x0 | ((x3 | ((x1 | x2 | ~x4 | ~x5) & (~x1 | x4 | (~x2 ^ x5)))) & (x1 | x2 | ~x3 | x4 | ~x5))) & (~x0 | x1 | ~x2 | x3 | x4 | x5);
  assign z030 = ~n474 | (~x1 & (~n467 | (~x0 & ~n466)));
  assign n466 = (x5 | x7 | (x2 ? (x3 ? x6 : (x4 | ~x6)) : (x3 ? (x4 | ~x6) : (~x4 | x6)))) & (x3 | ~x4 | ~x5 | ~x6 | ~x7);
  assign n467 = ~n468 & ~n469 & ~n472 & ~n473 & (n470 | ~n471);
  assign n468 = ~x2 & ((x3 & ~x5 & (x4 ? (x6 & x7) : (~x6 & ~x7))) | (~x3 & ~x4 & x5 & ~x6 & ~x7));
  assign n469 = ~x2 & ((x0 & x7 & (x3 ? (~x4 & ~x6) : (x4 & x6))) | (x4 & x6 & ~x7 & ~x0 & ~x3));
  assign n470 = (x2 | ~x3 | ~x5) & (~x4 | x5 | ~x2 | x3);
  assign n471 = x0 & x6 & ~x7;
  assign n472 = ~x0 & x2 & ~x3 & (x4 ? (x6 & ~x7) : (~x6 & x7));
  assign n473 = ~x7 & ~x6 & x5 & ~x4 & x2 & ~x3;
  assign n474 = (n215 | n475) & (~n152 | n476);
  assign n475 = x3 ? (~x5 | ((x1 | (x0 & (x2 | ~x7))) & (x0 | (x2 & x7)))) : (x5 | (x0 ? x1 : ~x7));
  assign n476 = x6 ? ((~x4 | (x3 ? (~x5 | x7) : ~x7)) & (x3 | ((x5 | x7) & (~x2 | ~x5 | ~x7)))) : ((~x3 | (x7 ? ((x4 | ~x5) & (~x2 | (x4 & ~x5))) : ((x4 | x5) & (x2 | (x4 & x5))))) & (x2 | x3 | x4 | x5 | ~x7));
  assign z031 = n478 | ~n483 | (~x2 & ~n480) | (~x0 & ~n482);
  assign n478 = ~n179 & ~n479;
  assign n479 = (x1 | ((~x0 | x3 | (x2 ? x5 : (~x4 | ~x5))) & (x2 | ~x4 | x5 | (x0 & ~x3)))) & (x0 | ~x5 | ((~x2 | ~x4) & (~x1 | (x2 & x3))));
  assign n480 = (x1 | n481) & (x0 | ~x1 | ~n264 | (~n388 & ~n186));
  assign n481 = (~x3 | ((~x0 | ((~x4 | ~x5 | ~x7) & (x6 | x7 | x4 | x5))) & (~x5 | x6 | x7 | x0 | ~x4))) & (x0 | ~x7 | ((x4 | x5 | ~x6) & (x3 | x6 | (~x4 ^ x5))));
  assign n482 = (~x6 | x7 | x1 | ~x5) & (x5 | ~x7 | (x1 ? (x2 | x6) : (x3 ? x6 : ~x2)));
  assign n483 = (~n153 | ~n486) & (~n171 | n484) & (n420 | n485);
  assign n484 = (~x1 | ((~x3 | ((~x6 | ~x7 | x4 | ~x5) & (x6 | x7 | ~x4 | x5))) & (x3 | ~x4 | x5 | x6 | ~x7))) & (~x5 | x6 | x7 | x1 | ~x3 | x4);
  assign n485 = x0 ? (x1 | ((x3 | x4) & (x2 | (x3 & x4)))) : (~x1 | (~x2 & (~x3 | x4)));
  assign n486 = ~x7 & ~x6 & ~x3 & ~x5;
  assign z032 = ~n490 | (~x1 & (x2 ? ~n489 : ~n488));
  assign n488 = x5 ? (x0 ? ((~x3 | (x4 ? ~x6 : (x6 | ~x7))) & (x3 | ~x4 | x6 | x7)) : ((x4 | x6 | x7) & (x3 | ~x6 | (~x4 ^ x7)))) : ((~x0 | ~x7 | (~x4 ^ x6)) & (x0 | ~x3 | ~x4 | x6 | x7));
  assign n489 = (~x0 | x3 | ~x4 | x5 | x6 | ~x7) & (x0 | ((x3 | ((x6 | x7 | x4 | ~x5) & (~x6 | ~x7 | ~x4 | x5))) & (~x7 | (x4 ? (~x5 | x6) : ((x5 | x6) & (~x3 | ~x5 | ~x6))))));
  assign n490 = x1 ? (x0 | (n492 & n493)) : n491;
  assign n491 = (~x6 | ((x7 | ((~x0 | x2 | (x3 & x4)) & (~x2 | x3 | x4) & (x0 | (~x2 & (~x3 | ~x4))))) & (x2 | x3 | ~x4 | ~x7) & (x0 | (x2 ? (x3 | x4) : (~x3 | ~x7))))) & (x3 | x6 | (x0 ^ x2) | (~x4 ^ x7));
  assign n492 = (x6 | ((x3 | (~x2 ^ x7)) & (x2 | (x4 ^ x7)))) & (~x2 | ~x6 | ~x7 | (~x3 & x4));
  assign n493 = x7 ? ((~x2 | x3 | ~x4 | (x5 ^ x6)) & (x2 | ~x3 | x4 | x5 | x6)) : ((~x3 | ((~x4 | ~x5 | x6) & (~x2 | x4 | (x5 ^ x6)))) & (x2 | x3 | ~x6 | (~x4 ^ x5)));
  assign z033 = ~n496 | ~n499 | (~n495 & (n152 | n207));
  assign n495 = (x3 | ((~x2 | (x4 ? (x5 | ~x7) : x7)) & (x5 | x7 | x2 | ~x4))) & (x2 | (x4 ? (~x5 | ~x7) : ((x5 | ~x7) & (~x3 | ~x5 | x7))));
  assign n496 = (n179 | n497) & (x5 | ~n147 | n498);
  assign n497 = (x1 | x2 | ~x3 | ~x4 | x5) & (x0 | ((x2 | ~x3 | ~x4 | x5) & (x1 | ~x2 | x3 | x4 | ~x5)));
  assign n498 = (~x2 | ~x4 | (~x6 ^ x7)) & (x1 | x2 | x4 | x6 | ~x7);
  assign n499 = (x0 | n501) & (~n500 | n502);
  assign n500 = ~x3 & x5;
  assign n501 = ((~x4 ^ x7) | ((~x2 | ~x3 | ~x5) & (x1 | x2 | x3 | x5))) & (x1 | (x2 ? (x5 | ((x4 | x7) & (x3 | ~x4 | ~x7))) : (~x5 | ((~x4 | ~x7) & (~x3 | x4 | x7))))) & (~x2 | ~x3 | x4 | x5 | x7);
  assign n502 = x2 ? (~x6 | ((x0 | ((~x4 | x7) & (~x1 | x4 | ~x7))) & (~x0 | x1 | x4 | ~x7))) : ((x0 | x4 | ~x6 | x7) & (x6 | (x0 & x1) | (~x4 ^ x7)));
  assign z034 = ~n508 | (~x1 & (n505 | ~n506 | (x5 & ~n504)));
  assign n504 = (~x0 | x4 | ~x6 | ((x3 | x7) & (x2 | ~x3 | ~x7))) & (x0 | ~x2 | ~x3 | ~x4 | x6 | ~x7);
  assign n505 = ~x3 & ((~x6 & ~x7 & x4 & x5) | (~x5 & x6 & x7 & x2 & ~x4));
  assign n506 = ~n507 & (~x6 | ~n271 | ~n303 | (x3 ^ ~x7));
  assign n507 = x7 & ~x6 & x5 & x4 & ~x2 & x3;
  assign n508 = ~n510 & (~x5 | ~n152 | n509) & (~x3 | n511);
  assign n509 = x3 ? (~x7 | (~x4 ^ x6)) : (x7 | ((~x4 | x6) & (~x2 | x4 | ~x6)));
  assign n510 = ~x3 & (~x0 | ~x1) & (x4 ? (~x5 & x6) : (x5 & ~x6));
  assign n511 = (x1 & (x0 | (~x4 & x5))) | (x0 & (x2 | (~x4 & x5))) | (x5 & ~x6) | (~x5 & x6 & (x4 | (~x0 & ~x1 & ~x2)));
  assign z035 = (~x0 & (x1 ? ~n514 : ~n515)) | ~n516 | (x0 & ~x1 & ~n513);
  assign n513 = (~x7 | ((x6 | (x2 & x3) | (~x4 ^ x5)) & (x5 | ~x6 | x2 | x4))) & (x2 | ~x4 | ~x5 | (x7 & (~x3 | ~x6)));
  assign n514 = (x6 | (x4 ? ((x5 | ~x7) & (~x2 | ~x3 | ~x5 | x7)) : (~x5 | ~x7))) & (x4 | x5 | ~x6 | ((x2 | x3) & ~x7));
  assign n515 = (~x4 | x5 | x6 | ~x7) & (x4 | ((~x2 | ((~x3 | x5 | ~x6) & (~x5 | x6 | ~x7))) & (x5 | ~x6 | x7) & (x6 | ~x7 | ~x3 | ~x5)));
  assign n516 = x7 ? n518 : n517;
  assign n517 = ((x2 & x3) | ((~x0 | x1 | x4 | ~x6) & (x0 | ~x4 | x6))) & (x1 | ~x2 | x3 | ~x4 | x6) & (x0 | (x1 ? (x4 | ~x6 | (~x2 & ~x3)) : (~x4 | x6)));
  assign n518 = (x0 | ((~x4 | ~x6) & (x1 | x2 | x3 | x4 | x6))) & (x1 | x2 | x3 | ~x4 | ~x6);
  assign z036 = ~n529 | n528 | n526 | n524 | n520 | n522;
  assign n520 = ~x2 & ~n521;
  assign n521 = (x1 | (x0 ? (~x4 | ((x6 | x7) & (~x5 | ~x6 | ~x7))) : (x4 | x7 | (~x5 ^ x6)))) & (x0 | ((~x4 | x5 | x6 | ~x7) & (~x6 | ((x4 | ~x5 | ~x7) & (~x1 | ((~x5 | ~x7) & (~x4 | x5 | x7)))))));
  assign n522 = ~n523 & ~x1 & x7;
  assign n523 = (~x4 | x5 | x6 | ~x0 | x2 | x3) & (x4 | ((~x2 | x3 | x5 | x6) & (x0 | ((~x5 | ~x6 | ~x2 | x3) & (x2 | ~x3 | x5 | x6)))));
  assign n524 = ~x4 & ~n525;
  assign n525 = (x1 | ((~x0 | x2 | ((x5 | ~x7) & (x3 | ~x5 | x7))) & (~x3 | ~x7 | x0 | ~x2))) & (x0 | ((~x2 | ~x3 | x5 | ~x7) & (~x1 | ((x2 | x3 | x5 | ~x7) & (~x2 | ~x3 | ~x5 | x7)))));
  assign n526 = ~n527 & (x0 ? (~x1 & (x4 ? (~x5 & x7) : (x5 & ~x7))) : ((x4 & x5 & ~x7) | (x1 & ((x5 & ~x7) | (~x4 & ~x5 & x7)))));
  assign n527 = ~x2 ^ x3;
  assign n528 = n171 & ((~x1 & ~x4 & x5 & ~x6 & ~x7) | (x4 & x7 & ((~x5 & ~x6) | (x1 & x5 & x6))));
  assign n529 = (n531 | ~n532) & (~n264 | ~n530 | ~n248 | ~n152);
  assign n530 = x4 & ~x5;
  assign n531 = x2 ? (~x3 | (~x1 & ~x5)) : (x3 | ~x5);
  assign n532 = ~x7 & ~x0 & x4;
  assign z037 = ~n544 | n542 | n540 | n538 | n534 | n536;
  assign n534 = ~x1 & ((~x0 & ~n535) | (n260 & n265 & x0 & n247));
  assign n535 = (~x3 | ((x2 | x4 | ~x5 | x6 | ~x7) & (x5 | ~x6 | x7 | (~x2 & ~x4)))) & (~x2 | ((~x4 | (x5 ? (x6 | ~x7) : (~x6 | x7))) & (x6 | ~x7 | x3 | ~x5)));
  assign n536 = ~x0 & ~n537;
  assign n537 = (~x3 | ((~x1 | ((~x5 | x6 | ~x2 | ~x4) & (x2 | x4 | x5 | ~x6))) & (x5 | x6 | x1 | ~x4))) & (x1 | ((~x4 | ((~x5 | ~x6) & (~x2 | x5 | x6))) & (x2 | x3 | x4 | ~x5 | x6)));
  assign n538 = ~n539 & (n245 | n246);
  assign n539 = (x0 | ~x1 | x2 | x3 | x4) & (x1 | (x0 ? (~x4 | (~x2 ^ x3)) : (x4 | (~x2 & ~x3))));
  assign n540 = ~n541 & (x4 ^ x7);
  assign n541 = (x0 | ~x1 | ~x2 | ((~x5 | ~x6) & (~x3 | x5 | x6))) & (~x0 | x1 | x2 | x5 | x6);
  assign n542 = ~n164 & ~n543;
  assign n543 = (~x0 | x1 | ~x2 | x3 | x4 | x5) & (x0 | x2 | ~x4 | (x1 ? ~x5 : (x3 | x5)));
  assign n544 = n548 & (n546 | n547) & (~n272 | ~n152 | ~n545);
  assign n545 = ~x7 & x6 & ~x4 & ~x5;
  assign n546 = x2 ? (x4 | ~x6) : (~x4 | x6);
  assign n547 = (x0 | ~x1 | x5) & (x3 | ~x5 | ~x0 | x1);
  assign n548 = (~x0 | x1 | x2 | x4 | ~x6) & (x3 | ~x4 | x6 | x0 | ~x1 | ~x2);
  assign z038 = n551 | ~n554 | (~x3 & ~n550);
  assign n550 = (x1 | ((~x0 | x5 | x7 | (~x2 ^ x4)) & (~x5 | ~x7 | ((~x2 | x4) & (x0 | x2 | ~x4))))) & (x0 | ~x1 | ((x2 | ~x5 | x7) & (x5 | ~x7 | (~x2 & x4))));
  assign n551 = ~x1 & ((n171 & ~n553) | (~x2 & ~n552));
  assign n552 = x0 ? ((x3 | x4 | x5 | x6 | x7) & (~x3 | ~x5 | ~x7 | (~x4 ^ x6))) : ((x3 | ((~x6 | ~x7 | x4 | ~x5) & (x6 | x7 | ~x4 | x5))) & (x4 | x5 | ~x6 | x7));
  assign n553 = x5 ? ((~x3 | x4 | x6 | x7) & (~x6 | ((~x4 | ~x7) & (~x3 | (~x4 & ~x7))))) : (x6 | ~x7);
  assign n554 = (~n152 | n557) & (n198 | n555) & (~n247 | n556);
  assign n555 = (x1 | ((x2 | ~x7 | ((x3 | x4) & (~x0 | (x3 & x4)))) & (x7 | ((~x2 | x3 | ~x4) & (x0 | (~x4 & (~x2 | x3))))))) & (x0 | ~x1 | ~x2 | ~x3 | ~x7);
  assign n556 = (~x0 | x1 | x5 | x7) & (x0 | (x1 ? ((x5 | ~x7) & (~x4 | ~x5 | x7)) : (~x5 | ~x7)));
  assign n557 = (x2 | ~x7 | ((x4 | ~x5 | ~x6) & (x3 | ~x4 | x5 | x6))) & (x7 | ((~x2 | ((~x5 | ~x6) & (x4 | x5 | x6))) & (~x3 | ((x4 | ~x5 | ~x6) & (~x2 | x5 | x6)))));
  assign z039 = n559 | n563 | n565 | ~n567 | (~n164 & ~n562);
  assign n559 = ~x0 & (x2 ? ~n561 : ~n560);
  assign n560 = (x4 | (x1 ? ((~x5 | ~x6 | ~x7) & (x6 | x7 | x3 | x5)) : (x5 | ~x7 | (~x3 ^ x6)))) & (~x5 | ~x6 | ~x7 | x1 | ~x3 | ~x4);
  assign n561 = (x3 | x4 | ~x6 | (x1 ? (~x5 | ~x7) : (x5 | x7))) & (~x1 | ~x4 | x5 | x7 | (~x3 & x6));
  assign n562 = (~x0 | x1 | ~x2 | x3 | ~x4 | x5) & (x0 | ((~x1 | ((~x2 | x3) & (x2 | ~x3 | x4 | ~x5))) & (~x2 | x3 | x4 | ~x5) & (x1 | x2 | ~x4 | (~x3 & ~x5))));
  assign n563 = ~n179 & ~n564;
  assign n564 = (x1 | ((~x3 | (x4 ^ x5) | (x0 ^ ~x2)) & (~x0 | x2 | x3 | (~x4 ^ x5)))) & (x3 | ~x4 | x5 | x0 | ~x1 | x2);
  assign n565 = ~x1 & ~n566;
  assign n566 = (x2 | ((x5 | ((~x0 | (x3 ? (~x4 | x6) : (x4 | ~x6))) & (x0 | x3 | ~x4 | x6))) & (x4 | ~x5 | x6 | (x0 & ~x3)))) & (x0 | ~x2 | ~x3 | ~x6 | (~x4 ^ x5));
  assign n567 = ~n569 & ~n570 & (~n261 | ~n447) & (~n152 | n568);
  assign n568 = (x2 | x6 | (x3 ? (x4 | x5) : ~x5)) & (~x2 | ~x3 | ~x4 | ~x5 | ~x6);
  assign n569 = ~x0 & ((~x1 & x2 & ~x3 & x4 & x6) | (x1 & x3 & (x2 ? (~x4 & x6) : (x4 & ~x6))));
  assign n570 = ~x6 & ~x4 & ~x3 & x2 & x0 & ~x1;
  assign z040 = n572 | n575 | (x7 ? ~n579 : ~n578);
  assign n572 = x2 & ((n319 & n573) | (~x0 & ~n574));
  assign n573 = x7 & x6 & ~x4 & x5;
  assign n574 = (x5 | ((~x6 | (x1 ? (x3 ? (x4 | x7) : (~x4 | ~x7)) : (x3 ? (~x4 | ~x7) : (~x4 ^ x7)))) & (~x1 | x3 | ~x4 | x6 | x7))) & (~x1 | x3 | x4 | ~x5 | (~x6 ^ x7));
  assign n575 = ~x2 & ((~x1 & ~n576) | (n152 & ~n577));
  assign n576 = x0 ? ((x3 | ~x4 | x6 | (~x5 ^ x7)) & (~x6 | ((~x3 | x4 | ~x5 | x7) & (x3 | (x4 ? (x5 ^ x7) : (x5 | ~x7)))))) : ((x3 | x4 | ~x5 | ~x6 | x7) & (~x3 | ((~x6 | ~x7 | x4 | ~x5) & ((x4 ^ x5) | (~x6 ^ x7)))));
  assign n577 = (~x5 | ((~x6 | (x3 ? (~x4 | ~x7) : (~x4 ^ x7))) & (x3 | x4 | x6 | x7))) & (x3 | x4 | x5 | (~x6 ^ x7));
  assign n578 = (x0 | ((~x3 | ((~x1 | (x5 ? ~x4 : x2)) & (~x2 | x4 | ~x5) & (x1 | ((x4 | ~x5) & (~x2 | ~x4 | x5))))) & (x1 | x3 | ~x4 | (~x2 ^ ~x5)))) & (x1 | ((x3 | x4 | ((~x2 | x5) & (~x0 | (~x2 & x5)))) & (~x3 | ~x4 | x5 | ~x0 | x2)));
  assign n579 = ((x4 ^ x5) | ((x2 | ~x3 | ~x0 | x1) & (x0 | (x1 ? (~x2 | x3) : (x2 ^ x3))))) & ((x0 ? (x1 | x3) : (~x1 | ~x3)) | (x2 ? (~x4 | x5) : (x4 | ~x5))) & (x0 | ((x1 | ((~x2 | x3 | x4 | ~x5) & (x2 | ~x3 | ~x4 | x5))) & (~x1 | x2 | x3 | ~x4 | x5)));
  assign z041 = (~x1 & (~n581 | (x0 & ~n582))) | ~n589 | (~x0 & ~n583);
  assign n581 = (x2 | ((~x0 | (x3 ? (x5 | ~x6) : (~x4 | x6))) & (x5 | x6 | x3 | ~x4) & (x0 | (x3 ? (x6 | (x4 ^ x5)) : (x5 | ~x6))))) & (x0 | ~x2 | x3 | ~x5 | (~x4 & ~x6));
  assign n582 = (x3 | ((x7 | ((x5 | ~x6 | x2 | x4) & (~x2 | ~x5 | (~x4 ^ x6)))) & (x5 | ~x6 | ~x7 | x2 | ~x4))) & (x2 | ~x3 | ~x5 | x6 | (~x4 ^ ~x7));
  assign n583 = (~n447 | ~n588) & (n585 | ~n587) & (~n584 | n586);
  assign n584 = ~x4 & ~x7;
  assign n585 = x1 ? (x2 | ~x5) : (~x2 | x5);
  assign n586 = (~x2 | x5 | (x1 ? (~x3 | x6) : (x3 | ~x6))) & (x1 | x2 | ~x5 | (x3 ^ x6));
  assign n587 = (~x4 ^ ~x7) & (x3 ^ ~x6);
  assign n588 = ~x3 & ~x1 & ~x2;
  assign n589 = (n590 | n594) & (~n152 | n592) & (n591 | n593);
  assign n590 = x5 ^ x6;
  assign n591 = x4 ? (x5 | ~x6) : (~x5 | x6);
  assign n592 = x2 ? (x4 | (x3 ? (~x5 | ~x6) : (~x5 ^ x6))) : ((~x3 | (x4 ? (~x5 | x6) : x5)) & (x5 | ((x4 | x6) & (x3 | ~x4 | ~x6))));
  assign n593 = (~x2 | x3 | ~x0 | x1) & (x0 | ~x3 | (~x1 ^ ~x2));
  assign n594 = (x1 | ((~x3 | ~x4 | x0 | ~x2) & (~x0 | x2 | (x3 ^ x4)))) & (x0 | ~x1 | ~x2 | x3 | ~x4);
  assign z042 = ~n601 | (~x1 & (n596 | n597 | ~n599));
  assign n596 = n366 & ((~x2 & (x3 ? (x4 & x5) : (~x4 & x6))) | (~x3 & ~x4 & x5 & x6) | (x3 & ~x5 & ~x6 & (x2 | ~x4)));
  assign n597 = ~n598 & (~x3 ^ x6);
  assign n598 = x0 ? (x2 | ((x5 | ~x7) & (~x4 | (x5 & ~x7)))) : (~x2 | x4 | (~x5 & x7));
  assign n599 = (~x0 | x2 | ~x3 | (~n196 & (x4 | n600))) & (x0 | ~x2 | x3 | ~x4 | n600);
  assign n600 = x5 ? (~x6 | ~x7) : (x6 | x7);
  assign n601 = (n420 | n604) & (n293 | n603) & (~n152 | n602);
  assign n602 = (x3 | ((x2 | x5 | (x6 ^ x7)) & (~x5 | ~x7 | (~x2 & (~x4 | ~x6))))) & (~x3 | ((~x6 | ~x7 | x4 | ~x5) & (~x2 | x5 | x6 | (~x4 ^ ~x7)))) & (~x6 | ~x7 | ~x2 | ~x5);
  assign n603 = x0 ? (x1 | ((~x2 | x3 | (~x4 ^ x6)) & (x4 | x6 | x2 | ~x3))) : (((x3 ^ x6) | (~x1 & (x2 | x4))) & (x1 | ~x4 | ((x3 | ~x6) & (x2 | ~x3 | x6))));
  assign n604 = (x1 | (x0 ? (x3 | x4) : (~x4 | (x2 ^ x3)))) & (x0 | x2 | ~x3 | (~x1 & x4));
  assign z043 = n606 | ~n610 | ~n616 | (~x3 & ~n609);
  assign n606 = ~x0 & ((~x1 & ~n607) | (x1 & ~x2 & n139 & ~n608));
  assign n607 = (~x7 | ((x4 | ~x5 | x6 | ~x2 | x3) & ((x3 ? (~x4 | ~x5) : (x4 | x5)) | (~x2 ^ ~x6)))) & (~x5 | x7 | ((~x2 | ~x3 | ~x4 | x6) & (x2 | ~x6 | (~x3 ^ x4))));
  assign n608 = x3 ? (~x6 | x7) : (~x6 ^ ~x7);
  assign n609 = x0 ? (x1 | ((~x2 | ~x4 | x5 | ~x7) & (x2 | ((~x5 | ~x7) & (x4 | x5 | x7))))) : (x1 ? ((~x2 | x5 | ~x7) & (x2 | ~x4 | ~x5 | x7)) : (x2 ? ((x5 | x7) & (~x4 | ~x5 | ~x7)) : (x4 ? (x5 | ~x7) : (~x5 | x7))));
  assign n610 = (n611 | n615) & (n612 | ~n613) & (n293 | n614);
  assign n611 = x3 ? (~x6 | ~x7) : (x6 | x7);
  assign n612 = (~x2 | x3 | ~x4 | x6 | x7) & (x2 | (~x6 ^ x7) | (~x3 ^ x4));
  assign n613 = ~x5 & x0 & ~x1;
  assign n614 = (x0 | ~x1 | x2 | ~x3 | ~x4) & (~x0 | x1 | (x2 ? (x3 | x4) : (~x3 | ~x4)));
  assign n615 = (x0 | ~x1 | ~x2 | x5) & (x2 | ~x5 | ~x0 | x1);
  assign n616 = (x0 | n618) & (~x3 | n617);
  assign n617 = (x4 | ((~x0 | x1 | x2 | ~x5 | x7) & (x0 | ~x7 | ((~x2 | ~x5) & (~x1 | x2 | x5))))) & (x0 | ~x1 | ~x2 | (x5 ^ x7));
  assign n618 = x1 ? (x3 | ((x2 | x5 | x6 | ~x7) & (~x2 | ~x5 | (~x6 ^ x7)))) : (~x3 | x5 | (x2 ? (~x6 | x7) : (x6 ^ x7)));
  assign z044 = n620 | (~n179 & ~n624) | (n152 & ~n625);
  assign n620 = ~x1 & (~n622 | (~x3 & ~n623) | (~x2 & x3 & ~n621));
  assign n621 = (~x0 | ((~x5 | ~x6 | x7) & (x6 | ~x7 | ~x4 | x5))) & (x0 | x4 | x5 | x6 | ~x7) & (~x5 | ((~x4 | ~x6 | x7) & (x0 | x6 | (~x4 ^ ~x7))));
  assign n622 = x3 ? (x0 ? (x2 | ((~x4 | x5 | ~x6) & (x6 | (x4 & ~x5)))) : ((~x2 | ~x5 | (~x4 ^ x6)) & (x5 | x6 | x2 | ~x4))) : (~x6 | (x0 ? (~x2 | x4) : (x2 ? ~x4 : (x4 | ~x5))));
  assign n623 = x0 ? ((x2 | x4 | x5 | ~x6 | ~x7) & (x6 | ((~x2 | (x4 ? (~x5 | x7) : (x5 | ~x7))) & (x2 | ~x4 | x5 | ~x7)))) : ((x4 | ((~x2 | ((~x6 | x7) & (~x5 | x6 | ~x7))) & (x5 | ((~x6 | x7) & (x2 | x6 | ~x7))))) & (x2 | ~x4 | (x5 ? (x6 | x7) : (~x6 | ~x7))));
  assign n624 = (x1 | (x0 ? (x3 | (x5 ? x2 : ~x4)) : (~x3 | x5 | (~x2 & x4)))) & (x0 | ~x1 | x2 | ~x3 | x4 | ~x5);
  assign n625 = (x2 & ((~x5 & x6 & x7) | (~x3 & (x6 | (~x5 & x7))))) | (x6 & ((~x2 & ~x4 & x5) | (~x3 & ~x5 & x7))) | (~x6 & ~x7 & ~x2 & x5) | (x3 & ((~x6 & (x4 | x5 | ~x7)) | (~x2 & (~x6 | (x5 & ~x7)))));
  assign z045 = (~x1 & ~n630) | (~x3 & ~n627) | n631 | (x3 & ~n632);
  assign n627 = (x1 | n628) & (x0 | ~x1 | n629);
  assign n628 = (x5 | ((~x0 | ~x7 | (x2 ? (x4 | ~x6) : x6)) & (x7 | ((x2 | x4 | ~x6) & (x0 | (~x2 ^ x6)))))) & (~x4 | ~x5 | ((x6 | (x0 ? (~x2 | x7) : (~x2 ^ ~x7))) & (x0 | x2 | ~x6 | ~x7)));
  assign n629 = ((~x2 ^ ~x7) | ((x5 | ~x6) & (x4 | ~x5 | x6))) & (x6 | x7 | ~x2 | x5) & (x2 | ~x7 | ((~x5 | ~x6) & (~x4 | x5 | x6)));
  assign n630 = x0 ? ((x2 | ~x3 | x5 | (~x4 ^ x7)) & (x3 | (x2 ? ((x4 | ~x5 | ~x7) & (x5 | x7)) : (~x5 | x7)))) : (x5 ? (x2 ? (x3 ? (~x4 | ~x7) : (x4 | x7)) : (x3 ? (~x4 | x7) : (x4 | ~x7))) : ((x2 | ~x3 | ~x4 | ~x7) & (~x2 | (~x3 ^ x7))));
  assign n631 = n152 & ((x5 & (x2 ? (x7 & (x3 | x4)) : (~x7 & (x3 ^ x4)))) | (x3 & ~x5 & (x2 ? (~x4 & ~x7) : x7)));
  assign n632 = (~x5 | (n634 & (x6 | n635))) & (n633 | ~n636) & (x5 | ~x6 | n635);
  assign n633 = x1 ? (~x2 | ~x4) : (x2 | x4);
  assign n634 = (~x0 | x1 | x2 | ~x6 | x7) & (x0 | ((~x1 | x7 | (x2 ? (x4 | x6) : (~x4 | ~x6))) & (x4 | ~x7 | ((x2 | ~x6) & (x1 | ~x2 | x6)))));
  assign n635 = (~x0 | x1 | x2 | ~x4 | ~x7) & (x0 | x7 | (x1 ? (~x2 | ~x4) : (x2 | x4)));
  assign n636 = x7 & ~x6 & ~x0 & ~x5;
  assign z046 = ~n640 | (x6 ? ~n638 : ~n639);
  assign n638 = (x2 | ((x4 | ~x5 | x0 | ~x3) & (x1 | (x0 ? (x3 ? ~x5 : (x4 | x5)) : (x3 ? x4 : (~x4 | ~x5)))))) & (x0 | ((~x1 | ((x3 | x5) & (~x4 | ~x5 | ~x2 | ~x3))) & (~x2 | x3 | ~x4 | x5)));
  assign n639 = (x1 | ((~x0 | x5 | ((x3 | ~x4) & (x2 | ~x3 | x4))) & (~x2 | ((x0 | ~x3 | ~x4) & (x3 | x4 | ~x5))) & (x0 | ~x5 | (x3 ^ x4)))) & (x0 | ~x1 | ~x3 | ((x4 | x5) & (x2 | (x4 & x5))));
  assign n640 = (x1 | (x6 ? n642 : n641)) & (x0 | ~x1 | n643);
  assign n641 = (x2 | ((~x0 | ~x5 | (x3 ? (x4 | ~x7) : x7)) & (x5 | x7 | x0 | ~x3))) & (x0 | x5 | (x3 ? (x4 | x7) : (~x7 | (~x2 & ~x4))));
  assign n642 = (x5 | ((~x0 | (x2 ? (x3 | (~x4 ^ x7)) : ((~x4 | ~x7) & (~x3 | x4 | x7)))) & (x0 | x2 | x3 | ~x4 | x7))) & (x0 | ~x2 | ((x3 | x4 | x7) & (~x5 | (x3 ? (~x4 ^ x7) : (~x4 | ~x7)))));
  assign n643 = x5 ? (x6 ? (((x2 ^ ~x4) | (x3 ^ ~x7)) & (x2 | x3 | x4 | x7)) : ((~x3 | ~x4 | ~x7) & (~x2 | (~x3 ^ ~x7)))) : ((x2 | x3 | x4 | x6 | ~x7) & (~x2 | ~x3 | ~x4 | ~x6 | x7));
  assign z047 = n645 | n649 | ~n653 | (~n293 & ~n648);
  assign n645 = x6 & ((~x3 & ~n646) | (n147 & ~n647));
  assign n646 = (x1 | ((~x4 | ((x5 | x7 | x0 | ~x2) & (~x0 | (x2 ? (x5 | ~x7) : (~x5 | x7))))) & (x0 | ~x5 | (x2 ? ~x7 : (x4 | x7))))) & (x0 | ((~x5 | ~x7 | ~x2 | x4) & (~x1 | ((x4 | x5 | x7) & (x2 | (x5 ^ x7))))));
  assign n647 = ((~x1 ^ x2) | (x5 ^ x7)) & (~x2 | ~x7 | ((x4 | ~x5) & (~x1 | ~x4 | x5)));
  assign n648 = (x1 | (x0 ? (~x6 | (x2 ? (x3 | x4) : ~x3)) : ((x3 | x6) & (x2 | (x6 & (x3 | ~x4)))))) & (x0 | x2 | x3 | x4 | x6);
  assign n649 = ~x6 & ((n650 & ~n652) | (~n217 & ~n651));
  assign n650 = ~x5 & ~x1 & x3;
  assign n651 = x0 ? (x1 | x2 | (x3 & x4)) : (~x1 | (~x2 & (~x3 | ~x4)));
  assign n652 = (x0 | ~x2 | x4 | ~x7) & (~x4 | x7 | ~x0 | x2);
  assign n653 = ~n657 & (~n152 | n656 | (~n654 & ~n655));
  assign n654 = x3 & ~x4;
  assign n655 = ~x3 & x4;
  assign n656 = x2 ? (x5 | ~x6) : (~x5 | x6);
  assign n657 = ~x1 & (x2 ^ x6) & (x0 ? (~x3 & ~x5) : (x3 & x5));
  assign z048 = n659 | n663 | ~n664 | ~n667 | (~n179 & ~n662);
  assign n659 = ~x0 & ((~x4 & ~n660) | (n142 & n260 & ~n661));
  assign n660 = x1 ? ((~x2 | ~x3 | ~x5 | ~x6 | ~x7) & (x2 | x3 | x5 | x6 | x7)) : ((~x5 | ((~x2 | x3 | x6 | x7) & (x2 | ~x7 | (~x3 ^ x6)))) & (~x2 | x5 | (x3 ? x6 : (~x6 | x7))));
  assign n661 = x1 ? (~x6 ^ x7) : (x6 | x7);
  assign n662 = (x1 | ((~x3 | ~x4 | ~x5 | ~x0 | x2) & (~x2 | (x0 ? (x3 | (x4 & x5)) : (~x3 | (~x4 ^ x5)))))) & (x0 | ~x1 | x2 | (x4 ? x3 : (~x3 & ~x5)));
  assign n663 = ~x0 & ((~x1 & x2 & ~x3 & x4 & ~x6) | (x6 & ((~x1 & ~x2 & ~x3 & x4) | (x1 & (x2 ? (~x3 & ~x4) : (x3 & x4))))));
  assign n664 = ~n665 & (~n153 | ~n655 | ~n265) & (~n233 | n666);
  assign n665 = ~x6 & ~x4 & x3 & ~x2 & x0 & ~x1;
  assign n666 = (x1 | ((x6 | ~x7 | ~x2 | x3) & (x2 | ~x3 | ~x6 | x7))) & (~x1 | x2 | x3 | x6 | ~x7);
  assign n667 = (n164 | n668) & (~x4 | ~n207 | n669);
  assign n668 = (x1 | x2 | x3 | x4) & (x0 | ((x1 | x2 | ~x3 | ~x4) & (~x1 | ~x2 | (~x3 ^ x4))));
  assign n669 = (x3 | ~x5 | x6 | x7) & (x2 | x5 | (x3 ? x6 : (~x6 | x7)));
  assign z049 = n671 | n676 | ~n677 | (x3 ? ~n675 : ~n674);
  assign n671 = ~x1 & ((n147 & ~n673) | (~x3 & ~n672));
  assign n672 = x0 ? (~x4 | ((~x6 | ~x7 | x2 | x5) & (x6 | x7 | ~x2 | ~x5))) : (x4 | ~x6 | (x2 ? (x5 | ~x7) : (x5 ^ x7)));
  assign n673 = x2 ? (~x4 | ~x5 | (x6 ^ x7)) : (x4 | x5 | (~x6 ^ x7));
  assign n674 = (x1 | (x0 ? (~x4 | ((x5 | x7) & (x2 | ~x5 | ~x7))) : (x4 | (x2 ? (x5 ^ x7) : (~x5 | x7))))) & (x0 | ~x1 | x2 | x4 | x5 | ~x7);
  assign n675 = (~x4 | ((x0 | x1 | ~x2 | x5 | x7) & ((~x5 ^ x7) | (x0 ? (x1 | x2) : (~x1 | ~x2))))) & (x0 | x4 | ((x5 | x7 | ~x1 | ~x2) & (x1 | ((~x5 | x7) & (~x2 | x5 | ~x7)))));
  assign n676 = n139 & n152 & ((~x2 & ~x3 & (x6 ^ x7)) | (x3 & ((x6 & x7) | (x2 & ~x6 & ~x7))));
  assign n677 = ((x0 ? (x1 | x4) : (~x1 | ~x4)) | ((x3 | x7) & (x2 | ~x3 | ~x7))) & (x0 | (x1 ? (x4 | (x2 ? (x3 | ~x7) : (~x3 | x7))) : (~x4 | ((x3 | ~x7) & (x2 | ~x3 | x7)))));
  assign z050 = ~n683 | (~x0 & (~n681 | n682 | (n679 & n680)));
  assign n679 = ~x3 & ~x1 & x2;
  assign n680 = x7 & x6 & ~x4 & ~x5;
  assign n681 = (x6 | ((~x1 | ~x2 | ~x3 | ~x4) & (x1 | ((x2 | ~x4) & (x4 | ~x5 | ~x2 | x3))))) & (x4 | ((x2 | ~x3) & (~x1 | (x2 & (~x3 | ~x5 | ~x6))))) & (~x4 | ((~x5 | ~x6 | ~x2 | ~x3) & (x2 | (x3 & x5))));
  assign n682 = n408 & ((~x1 & x6 & (x3 ? (x4 & ~x7) : (~x4 & x7))) | (x1 & x3 & x4 & ~x6 & ~x7));
  assign n683 = x2 | ~n207 | (x3 & (x4 | (x5 & ~n140)));
  assign z051 = n685 | n689 | n690 | ~n691 | (~x0 & ~n688);
  assign n685 = x5 & ((~x1 & ~n687) | (x4 & n152 & n686));
  assign n686 = ~x6 & (x2 ? (~x3 & ~x7) : (x3 & x7));
  assign n687 = (x2 | ((x4 | ((~x0 | x6 | (~x3 ^ ~x7)) & (~x6 | ~x7 | x0 | x3))) & (~x4 | ~x6 | ~x7 | x0 | ~x3))) & (x0 | ~x2 | x7 | (x3 ? (x4 | x6) : (~x4 | ~x6)));
  assign n688 = x1 ? ((~x4 | x5 | x6 | ~x2 | ~x3) & (~x5 | (~x3 ^ ~x6) | (x2 ^ ~x4))) : ((x4 | (x2 ? (x3 | (x5 ^ x6)) : (~x3 | (~x5 ^ x6)))) & (~x2 | ~x4 | ~x5 | (~x3 ^ ~x6)));
  assign n689 = x2 & ((x0 & ~x1 & ~x3 & ~x4 & ~x5) | (~x0 & ((~x3 & x4 & ~x5) | (x1 & (x3 ? (x4 & x5) : ~x5)))));
  assign n690 = ~x2 & ((~x1 & (x0 ? (x3 ? x4 : (~x4 & ~x5)) : (~x3 & x4))) | (~x0 & ~x3 & (x4 ? ~x5 : x1)));
  assign n691 = ~x6 | (x5 ? (~n153 | ~n654) : (~n692 | n693));
  assign n692 = ~x1 & ~x3;
  assign n693 = (x0 | ~x2 | x4 | x7) & (~x4 | ~x7 | ~x0 | x2);
  assign z052 = ~n697 | (~x1 & (x2 ? ~n696 : ~n695));
  assign n695 = ((~x3 ^ ~x4) | ((x6 | x7 | ~x0 | x5) & (~x6 | ~x7 | x0 | ~x5))) & (~x0 | x4 | ~x5 | x6 | ~x7) & (x0 | x5 | ((~x4 | ~x6 | x7) & (x3 | x4 | x6 | ~x7)));
  assign n696 = (x3 | ~x4 | ((x6 | x7 | ~x0 | x5) & (~x6 | ~x7 | x0 | ~x5))) & (x0 | x4 | ((x5 | ~x6 | x7) & (x6 | ~x7 | ~x3 | ~x5)));
  assign n697 = (~n154 | n700) & (~n152 | n698) & (~x5 | n699);
  assign n698 = (x6 | (x2 ? ((x3 | ~x4 | ~x5 | ~x7) & (~x3 | x4 | x5 | x7)) : (~x4 | ((~x3 | ~x5 | ~x7) & (x5 | x7))))) & (x2 | x4 | ~x6 | (x3 ? (~x5 | ~x7) : (x5 | x7)));
  assign n699 = (x1 | ((~x0 | x2 | ~x4) & (x4 | ((x2 | ~x3 | ~x6) & (x3 | ((~x2 | ~x6) & (~x0 | (~x2 & ~x6)))))))) & (x0 | ((~x2 | ~x3 | (~x6 & (~x1 | ~x4))) & (~x1 | ~x6 | (x3 & ~x4))));
  assign n700 = (x2 & (x0 | (x1 & x3 & ~x4))) | (x0 & (x3 | ~x4)) | (~x1 & ~x2 & ~x3 & ~x4) | (x1 & x4 & (~x2 | ~x3));
  assign z053 = n702 | n706 | n707 | n709 | (~x3 & ~n705);
  assign n702 = ~x2 & ((~x1 & ~n703) | (n152 & ~n704));
  assign n703 = x6 ? ((x3 | ((x4 | ~x5 | ~x7) & (x5 | x7 | ~x0 | ~x4))) & (~x7 | ((~x3 | ~x4 | x5) & (x0 | ((~x4 | x5) & (~x3 | (~x4 & x5))))))) : (x7 | ((x0 | ~x4 | x5) & (~x3 | (x4 ^ x5))));
  assign n704 = (~x6 | ~x7 | (x3 ? (~x4 | ~x5) : x5)) & (x4 | x7 | ((~x5 | x6) & (x3 | (~x5 & x6))));
  assign n705 = (x0 | ((~x4 | x5 | x6 | ~x1 | ~x2) & (~x6 | ((~x1 | (x2 ? x4 : (~x4 | ~x5))) & (~x2 | x4 | ~x5) & (x1 | x5 | (x2 ^ x4)))))) & (x1 | x6 | (x2 ? (x4 | x5) : (~x4 | ~x5)));
  assign n706 = n147 & ((x6 & ((~x1 & x2 & x4) | (~x4 & (x1 ? (x2 ^ ~x5) : (~x2 & x5))))) | (x1 & x2 & x4 & x5 & ~x6));
  assign n707 = ~n164 & ~n708;
  assign n708 = (x1 | ((~x2 | ((x4 | ~x5 | x0 | ~x3) & (~x4 | x5 | ~x0 | x3))) & (x2 | ((~x3 | x4 | x5) & (~x0 | (x4 & (~x3 | x5))))) & (x4 | ~x5 | ~x0 | x3))) & (x0 | ~x1 | (x2 ? (x3 ? (x4 | x5) : (~x4 | ~x5)) : (~x4 | (~x3 & x5))));
  assign n709 = x2 & ((n139 & n140 & n319) | (~x0 & ~n710));
  assign n710 = (~x3 | x4 | x5 | ((~x6 | ~x7) & (x1 | x6 | x7))) & (x1 | x3 | ~x4 | ~x5 | (x6 ^ x7));
  assign z054 = n712 | n716 | n719 | ~n721 | (~x4 & ~n718);
  assign n712 = x7 & ((~x4 & ~n713) | n715 | (~n369 & ~n714));
  assign n713 = (x3 | ~x5 | ~x6 | x0 | ~x1 | ~x2) & (x5 | ((~x0 | x1 | x2 | ~x3 | ~x6) & (x0 | ((~x1 | ~x3 | (~x2 ^ x6)) & (x1 | ~x2 | x3 | ~x6)))));
  assign n714 = (~x0 | x1 | x3 | x4 | ~x5) & (x0 | ~x1 | ~x4 | (x3 ^ x5));
  assign n715 = ~x6 & x4 & x3 & ~x2 & x0 & ~x1;
  assign n716 = ~n717 & ~x1 & ~x7;
  assign n717 = (x2 | ((x4 | (x0 ? (x3 ? (x5 | x6) : (~x5 | ~x6)) : (x3 | (~x5 ^ x6)))) & (~x4 | ~x6 | ~x0 | ~x3))) & (~x0 | ~x2 | x3 | x4 | ~x5 | x6);
  assign n718 = (x2 | ~x7 | ((x0 | ~x1 | ~x3 | ~x5) & (x1 | (x0 ? (x3 ^ x5) : (x3 | ~x5))))) & (x0 | ~x2 | x7 | ((x3 | x5) & (~x1 | ~x3 | ~x5)));
  assign n719 = ~n720 & ((~x0 & (x2 ? (~x3 & x5) : (x3 & ~x5))) | (~x1 & ((~x0 & ~x2 & x3) | (~x3 & ~x5 & x0 & x2))));
  assign n720 = x4 ^ x7;
  assign n721 = ~n723 & ~n724 & (~x4 | ~n722 | n725);
  assign n722 = ~x0 & ~x3;
  assign n723 = ~x0 & ((x2 & x3 & ((x4 & ~x7) | (~x1 & ~x4 & x7))) | (x1 & ~x2 & ~x3 & ~x4 & x7));
  assign n724 = ~x7 & x4 & ~x3 & ~x2 & x0 & ~x1;
  assign n725 = x2 ? (x5 | x7) : ((~x5 | x7) & (x1 | x5 | ~x7));
  assign z055 = ~n737 | n735 | n734 | n732 | n727 | n730;
  assign n727 = ~x3 & ((n233 & ~n729) | (x4 & ~n728));
  assign n728 = (x1 | ((x0 | x2 | x5 | x6 | ~x7) & (~x0 | x7 | (x2 ? (~x5 | x6) : (x5 | ~x6))))) & (x0 | ~x1 | ~x6 | (x5 ^ x7));
  assign n729 = (~x6 | ((~x2 | x5 | ~x7) & (~x1 | ((x5 | ~x7) & (~x2 | ~x5 | x7))))) & (x1 | x2 | x6 | (~x5 ^ x7));
  assign n730 = ~x1 & ~n731;
  assign n731 = (x5 | (x0 ? ((~x2 | x3 | ~x6) & (x2 | ~x3 | ~x4 | x6)) : (x3 | (x2 ? (~x4 | x6) : (x4 | ~x6))))) & (x2 | ~x3 | ~x5 | ~x6 | (~x0 ^ x4));
  assign n732 = ~n733 & ((x0 & ~x1 & ~x2 & ~x3 & x6) | (x3 & ((~x0 & (~x6 | (~x1 & x2))) | (~x1 & ~x2 & ~x6))));
  assign n733 = x4 ^ x5;
  assign n734 = ~x0 & ((~x4 & x5 & ~x1 & x3) | (~x3 & ((~x5 & x6 & ~x1 & x4) | (x1 & ~x6 & (x4 ^ x5)))));
  assign n735 = x3 & x6 & n152 & ~n736;
  assign n736 = x4 ? (~x5 ^ x7) : ((x5 | x7) & (~x2 | ~x5 | ~x7));
  assign n737 = x6 | ((x4 | ~x5 | ~n319) & (~x3 | ~x4 | x5 | ~n738));
  assign n738 = x2 & ~x0 & x1;
  assign z056 = (~x0 & (~n744 | (x3 & ~n743))) | n745 | (~x3 & ~n740);
  assign n740 = (x6 | n741) & (x0 | ~x6 | n742);
  assign n741 = (x1 | (x0 ? ((x2 | x4 | x5 | ~x7) & (~x2 | ~x4 | ~x5 | x7)) : (x2 | x7 | (~x4 ^ x5)))) & (x0 | ~x1 | ~x7 | (~x2 & x4 & ~x5));
  assign n742 = (~x1 | x7 | (~x2 & ~x4 & x5)) & (x1 | x2 | x4 | ~x7);
  assign n743 = (~x7 | ((x2 | ((~x1 | x6) & (x5 | ~x6 | x1 | x4))) & (~x1 | x6 | (x4 & ~x5)))) & (~x1 | ~x6 | x7);
  assign n744 = x1 ? ((~x4 | x5 | x6 | ~x2 | ~x3) & (x2 | x3 | x4 | ~x5 | ~x6)) : (~x6 | (~x2 & ~x4 & (~x3 | ~x5)));
  assign n745 = (~x2 | (~x3 & (~x4 | ~x5))) & n226 & (x2 | x3 | x4 | x5);
  assign z057 = ~n751 | (~x0 & (~n747 | (x5 & ~n750)));
  assign n747 = (x5 | n748) & (~x5 | n749 | ~x1 | x4);
  assign n748 = (~x4 | ((x2 | x3 | (x1 ? (x6 | ~x7) : (x6 ^ x7))) & (~x1 | ~x2 | ~x3 | (~x6 ^ x7)))) & (x2 | ((x1 | x4 | ((~x6 | x7) & (~x3 | x6 | ~x7))) & (~x6 | x7 | ~x1 | x3)));
  assign n749 = (~x2 | ~x3 | ~x6 | ~x7) & (x2 | x3 | (x6 ^ x7));
  assign n750 = (~x4 | ((x1 | x2 | x3 | ~x7) & (~x1 | x7 | (~x2 ^ ~x3)))) & (x1 | x2 | x4 | (x3 ^ x7));
  assign n751 = n754 & (~n261 | ~n448) & (~n190 | (~n752 & ~n753));
  assign n752 = x7 & ~x3 & ~x4;
  assign n753 = x7 & ~x5 & ~x3 & x4;
  assign n754 = (x0 | ((~x2 | (x1 ? (x3 | x7) : ~x7)) & (~x1 | ~x3 | x7 | (x2 & x4)))) & (x1 | x2 | ~x7 | (~x0 & (~x3 | ~x4)));
  assign z058 = n757 | n758 | (~x0 & ~n756) | ~n761;
  assign n756 = (~x1 | ((~x6 | ((x2 | x3 | x4 | ~x5) & (~x2 | x5 | (x3 & ~x4)))) & (~x2 | ~x3 | x4 | ~x5 | x6))) & (x5 | ((x2 | ((x3 | ~x4 | x6) & (x1 | x4 | ~x6))) & (~x2 | x3 | ~x4 | ~x6)));
  assign n757 = ~x1 & (x2 ? (x0 ? (~x3 & (x4 ^ x5)) : (x3 | (x4 & x5))) : ((~x0 & ~x3 & ~x4 & x5) | (x4 & ~x5 & x0 & x3)));
  assign n758 = ~x4 & ((x6 & ~n759) | (~x3 & ~x5 & ~x6 & ~n760));
  assign n759 = (~x3 | ~x5 | ~x7 | ~x0 | x1 | x2) & (x0 | ~x2 | x7 | (x1 ? (~x3 | ~x5) : (x3 | x5)));
  assign n760 = (x0 & (x1 | (~x2 & x7))) | (x1 & ~x2 & x7) | (~x7 & (x2 | (~x0 & ~x1)));
  assign n761 = ~n764 & (~n196 | ~n763) & (~n186 | ~n762 | ~n190);
  assign n762 = ~x5 & x6;
  assign n763 = ~x3 & x2 & x0 & ~x1;
  assign n764 = ~x0 & x1 & x2 & ((x3 & ~x4 & ~x5) | (x5 & (~x3 | x4)));
  assign z059 = x3 ? (n770 | ~n772) : ~n766;
  assign n766 = n769 & (x1 | n767) & (x0 | ~x1 | x4 | n768);
  assign n767 = (~x5 | ~x6 | ~x7 | ~x0 | x4) & (x7 | ((~x0 | x2 | ~x4 | x5 | ~x6) & (x6 | ((~x2 | x4 | x5) & (~x0 | ((x4 | x5) & (~x2 | ~x4 | ~x5)))))));
  assign n768 = (x5 | x6 | x7) & (~x2 | ~x5 | ~x6 | ~x7);
  assign n769 = (x0 | (x4 ? (x5 | x6) : (~x5 | (x1 & (x2 | ~x6))))) & (x1 | ~x4 | x5 | (x6 & (~x0 | ~x2)));
  assign n770 = ~x4 & (x5 ? (n264 & ~n771) : (n265 & (n141 | ~n771)));
  assign n771 = x0 ? (x1 | x2) : ~x1;
  assign n772 = (~x4 & ((x5 & x6) | (~x0 & ~x1 & ~x6))) | (~x5 & (~x6 | (x0 & x4))) | (x0 & (x1 | x2));
  assign z060 = n774 | n777 | n779 | ~n781 | (~n590 & ~n776);
  assign n774 = x5 & ((n140 & n655 & n190) | (x7 & ~n775));
  assign n775 = (x0 | ((x2 | ((~x3 | x4 | ~x6) & (~x1 | (x6 ? x4 : x3)))) & (~x4 | x6) & (x1 | ~x2 | x4 | ~x6))) & (x1 | x2 | x6 | (~x4 & (~x0 | x3)));
  assign n776 = (x1 | (x0 ? (x4 | x7 | (x2 & x3)) : (x2 ? (~x3 | ~x4) : (x3 | ~x7)))) & (x0 | ((~x4 | ~x7 | x2 | x3) & (~x1 | x4 | x7 | (~x2 & ~x3))));
  assign n777 = ~n778 & (x3 ? ~x2 : (x2 | ~x7));
  assign n778 = x0 ? (x1 | (x4 ? (x5 | ~x6) : (~x5 | x6))) : ((~x4 | (x5 ^ x6)) & (~x1 | x4 | ~x5 | x6));
  assign n779 = ~n780 & ~x5 & n233;
  assign n780 = (~x1 | x2 | x3 | x6 | x7) & (x1 | ((~x3 | x6 | x7) & (~x2 | ((x6 | x7) & (x3 | ~x6 | ~x7)))));
  assign n781 = (~x6 | n782) & (~n654 | ~n738 | ~x5 | x6);
  assign n782 = (x0 | ((~x1 | ~x2 | ~x3 | ~x4 | ~x5) & (x1 | x2 | x4 | x5))) & (~x0 | x1 | x2 | ~x4 | ~x5);
  assign z061 = n785 | ~n787 | (n784 & ~n786);
  assign n784 = ~x1 & ~x4;
  assign n785 = ~x7 & n154 & ((~x1 & ~x2 & (x0 ^ x4)) | (~x0 & ~x4 & (x1 | x2)));
  assign n786 = (x0 | x2 | ~x3 | x5 | x6 | x7) & (~x0 | ~x2 | x3 | (x5 ? (x6 | ~x7) : x7));
  assign n787 = ((~x5 | ~x7) & (x4 ^ ~x6)) | (~x5 & ~x7 & (~x6 | n788)) | (n788 & (~n763 | (x5 & x7))) | (x5 & x7 & (~x4 ^ ~x6));
  assign n788 = x0 & (x1 | x2);
  assign z062 = ~n792 | (n692 & ~n791) | (~x7 & n784 & ~n790);
  assign n790 = (~x0 | ~x2 | x3 | ~x5 | ~x6) & (x0 | x6 | (x2 ? (x3 | ~x5) : ~x3));
  assign n791 = (x0 | x2 | ~x5 | x6 | x7) & (~x0 | ~x2 | x5 | (x6 & ~x7));
  assign n792 = (x0 & (x1 | x2)) | (x5 & (~x6 | x7)) | (~x7 & ((~x5 & x6) | (~x0 & ~x1 & ~x2 & ~x6)));
  assign z063 = (~n179 & ~n794) | (~x1 & (n796 | (~x3 & ~n795)));
  assign n794 = x0 ? (x1 | (x2 & (x3 | (x4 & x5)))) : (~x1 & ((~x2 & (x4 ^ x5)) | (~x3 & (~x2 | (~x4 & x5)))));
  assign n795 = (x0 | ~x6 | ((x2 | (x5 & ~x7)) & (x4 | (x2 & (~x5 | ~x7))))) & (~x5 | x6 | x7 | ~x0 | ~x2 | ~x4);
  assign n796 = x3 & x6 & n303 & (~x4 ^ (~x5 & x7));
  assign z064 = ~n801 | (~x1 & (~n798 | ~n799));
  assign n798 = (x0 | x2 | x3 | x5 | ~x7) & (x7 | ((~x2 | ((~x0 | x3 | (x4 & x5)) & (x4 | ~x5 | x0 | ~x3))) & (x0 | x2 | ~x3 | ~x4 | ~x5)));
  assign n799 = (~x7 | ~n233 | n527 | ~n762) & (x7 | n800);
  assign n800 = (x3 | ~x5 | ((~x0 | ~x2 | ~x4 | x6) & (x0 | ~x6 | (x2 ^ ~x4)))) & (x0 | x2 | ~x3 | x5 | (x4 ^ x6));
  assign n801 = (x1 | x2 | ((~x0 | x7) & (x0 | x4 | ~x5 | ~x7))) & (x0 | x7 | (~x1 & (~x2 | (~x4 & x5))));
  assign z065 = ~x0 & (~n804 | (~x3 & ~n803));
  assign n803 = (~x2 | x4 | x5 | ~x6 | x7) & (~x5 | ((~x1 | ~x2 | ~x4 | ~x6 | x7) & (x1 | x6 | ~x7 | (~x2 ^ x4))));
  assign n804 = ~n805 & ~n806 & n807 & (x1 | ~n247 | ~n241);
  assign n805 = ~x5 & ((x1 & x2 & (x3 ? (x4 & x6) : ~x6)) | (~x1 & ~x2 & x3 & ~x4 & ~x6));
  assign n806 = (x1 | x2 | (x3 & x4)) & (~x5 | ~x6) & (x5 | x6) & (~x2 | (x3 ? ~x1 : x4));
  assign n807 = (~x1 & ~x2 & (~x4 | ~x6)) | (x1 & x2) | (~x5 & x6) | (x5 & ~x6);
  assign z066 = n810 | n813 | (~x0 & ~n809) | ~n814;
  assign n809 = (x2 | ((x3 | ((~x5 | ~x6 | x1 | ~x4) & (~x1 | (x4 ? (x5 | x6) : (~x5 | ~x6))))) & (x1 | ~x3 | ~x4 | x5 | ~x6))) & (x4 | x5 | x6 | x1 | ~x3) & (~x2 | ((x6 | ((~x4 | x5 | ~x1 | ~x3) & (x1 | ((x4 | x5) & (~x3 | ~x4 | ~x5))))) & (x4 | ~x5 | ~x6 | x1 | x3)));
  assign n810 = ~x3 & ((~x1 & ~n811) | (x7 & ~n733 & n812));
  assign n811 = (x5 | ((x0 | ~x2 | x4 | ~x6 | x7) & (~x0 | ((x2 | ~x4 | ~x6 | ~x7) & (~x2 | x4 | x6 | x7))))) & (x0 | ~x5 | x6 | ~x7 | (~x2 ^ x4));
  assign n812 = x6 & x2 & ~x0 & x1;
  assign n813 = x5 & ((~x0 & x2 & (x1 ? (~x3 ^ x4) : (x3 & ~x4))) | (~x1 & ~x2 & x4 & (x0 | x3)));
  assign n814 = ~n816 & n815 & (~n177 | n817 | ~x3 | x6);
  assign n815 = (~x0 | x1 | x2 | x3 | x4) & (x0 | ~x2 | (x1 ? (~x3 | x4) : (x3 | ~x4)));
  assign n816 = ~x1 & x3 & ~x5 & (x0 ? (~x2 & ~x4) : (x2 & x4));
  assign n817 = (x0 | ~x4 | x5 | ~x7) & (~x5 | x7 | ~x0 | x4);
  assign z067 = ~n824 | (~x1 & (~n820 | ~n823 | (~x2 & ~n819)));
  assign n819 = (~x3 | ((x0 | x4 | x5 | ~x6 | x7) & (~x0 | ((x4 | ~x5 | x6 | ~x7) & (~x4 | x5 | ~x6 | x7))))) & (x0 | x3 | x6 | ~x7 | (x4 ^ x5));
  assign n820 = (x5 | x6 | ~x7 | n821) & (~x5 | ((~x6 | x7 | n821) & (x4 | x6 | ~x7 | ~n822)));
  assign n821 = (~x0 | ~x2 | x3 | x4) & (x0 | x2 | ~x3 | ~x4);
  assign n822 = ~x3 & ~x0 & x2;
  assign n823 = (x2 | (x0 ? ((~x5 | ~x6 | ~x3 | x4) & (x5 | x6 | (x3 & ~x4))) : ((~x5 | ~x6 | x3 | ~x4) & (x5 | x6 | ~x3 | x4)))) & (x0 | ~x2 | ((x3 | ~x4 | x5) & (~x5 | ~x6 | (~x3 & x4))));
  assign n824 = (n198 | n825) & (~n152 | (n826 & n827));
  assign n825 = (x1 | ((~x3 | ~x4 | x0 | x2) & (x3 | (x0 ? (~x2 ^ x4) : (x2 | x4))))) & (x0 | ((~x2 | ~x3 | x4) & (x3 | ~x4 | ~x1 | x2)));
  assign n826 = x2 ? (x3 ? (x4 ? ~x5 : (x5 | x6)) : (x4 | ~x5)) : (x3 ? (~x4 | x5) : (x4 ? (~x5 | ~x6) : x5));
  assign n827 = ((x5 ? (~x6 | ~x7) : (x6 | x7)) | (x2 ? (x3 | ~x4) : (~x3 | x4))) & (x5 | ~x6 | ~x7 | ~x2 | x3 | x4) & (~x5 | x6 | x7 | x2 | ~x3 | ~x4);
  assign z068 = ~n834 | (~n590 & ~n833) | (~x0 & (~n829 | ~n830));
  assign n829 = x1 ? (x5 ? ((x3 | x4 | x6) & (x2 | (x3 ? (~x4 | ~x6) : x6))) : ((x3 | ~x4 | ~x6) & (~x2 | ~x3 | x4 | x6))) : (x2 ? ((x5 | x6 | x3 | x4) & (~x5 | ~x6 | ~x3 | ~x4)) : (x3 ? (x4 ? (x5 | ~x6) : (~x5 | x6)) : ((~x5 | ~x6) & (~x4 | x5 | x6))));
  assign n830 = x4 ? n832 : n831;
  assign n831 = (~x2 | (~x3 ^ x7) | (x1 ? (x5 | ~x6) : (~x5 | x6))) & (x1 | x2 | x5 | (x3 ? (~x6 | ~x7) : (~x6 ^ x7)));
  assign n832 = (x1 | ((x2 | x3 | ~x5 | x6 | ~x7) & (~x2 | ~x6 | x7 | (~x3 ^ x5)))) & (~x1 | x2 | ~x3 | ~x5 | x6 | ~x7);
  assign n833 = (~x7 | ((~x0 | x1 | ~x2 | x3 | x4) & (x0 | ((x1 | x2 | ~x3 | ~x4) & (~x1 | (x2 ? (x3 | ~x4) : (~x3 | x4))))))) & (x0 | ~x1 | x7 | (x2 ? (~x3 | ~x4) : (x3 | x4)));
  assign n834 = (~n184 | n837) & (~n153 | ~n835) & (n215 | n836);
  assign n835 = x6 & x5 & ~x3 & x4;
  assign n836 = (x0 | ~x1 | ~x3 | (x2 ^ x5)) & (x1 | (x0 ? ((x3 | x5) & (x2 | ~x3 | ~x5)) : (~x2 | (~x3 ^ x5))));
  assign n837 = (~x3 | x4 | x5 | x6 | x7) & ((~x3 ^ ~x7) | (x4 ? (x5 | ~x6) : (~x5 | x6)));
  assign z069 = ~n844 | (~n179 & ~n843) | (~x3 & ~n839);
  assign n839 = n842 & (x0 | n840) & (~x7 | n841 | ~x0 | x1);
  assign n840 = (x4 | ~x6 | ((x7 | (x1 ? (~x2 ^ ~x5) : (x2 ^ ~x5))) & (x1 | x2 | x5 | ~x7))) & (x1 | ~x4 | x6 | (x2 ? x5 : (~x5 | ~x7)));
  assign n841 = (~x5 | x6 | ~x2 | x4) & (x2 | x5 | (x4 ^ ~x6));
  assign n842 = (x0 | ~x1 | ~x2 | ~x4 | x6 | ~x7) & (x4 | ~x6 | x7 | ~x0 | x1 | x2);
  assign n843 = x0 ? (x1 | ((~x2 | x3 | x4 | ~x5) & (~x4 | ((x3 | x5) & (x2 | (x3 & x5)))))) : (x4 ? ((x1 | ~x3 | (~x2 & ~x5)) & (~x2 | ~x5) & (~x1 | x2 | x3 | x5)) : (((~x2 ^ x5) | (~x1 & x3)) & (~x1 | x3 | ~x5) & (x1 | x2 | ~x3 | x5)));
  assign n844 = (n164 | n847) & (~n147 | n845) & (n437 | n846);
  assign n845 = (~x2 | ((x1 | x4 | x5 | ~x6 | x7) & (~x1 | ((~x4 | x5 | x6 | ~x7) & (x4 | ~x5 | ~x6 | x7))))) & (x1 | x2 | ~x5 | (x4 ? (x6 | ~x7) : (~x6 | x7)));
  assign n846 = (x1 | ((~x3 | ~x5 | x0 | ~x2) & (~x0 | (x2 ? (x3 | x5) : ~x5)))) & (x0 | ((x2 | x3 | x5) & (~x1 | ((x3 | x5) & (x2 | (x3 & x5))))));
  assign n847 = (~x3 | x4 | x5 | ~x0 | x1 | x2) & (x0 | ((x1 | ((~x2 | x3 | x4 | ~x5) & (x2 | ~x3 | ~x4 | x5))) & (~x1 | x2 | ~x3 | ~x4 | ~x5)));
  assign z070 = n849 | ~n854 | (~n179 & ~n852) | (~n164 & ~n853);
  assign n849 = ~x1 & (x0 ? ~n851 : ~n850);
  assign n850 = (x4 | ((x2 | x5 | (x3 ? (x6 | x7) : (~x6 | ~x7))) & (~x2 | ~x3 | ~x6 | x7))) & (~x2 | x3 | ((~x5 | ~x7) & (~x4 | x5 | x7)));
  assign n851 = (~x4 | x6 | ((x2 | ~x3 | x5 | ~x7) & (~x2 | x3 | ~x5 | x7))) & (x2 | x3 | ((x5 | ~x6 | x7) & (x4 | (x5 ^ x7))));
  assign n852 = (x1 | ((~x0 | ((x2 | ~x3 | x5) & (~x2 | x3 | x4 | ~x5))) & (x2 | x3 | ~x4 | x5) & (~x3 | ((x2 | ~x4 | ~x5) & (x0 | (~x2 ^ x5)))))) & (x0 | ~x1 | ((~x2 | (x3 ? ~x5 : (x4 | x5))) & (x3 | ~x4 | ~x5) & (x2 | (x3 ? (~x4 | x5) : ~x5))));
  assign n853 = (x3 | ((x0 | (x1 ? (x2 ? (x4 | ~x5) : (~x4 | x5)) : (x2 | ~x5))) & (x1 | (x2 ? (x5 | (~x0 & x4)) : (~x4 | ~x5))))) & (~x3 | ~x4 | x5 | x0 | ~x1 | ~x2);
  assign n854 = (~n152 | n856) & (n855 | (x5 ? (~x6 | x7) : (x6 | ~x7)));
  assign n855 = (x1 | x2 | ~x3 | x4) & (x0 | (x1 ? (~x2 | (~x3 ^ x4)) : (~x3 | ~x4)));
  assign n856 = (x5 | ((~x2 | x3 | ~x4 | ~x6 | ~x7) & (x2 | (x3 ? (~x6 | x7) : (x4 | ~x7))))) & (~x3 | ~x5 | x6 | (x4 ? ~x7 : x2));
  assign z071 = ~n862 | (~x3 & ~n861) | (~x1 & ~n858);
  assign n858 = (n293 | n860) & (~n545 | ~n822) & (~x3 | n859);
  assign n859 = x7 ? ((~x0 | x2 | x4 | x6) & (x0 | (x2 ? (x6 | (~x4 & ~x5)) : ~x6))) : ((x2 | (x0 ? (~x6 | (x4 & x5)) : (~x4 | x6))) & (x0 | ~x2 | (x4 ? ~x6 : (x5 | x6))));
  assign n860 = (x0 | ~x2 | ~x3 | x4 | ~x6) & (x2 | ((x4 | x6 | x0 | ~x3) & (~x0 | ~x4 | (~x3 ^ x6))));
  assign n861 = (x1 | (x0 ? (x4 | (~x2 ^ ~x6)) : (x2 ? (~x5 | x6) : ~x6))) & (x0 | ((~x1 | x4 | ~x5 | (x2 & ~x6)) & (~x4 | (x2 ? x6 : (x5 | ~x6)))));
  assign n862 = (~x4 | n863 | ~x0 | x1) & (x0 | ~x1 | (n864 & (x4 | n863)));
  assign n863 = (x5 | ~x6 | ~x2 | x3) & (x2 | (x3 ? (~x5 | ~x6) : (x5 | x6)));
  assign n864 = (~x4 | ((~x6 | (x2 ? (x3 ? x7 : (~x5 | ~x7)) : (x3 ? ~x7 : (~x5 | x7)))) & (~x3 | x6 | ((x7 | (x2 & x5)) & (~x2 | ~x5 | ~x7))))) & (~x3 | x4 | (x2 ? (x6 ^ x7) : ((x6 | ~x7) & (x5 | ~x6 | x7))));
  assign z072 = n867 | n868 | n869 | ~n870 | (n260 & ~n866);
  assign n866 = (~x7 | (~x3 ^ x6) | (x0 ? (x1 | x2) : ~x1)) & (~x0 | x1 | x7 | ((x3 | x6) & (x2 | ~x3 | ~x6)));
  assign n867 = (~x1 | (~x0 & ~x4)) & (~x0 | (~x2 & ~x4)) & (x3 | ~x7) & (~x3 | x7) & (x0 | x1 | x2 | x4);
  assign n868 = n530 & ((~x0 & x1 & x3 & x7) | (x0 & ~x1 & ((~x3 & ~x7) | (~x2 & x3 & x7))));
  assign n869 = ~x0 & ((x4 & ~x7 & x1 & ~x3) | (~x1 & ~x2 & x3 & ~x4 & x7));
  assign n870 = ~n873 & (~n545 | ~n872) & (~n186 | ~n871 | ~n404);
  assign n871 = x5 & ~x7;
  assign n872 = ~x3 & ~x2 & ~x0 & ~x1;
  assign n873 = ~x7 & ~x4 & ~x3 & x2 & x0 & ~x1;
  assign z073 = n875 | n878 | ~n880 | (~x0 & ~n879);
  assign n875 = ~x1 & (n877 | (~x5 & ~n876));
  assign n876 = (~x0 | ~x2 | x3 | x4) & (x0 | x2 | x6 | x7 | (~x3 ^ x4));
  assign n877 = ~x6 & x5 & ~x4 & x0 & x2 & ~x3;
  assign n878 = ~x1 & ((~x2 & ((~x4 & (x5 ^ x6)) | (x0 & (x4 ? (x5 & x6) : ~x6)))) | (~x0 & ~x4 & (x2 | x6)));
  assign n879 = (x1 | x2 | x4 | x5 | x6 | ~x7) & (~x1 | ~x5 | ~x6 | (~x4 ^ ~x7));
  assign n880 = x4 | ~n152 | (x5 & x6 & (~x7 | ~n272));
  assign z074 = n883 | ~n886 | (~x1 & ~n884) | (~x0 & ~n882);
  assign n882 = x1 ? (~x6 | (x5 ? (~x7 | (~x2 & ~x4)) : x7)) : (x2 | x6 | ((x5 | ~x7) & (x4 | ~x5 | x7)));
  assign n883 = ~x1 & (x0 ? (~x2 & (~x5 ^ x6)) : (~x5 & (x2 | x6)));
  assign n884 = (x0 | x2 | ~x3 | x7 | ~n154) & (~x0 | ~x2 | x3 | (~n154 & ~n885));
  assign n885 = x6 & ~x4 & x5;
  assign n886 = x0 | ~x1 | (~n154 & (~n247 | ~n573));
  assign z075 = ~n891 | (~x0 & (n889 | ~n890 | (~x2 & ~n888)));
  assign n888 = x1 ? (~x3 | ((~x6 | ~x7 | x4 | ~x5) & (x6 | x7 | ~x4 | x5))) : (x3 | ((x5 | ((x6 | ~x7) & (~x4 | ~x6 | x7))) & (x4 | ~x5 | ~x6 | x7)));
  assign n889 = ~x4 & (x1 ? (x6 ? (x7 & (x2 | ~x5)) : ~x7) : (~x2 & (x5 ? (~x6 & x7) : (x6 & ~x7))));
  assign n890 = ~x1 | ~x4 | (~n230 & (~n140 | (~x5 & ~n248)));
  assign n891 = (~n892 | ~n894) & (~n261 | ~n448) & (x1 | n893);
  assign n892 = ~x2 & ~x0 & x1;
  assign n893 = x6 ? (~x0 | (x2 & (x3 | (x4 & x5)))) : (x0 | (~x2 & (x5 ? ~x4 : ~x3)));
  assign n894 = ~x6 & ~x5 & ~x3 & x4;
  assign z076 = n896 | ~n901 | (~n304 & ~n899) | (n147 & ~n900);
  assign n896 = ~x3 & (x7 ? (n303 & ~n898) : ~n897);
  assign n897 = (x1 | ((~x4 | ~x5 | x0 | x2) & (~x0 | ((x2 | ~x4 | x5 | ~x6) & (~x2 | x4 | ~x5 | x6))))) & (x0 | ~x1 | x2 | (x4 ? (x5 | x6) : (~x5 | ~x6)));
  assign n898 = (x1 | ~x4 | x5 | x6) & (~x1 | (x4 ? (~x5 | x6) : (x5 | ~x6)));
  assign n899 = (x1 | (x2 ? (x7 | (x0 & (x3 | x5))) : ((~x3 | x5 | x7) & (~x0 | ((~x5 | x7) & (x3 | x5 | ~x7)))))) & (x0 | ~x1 | (~x7 & (x2 | x3 | x5)));
  assign n900 = (~x6 | ((x1 | x2 | ((~x5 | x7) & (x4 | x5 | ~x7))) & (~x1 | ~x2 | x4 | x5 | ~x7))) & (~x1 | ~x2 | ~x4 | x6 | (x5 ^ x7));
  assign n901 = (n215 | n902) & (x2 | ~n141 | n903);
  assign n902 = (x0 | (x1 ? (~x7 | (~x2 ^ x3)) : (~x2 | x7))) & (x1 | x7 | (x2 ? x3 : ~x0));
  assign n903 = (~x3 | ~x4 | x6 | x7) & (x3 | x4 | ~x7);
  assign z077 = n906 | ~n907 | (~x0 & (~n905 | ~n908 | ~n909));
  assign n905 = (~x1 | ((x2 | ~x3) & (~x2 | x3 | ~x4 | x5))) & (x2 | ~x4 | (~x3 & ~x5)) & (x1 | ~x2 | x3 | x4 | ~x5);
  assign n906 = ~x3 & ~x5 & n207 & (x2 ? (~x4 & ~x6) : (x4 ^ x6));
  assign n907 = x2 | ~n207 | ((~x3 | x4) & ~x5 & (x3 | ~x4 | ~n264));
  assign n908 = (x5 | (x1 ? ((x2 | x3 | x4 | ~x6) & (~x2 | ~x3 | ~x4 | x6)) : (x6 | (x2 ? (x3 | ~x4) : (~x3 | x4))))) & (x2 | x4 | ~x5 | (x1 ? (x3 | x6) : (~x3 | ~x6)));
  assign n909 = (n910 | n912) & (~n679 | ~n448) & (~n230 | n911);
  assign n910 = ~x2 ^ x7;
  assign n911 = (x1 | ~x2 | x3 | x4 | x5) & (~x1 | ((x2 | x3 | ~x4 | x5) & (x4 | ~x5 | ~x2 | ~x3)));
  assign n912 = (~x1 | x3 | x4 | x5 | x6) & (x1 | ((x5 | ~x6 | x3 | ~x4) & (~x3 | x4 | ~x5 | x6)));
  assign z078 = n915 | n918 | n919 | ~n921 | (n914 & n920);
  assign n914 = ~x4 & ~x2 & x0 & ~x1;
  assign n915 = ~x0 & ((n139 & ~n917) | (~x5 & ~n916));
  assign n916 = ((~x3 ^ x7) | ((x1 | ~x4 | ~x6) & (x4 | x6))) & (x2 | x3 | ~x4 | ~x6 | ~x7);
  assign n917 = x1 ? (~x6 | ((~x3 | ~x7) & (~x2 | x3 | x7))) : (x6 | (x3 ^ x7));
  assign n918 = ~x0 & ((~x1 & x3 & (x4 ? (~x5 & ~x6) : (x5 & x6))) | (~x3 & ~x4 & ((~x5 & x6) | (x1 & x5 & ~x6))));
  assign n919 = x4 & ((~x0 & ((~x3 & x5) | (x1 & x3 & ~x5))) | (~x1 & ~x2 & ((~x3 & x5) | (x0 & x3 & ~x5))));
  assign n920 = ~x6 & (x3 ^ x5);
  assign n921 = (~n261 | ~n923) & (~n922 | ~n319) & (~n389 | ~n190);
  assign n922 = x6 & ~x4 & ~x5;
  assign n923 = ~x7 & x6 & ~x4 & x5;
  assign z079 = ~n929 | (~x1 & (n926 | ~n927 | (x6 & ~n925)));
  assign n925 = (~x4 | ~x5 | x7 | ~x0 | x2 | x3) & (x0 | ~x2 | ~x3 | x4 | x5 | ~x7);
  assign n926 = ~n164 & ((~x0 & x2 & n271) | (x3 & n260 & x0 & ~x2));
  assign n927 = ~n928 & (n591 | ((x0 | ~x7) & (~x0 | ~x2 | x3 | x7)));
  assign n928 = ~x2 & ~x6 & ((x0 & x5 & ~x7) | (~x0 & ~x4 & ~x5 & x7));
  assign n929 = (n215 | n930) & (~n152 | n931);
  assign n930 = (x1 | ((~x0 | x5 | (x2 & x3)) & (~x5 | (x0 & (x2 | x3 | ~x7))))) & (x0 | ((~x1 | ((x5 | x7) & (~x2 | ~x3 | ~x7))) & (~x5 | (~x7 & (x2 | x3)))));
  assign n931 = (x5 | ~x7 | ((x2 | (x4 & (x3 | ~x6))) & (x4 | (x3 & x6)))) & (~x4 | ~x5 | x7 | (~x2 & (~x3 | x6)));
  assign z080 = n937 | ~n938 | (~x0 & (~n933 | ~n936));
  assign n933 = x3 ? n934 : n935;
  assign n934 = (x6 | ((~x7 | ((x1 | (x4 ? x5 : ~x2)) & (x5 | (x4 ? x2 : ~x1)))) & (~x1 | x7 | (x2 ? (~x4 | x5) : (x4 | ~x5))))) & (~x5 | ~x6 | x7 | (x1 & (x2 | ~x4)));
  assign n935 = x4 ? ((~x6 | x7 | x2 | ~x5) & (x6 | ~x7 | ~x2 | x5)) : ((x5 | ((x1 | x2 | ~x6 | ~x7) & (~x1 | ((x6 | ~x7) & (x2 | ~x6 | x7))))) & (x1 | ~x5 | ((~x6 | x7) & (~x2 | x6 | ~x7))));
  assign n936 = (x3 | (x1 ? (x2 | (x4 ? (x5 | ~x7) : (~x5 | x7))) : (~x2 | (x4 ? (~x5 | x7) : (x5 | ~x7))))) & (x1 | x2 | ~x3 | x4 | x5 | ~x7);
  assign n937 = ~n420 & ((~x1 & ((~x2 & ~x4) | (x0 & (x3 ? ~x2 : ~x4)))) | (~x0 & ~x4 & (x2 ? x1 : x3)));
  assign n938 = (n179 | n940) & (~n261 | ~n573) & (~n153 | ~n939);
  assign n939 = ~x7 & ~x5 & ~x3 & x4;
  assign n940 = (x0 | ((x1 | ~x4 | x5) & (~x5 | ((~x2 | ~x3 | ~x4) & (~x1 | (~x2 & ~x4)))))) & (x1 | ~x4 | (x2 ? (x3 | x5) : (x5 ? ~x0 : ~x3)));
  assign z081 = n942 | n946 | ~n948 | (~n293 & ~n945);
  assign n942 = ~x2 & ((~x1 & ~n943) | (n152 & ~n944));
  assign n943 = x4 ? ((~x3 | ((~x5 | ~x6 | ~x7) & (x0 | x6 | x7))) & (~x6 | x7 | ~x0 | x5) & (x0 | ((x5 | x6 | x7) & (x3 | ~x6 | ~x7)))) : (x0 ? ((x5 | x6 | x7) & (~x6 | ~x7 | x3 | ~x5)) : (x5 ? (x6 | ~x7) : (~x6 | x7)));
  assign n944 = (x6 | ~x7 | ~x4 | ~x5) & (~x6 | ((~x4 | x5 | x7) & (~x3 | (x4 ? x7 : (~x5 | ~x7)))));
  assign n945 = (x0 | (x4 ? (~x6 | (x1 ^ (~x2 & ~x3))) : ((~x2 | x6) & (~x1 | (x6 & (~x2 | ~x3)))))) & (x1 | ((x2 | x3 | ~x4 | x6) & (~x0 | (x2 & x3) | (~x4 ^ x6))));
  assign n946 = x2 & ((n139 & n265 & n319) | (~x0 & ~n947));
  assign n947 = ((x5 ? (~x6 | ~x7) : (x6 | x7)) | (x1 ? x4 : (x3 | ~x4))) & (x1 | x4 | x5 | ~x6 | x7) & (~x1 | ((x3 | ~x7 | (~x4 ^ x6)) & (~x4 | ((~x3 | ~x5 | x6) & (x5 | ~x6 | x7)))));
  assign n948 = (x1 | n949) & (~x5 | ~x7 | ~n186 | ~n892);
  assign n949 = x0 ? (x3 | ((~x5 | ~x7 | x2 | ~x4) & (x5 | x7 | ~x2 | x4))) : (~x2 | ((x4 | ~x5 | ~x7) & (x5 | x7 | ~x3 | ~x4)));
  assign z082 = n952 | ~n954 | n959 | (~x0 & ~n951) | n961;
  assign n951 = (~x1 | x2 | ~x3 | x4 | x5 | x6) & (x3 | ((x1 | x2 | ~x4 | ~x5 | ~x6) & (~x2 | ((x1 | x4 | x5 | ~x6) & (~x1 | ~x5 | (~x4 ^ x6))))));
  assign n952 = ~n217 & ~n953;
  assign n953 = (x1 | ((x2 | ((~x0 | x6 | (x3 & x4)) & (~x6 | (x3 ? x0 : x4)))) & (x0 | ~x2 | x6 | (~x3 & ~x4)))) & (x0 | ((~x4 | ~x6 | ~x2 | x3) & (~x1 | ((~x2 | ~x3 | ~x6) & (x4 | x6 | x2 | x3)))));
  assign n954 = ~n956 & ~n958 & (~n692 | n957) & (~n153 | ~n955);
  assign n955 = x6 & ~x5 & ~x3 & x4;
  assign n956 = ~x1 & ((x3 & x5 & ~x6 & ~x0 & ~x2) | (x0 & ~x5 & (x2 ? (~x3 & ~x6) : (x3 & x6))));
  assign n957 = (x0 | ~x2 | x4 | ~x5 | x6 | ~x7) & (~x0 | ~x4 | ~x6 | (x2 ? (x5 | ~x7) : (~x5 | x7)));
  assign n958 = x6 & x5 & x3 & ~x2 & ~x0 & x1;
  assign n959 = ~n293 & ~n960;
  assign n960 = (~x0 | x1 | ~x2 | x3 | x4 | ~x6) & (x0 | (x1 ? (x2 ? (x4 | x6) : (x6 ? x3 : ~x4)) : ((x2 | x3 | x6) & (~x4 | ~x6 | ~x2 | ~x3))));
  assign n961 = x3 & ((~x1 & ~n962) | (x7 & n152 & ~n963));
  assign n962 = (x0 | ~x2 | x4 | ~x6 | x7) & (x2 | ((x0 | x4 | x5 | x6 | ~x7) & (~x0 | ~x4 | x7 | (x5 ^ x6))));
  assign n963 = (~x2 | ~x4 | x6) & (x2 | x4 | x5 | ~x6);
  assign z083 = n965 | ~n970 | (~n164 & ~n968) | (n152 & ~n969);
  assign n965 = ~x1 & (x7 ? ~n967 : ~n966);
  assign n966 = ((x0 ? (x2 | x5) : (~x2 | ~x5)) | (x3 ? (x4 | x6) : (~x4 | ~x6))) & (~x4 | ~x5 | x6 | ~x0 | x3) & (x0 | x4 | ((~x2 | x5 | (~x3 ^ ~x6)) & (x2 | x3 | ~x5 | x6)));
  assign n967 = (x2 | ((x4 | x5 | x0 | ~x3) & (~x4 | ~x5 | x6 | ~x0 | x3))) & (x0 | ~x3 | x4 | ((x5 | ~x6) & (~x2 | ~x5 | x6)));
  assign n968 = (x1 | ((x0 | x3 | ~x4 | x5) & (x2 | (x0 ? (~x3 | (x4 & x5)) : (x3 | ~x4))))) & (x0 | ((x3 | x4 | ((~x2 | ~x5) & (~x1 | (~x2 & ~x5)))) & (~x1 | ~x3 | ~x4 | (x2 & x5))));
  assign n969 = (~x4 | ((~x2 | ~x5 | (x3 ? ~x6 : (x6 | x7))) & (x2 | x3 | x5 | ~x6 | x7))) & (x2 | x4 | x6 | (x3 ? (~x5 | x7) : x5));
  assign n970 = (~x7 | ((~n722 | n972) & (~x6 | n971))) & n973 & (x6 | x7 | n971);
  assign n971 = (x1 | ((~x0 | ~x2 | x3 | (x4 & x5)) & (x2 | ~x3 | ((~x4 | ~x5) & (x0 | (~x4 & ~x5)))))) & (x0 | ~x1 | (x2 ? (~x4 | x5) : (x4 | (~x3 ^ x5))));
  assign n972 = (~x4 | ~x6 | ~x1 | x2) & (x1 | (x2 ? (~x4 | ~x6) : (x4 | x6)));
  assign n973 = (~x0 | x1 | x2 | x3 | x4 | ~x6) & (x0 | ~x2 | ~x3 | x6 | (~x1 ^ x4));
  assign z084 = n976 | n977 | ~n978 | (n655 & ~n975);
  assign n975 = (~x5 | x6 | x7 | ~x0 | x1 | ~x2) & (x0 | ((x1 | ~x2 | x5 | x6 | x7) & (~x6 | ((x1 | ~x2 | x5 | ~x7) & (~x1 | ~x5 | (~x2 ^ ~x7))))));
  assign n976 = ~x2 & ((~x7 & ((~x1 & x3 & x4) | (~x0 & (x3 | (~x1 & x4))))) | (~x3 & x7 & (x0 ? ~x1 : ~x4)));
  assign n977 = x2 & ((~x4 & ~x7 & ~x1 & ~x3) | (~x0 & ((x3 & x7) | (x1 & ~x3 & ~x7))));
  assign n978 = (x1 | n981) & (~n979 | ~n980) & (~n753 | ~n892);
  assign n979 = x3 & ~x2 & x0 & ~x1;
  assign n980 = ~x4 & ~x5 & (x6 ^ x7);
  assign n981 = (~x4 | ~x5 | ~x7 | x0 | ~x2 | x3) & (~x0 | x7 | ((x4 | ~x5 | x2 | ~x3) & (~x2 | x3 | ~x4 | x5)));
  assign z085 = ~n983 | (~n369 & ~n988) | (~x1 & ~x5 & ~n987);
  assign n983 = ~n984 & n986 & (~n985 | (~x3 & ~x6) | ~x5 | (x3 & x6));
  assign n984 = ~x0 & ((~x1 & ~x2 & ~x3 & x4) | (x3 & (~x4 | (x1 & x2))));
  assign n985 = x4 & ~x2 & ~x0 & x1;
  assign n986 = (x1 | ((x3 | ~x4 | ~x5 | x0 | ~x2) & (~x0 | x2 | ~x3 | (~x4 & ~x5)))) & (~x3 | ~x4 | x5 | x0 | ~x1 | x2);
  assign n987 = x0 ? (x4 | (x2 ? (x3 | x6) : (~x3 | ~x6))) : (~x2 | ~x4 | (~x3 ^ x6));
  assign n988 = (x4 | x5 | x7 | ~x0 | x1 | x3) & (x0 | ~x4 | ((~x5 | ~x7 | ~x1 | x3) & (x1 | ~x3 | x5 | x7)));
  assign z086 = n990 | n992 | n994 | ~n996 | (~x1 & ~n995);
  assign n990 = x3 & ((n153 & n923) | (~x0 & ~n991));
  assign n991 = (x5 | ~x6 | ~x7 | x1 | ~x2 | ~x4) & (x2 | ((~x1 | ((~x6 | ~x7 | x4 | ~x5) & (x6 | x7 | ~x4 | x5))) & (x1 | ~x4 | x5 | x6 | ~x7)));
  assign n992 = ~x3 & ((n152 & ~n188 & ~n369) | (~x1 & ~n993));
  assign n993 = x2 ? ((~x6 | ~x7 | x4 | x5) & (x0 | ~x5 | x7 | (x4 ^ x6))) : ((x4 | x5 | x6 | ~x7) & (~x4 | ((~x5 | x6 | x7) & (~x6 | ~x7 | ~x0 | x5))));
  assign n994 = n152 & ((~x5 & ((~x2 & x3 & ~x4 & ~x6) | (x2 & (x3 ? (x4 & x6) : ~x6)))) | (~x2 & x5 & x6 & (~x3 | x4)));
  assign n995 = ((~x5 ^ x6) | ((~x0 | x2 | x4) & (x0 | ~x2 | x3 | ~x4))) & (~x3 | ((~x5 | x6 | x2 | ~x4) & (x0 | ((x2 | x5 | ~x6) & (~x5 | x6 | ~x2 | x4)))));
  assign n996 = (~x0 | x1 | ~x2 | x3 | x4 | ~x5) & (x0 | ((~x3 | x4 | x5 | ~x1 | ~x2) & (x1 | ~x4 | (x2 ? (~x3 | ~x5) : (x3 | x5)))));
  assign z087 = n998 | ~n1003 | (~x1 & ~n1001) | (~n179 & ~n1002);
  assign n998 = ~x0 & (x3 ? ~n1000 : ~n999);
  assign n999 = (x2 | (((~x6 ^ x7) | ((~x4 | ~x5) & (~x1 | x4 | x5))) & (~x5 | x6 | x7 | x1 | x4))) & (x1 | ~x2 | x4 | x6 | (x5 ^ x7));
  assign n1000 = (x2 | ~x4 | x5 | (~x6 ^ x7)) & (~x5 | ~x6 | x7 | ~x1 | ~x2 | x4);
  assign n1001 = x6 ? ((x2 | ((~x3 | ~x4 | ~x5) & (x4 | (x0 ? (~x3 ^ x5) : (x3 | x5))))) & (x0 | ~x2 | ((x4 | ~x5) & (x3 | ~x4 | x5)))) : (x2 ? (x0 ? (x3 | (~x4 ^ x5)) : (~x3 | (x4 ^ x5))) : ((x0 | (x3 ? (x4 | ~x5) : (~x4 | x5))) & (~x4 | x5 | ~x0 | ~x3)));
  assign n1002 = (x1 | ((~x0 | x4 | (x2 ? (x3 | x5) : (~x3 | ~x5))) & (~x3 | ~x4 | x5 | x0 | ~x2))) & (x0 | ~x2 | x3 | ((~x4 | ~x5) & (~x1 | x4 | x5)));
  assign n1003 = (x0 | ~x1 | n1004) & (~x0 | x1 | x3 | n1005);
  assign n1004 = (~x4 | ((x5 | ~x6 | ~x2 | x3) & (x2 | (x3 ? (~x5 | ~x6) : (x5 | x6))))) & (x2 | ~x3 | x4 | x5 | ~x6) & (~x2 | x6 | ((x4 | ~x5) & (~x3 | (x4 & ~x5))));
  assign n1005 = (x2 | (~x6 ^ x7) | (~x4 ^ ~x5)) & (~x2 | ~x4 | x5 | ~x6 | x7);
  assign z088 = ~n1011 | (x1 ? (~x0 & ~n1016) : (~n1007 | ~n1015));
  assign n1007 = (x3 | (n1009 & (x6 | n1010))) & (~n1008 | ~n448) & (~x3 | ~x6 | n1010);
  assign n1008 = x3 & ~x0 & ~x2;
  assign n1009 = (x0 | x2 | x4 | x5 | ~x6) & (~x0 | x7 | ((x2 | x4 | ~x5 | ~x6) & (~x2 | ~x4 | x5 | x6)));
  assign n1010 = (~x5 | ~x7 | x0 | x4) & (~x0 | x2 | ~x4 | x5 | x7);
  assign n1011 = (~n152 | n1014) & (n733 | n1012) & (n293 | n1013);
  assign n1012 = x0 ? (x1 | x2 | (~x3 ^ x7)) : ((~x2 | x3 | ~x7) & (~x1 | ((x3 | ~x7) & (~x2 | ~x3 | x7))));
  assign n1013 = (~x0 | x1 | ~x2 | x3 | x4) & (x0 | ~x3 | ~x4 | (x1 & x2));
  assign n1014 = (x3 | ~x4 | x5 | x7) & (~x3 | x4 | ((~x5 | ~x7) & (x2 | x5 | x7)));
  assign n1015 = (~x7 | ((~x0 | ((x3 | ~x4 | x5) & (x4 | ~x5 | x2 | ~x3))) & (x0 | x2 | x3 | ~x4 | ~x5))) & (x0 | x7 | (x3 ? (x4 | (~x2 & ~x5)) : (~x4 | x5)));
  assign n1016 = (~x3 | x4 | ~x5 | x6 | x7) & (~x2 | x3 | ~x6 | (x4 ? (x5 | ~x7) : (~x5 | x7)));
  assign z089 = ~n1018 | n1026 | (~x1 & (n1021 | n1022 | ~n1023));
  assign n1018 = (x1 | n1020) & (~n1019 | ((~x2 | x4 | ~x7) & (~x4 | (x2 & x7))));
  assign n1019 = x6 & ~x0 & x1;
  assign n1020 = (x3 | ((~x0 | ((x4 | ~x6 | ~x7) & (x6 | x7 | ~x2 | ~x4))) & (x0 | x2 | x4 | x6 | ~x7))) & (~x6 | ((x0 | (~x4 & (x2 | x7))) & (x2 | ~x7 | (x4 ? ~x3 : ~x0))));
  assign n1021 = ~x0 & x2 & ((x4 & ~x5 & ~x6 & x7) | (~x4 & x5 & (x6 ^ x7)));
  assign n1022 = ~x4 & ~n656 & (x0 ? (~x3 & ~x7) : (x3 & x7));
  assign n1023 = ~n1025 & (~x7 | ~n1024 | (~x2 ^ x5));
  assign n1024 = x6 & x4 & x0 & ~x3;
  assign n1025 = x0 & ~x2 & ~x7 & (x4 ? (~x5 ^ x6) : (~x5 & x6));
  assign n1026 = n152 & ~n1027;
  assign n1027 = x5 ? ((x4 | x7 | ((x2 | x3) & x6)) & (~x6 | ~x7 | ~x2 | ~x4)) : (x7 ? ((x3 | ~x4 | x6) & (x2 | (~x4 ^ x6))) : ((~x3 | x4 | ~x6) & (~x2 | ((x4 | ~x6) & (~x3 | ~x4 | x6)))));
  assign z090 = (~x7 | ~n1032) & (x7 | n1029 | n1030 | ~n1031);
  assign n1029 = ~n215 & ((~x0 & ~x2 & ~x3 & ~x5) | (~x1 & (x0 ? (x5 & (~x2 | ~x3)) : ~x5)));
  assign n1030 = n272 & ((x6 & n152 & x4 & ~x5) | (~x4 & x5 & ~x6 & n207));
  assign n1031 = (~x4 | x5 | (x0 ? (x1 | (x2 & x3)) : (~x1 | (~x2 & ~x3)))) & (x0 | x4 | ~x5);
  assign n1032 = n1034 & (x0 | x5 | n1033);
  assign n1033 = x1 ? ((x3 | x4 | x6) & (x2 | (x4 ^ x6))) : (~x2 | ((~x4 | ~x6) & (~x3 | x4 | x6)));
  assign n1034 = (x1 | ((~x0 | x4 | x5 | (x2 & x3)) & (x2 | ~x4 | (x0 & ~x5)))) & (x0 | ((~x4 | ~x5) & (~x3 | x4 | x5 | ~x1 | ~x2)));
  assign z091 = n1037 | n1038 | (~x0 & ~n1036) | ~n1039;
  assign n1036 = (~x1 & (x6 ? x5 : x7)) | (~x3 & (x2 | (x5 & x6 & x7))) | (~x2 & x3) | (~x5 & (x1 | ~x6));
  assign n1037 = ~n527 & ((x0 & ~x1 & ~x5 & ~x6 & ~x7) | (~x0 & ((~x1 & ~x5 & x6) | (x5 & ((~x6 & ~x7) | (x1 & (~x6 | ~x7)))))));
  assign n1038 = x7 & ~x6 & x5 & x2 & ~x0 & ~x1;
  assign n1039 = ~n1040 & (x3 | ((~n738 | ~n447) & (x4 | n1041)));
  assign n1040 = ~x2 & ((~x1 & ((~x0 & ~x5 & ~x6 & x7) | (x0 & x5 & (x6 | x7)))) | (~x0 & x1 & ~x5 & x6 & x7));
  assign n1041 = x0 ? (x1 | ~x5 | (~x2 ^ (~x6 & ~x7))) : (x5 | ((x1 | ~x2 | x6 | ~x7) & (~x1 | ~x6 | (~x2 ^ ~x7))));
  assign z092 = (x1 | n1043 | n1044 | ~n1045) & (~x1 | (~x0 & ~n1046));
  assign n1043 = ~n164 & (x2 ? (~x3 & ((~x4 & ~x5) | (x0 & (~x4 | ~x5)))) : (~x0 | x3 | (x4 & x5)));
  assign n1044 = ~x3 & ((~x0 & x2 & ~x4 & x5 & x6) | (x4 & ~x5 & ~x6 & x0 & ~x2));
  assign n1045 = (x3 | ((~x0 | x2 | x4 | x6) & (x0 | ~x2 | ~n680))) & (x0 | ~x2 | ~x6 | (~x3 & ~x4));
  assign n1046 = x6 ? ((x3 | x4 | ~x7) & (x2 | (~x7 & (x3 | x4 | x5)))) : ((~x2 | x7) & ((~x3 & ~x4) | (~x2 & x7)));
  assign z093 = ~n1051 | (~x3 & (~n1048 | n1049 | (n153 & n1050)));
  assign n1048 = (x7 | ((x2 | ~x4 | x5 | ~x0 | x1) & (x0 | x4 | (x1 ? (x2 | x5) : (~x2 | ~x5))))) & (~x0 | x1 | ~x4 | ~x7 | (~x2 ^ x5));
  assign n1049 = n233 & ((x5 & ~n179 & x1 & ~x2) | (~x1 & x2 & ~x5 & n265));
  assign n1050 = x7 & x6 & x4 & ~x5;
  assign n1051 = (x1 | ((~x0 | x3 | x4 | (~x2 ^ ~x7)) & (x2 | ~x7 | (x0 & ~x3)))) & (x0 | (((~x2 ^ x7) | (~x3 & ~x4)) & (~x1 | ~x2 | x3 | x4 | ~x7)));
  assign z094 = n1054 | n1056 | (~x0 & ~n1053) | ~n1057;
  assign n1053 = x1 ? ((x2 | x3 | x4 | ~x5 | x6) & (~x2 | ~x3 | ~x4 | x5 | ~x6)) : (x4 | x5 | (x2 ? (x3 | x6) : (~x3 | ~x6)));
  assign n1054 = ~n1055 & ~x7 & n692;
  assign n1055 = (~x0 | ~x4 | (x2 ? (~x5 | x6) : (x5 | ~x6))) & (x0 | ~x2 | x4 | x5 | ~x6);
  assign n1056 = ~x1 & ((x0 & ~x3 & (~x4 | (x2 & ~x5))) | (x3 & ((~x2 & x4 & x5) | (~x0 & (x4 | x5)))));
  assign n1057 = ~n1058 & (~n153 | ~n894) & (~n247 | ~n152 | ~n573);
  assign n1058 = ~x0 & x1 & (x3 ? (x4 & (~x2 | x5)) : (~x4 & (x2 | ~x5)));
  assign z095 = ~n1062 | ~n1064 | (~x0 & (n1061 | (n265 & ~n1060)));
  assign n1060 = (~x1 | ~x2 | ~x3 | x4 | x5) & (x1 | ~x4 | (x2 ? (~x3 | ~x5) : (x3 | x5)));
  assign n1061 = x6 & ~n720 & ((~x1 & x2 & ~x3 & ~x5) | (x3 & x5 & x1 & ~x2));
  assign n1062 = (~x5 | (n1063 & (~x2 | x4 | ~n152))) & (x4 | x5 | (x2 & x3) | ~n152);
  assign n1063 = (~x0 | x1 | ~x2 | x3 | x4 | ~x6) & (x0 | ((x1 | ~x2 | ~x3 | ~x4 | ~x6) & (~x1 | x2 | ((x3 | ~x4 | ~x6) & (x4 | x6)))));
  assign n1064 = ~n1066 & (~n207 | n1065) & (x5 | n1067);
  assign n1065 = (x5 | ~x6 | ~x7 | x2 | ~x3 | x4) & (x3 | ((~x2 | ~x5 | x6 | (~x4 ^ x7)) & (x5 | ~x6 | x7 | x2 | ~x4)));
  assign n1066 = ~x1 & (x5 ? (x0 ? (~x2 & ~x4) : (x4 & (~x2 | ~x3))) : ((x3 & ~x4 & ~x0 & x2) | (x0 & x4 & (x2 ^ x3))));
  assign n1067 = (((x2 | x3 | ~x0 | x1) & (x0 | ~x1 | ~x2 | ~x3)) | (~x4 ^ x6)) & (x0 | x1 | ((x4 | x6 | ~x2 | x3) & (x2 | ((~x4 | ~x6) & (~x3 | x4 | x6)))));
  assign z096 = n1079 | n1077 | n1075 | ~n1071 | n1069 | n1070;
  assign n1069 = ~x0 & ((~x3 & ((~x1 & ~x2 & x5 & x6) | (x1 & (x2 ? (x5 & ~x6) : (~x5 & x6))))) | (~x1 & x3 & ~x5 & (x2 ^ ~x6)));
  assign n1070 = ~x0 & ((~x1 & x2 & ~x5 & ~x6) | (x1 & x5 & (~x2 ^ x6)));
  assign n1071 = (~x2 | x6 | (x7 ? ~n1072 : n1073)) & n1074 & (x2 | ~x6 | (x7 ? n1073 : ~n1072));
  assign n1072 = x5 & x3 & ~x0 & x1;
  assign n1073 = (x0 | ~x1 | ~x3 | x5) & (x3 | ~x5 | ~x0 | x1);
  assign n1074 = ~x0 | x1 | x5 | (x2 ? (x3 | ~x6) : x6);
  assign n1075 = n207 & ~n1076;
  assign n1076 = (x5 | x6 | x7 | ~x2 | x3 | x4) & (x2 | ~x6 | ((x3 | x7 | (~x4 ^ x5)) & (~x3 | ~x4 | x5 | ~x7)));
  assign n1077 = ~x1 & ~n1078;
  assign n1078 = (x5 | ((x0 | ~x2 | x3 | ~x6 | x7) & (~x0 | ((~x2 | x3 | x6 | ~x7) & (x2 | ~x3 | ~x6 | x7))))) & (x0 | x2 | ~x5 | ~x7 | (x3 ^ x6));
  assign n1079 = ~x0 & ((n784 & ~n1080 & x5 & x6) | (~x6 & ~n1081));
  assign n1080 = x2 ? (x3 | ~x7) : (~x3 | x7);
  assign n1081 = ((x2 ? (~x3 | ~x4) : (x3 | x4)) | (x1 ? (x5 | ~x7) : (~x5 | x7))) & (~x4 | x5 | x7 | x1 | x2 | x3);
  assign z097 = ~n1093 | n1091 | n1090 | n1088 | n1083 | n1086;
  assign n1083 = ~x2 & ((~x1 & ~n1084) | (~x4 & n152 & ~n1085));
  assign n1084 = (x0 | ~x3 | x4 | x5 | x6 | ~x7) & (~x5 | (x0 ? ((~x3 | x4 | x6 | ~x7) & (x3 | ~x4 | ~x6 | x7)) : ((~x3 | ~x4 | ~x6 | x7) & (x3 | (x4 ? (x6 | x7) : (~x6 | ~x7))))));
  assign n1085 = (x3 | ~x5 | x6 | ~x7) & (~x6 | x7 | ~x3 | x5);
  assign n1086 = ~x1 & ~n1087;
  assign n1087 = x2 ? (~x6 | ((x4 | x5 | ~x0 | x3) & (x0 | ~x4 | (~x3 ^ x5)))) : ((x0 | x3 | x4 | x5 | ~x6) & (~x5 | ((~x0 | (x3 ? (x4 | ~x6) : (~x4 | x6))) & (x4 | x6 | x0 | ~x3))));
  assign n1088 = ~n164 & ~n1089;
  assign n1089 = (x1 | ((x3 | x4 | x0 | ~x2) & (x5 | (x0 ? (x2 | (~x3 ^ x4)) : (~x2 | x3))))) & (x0 | ~x1 | x2 | ~x3 | (~x4 & ~x5));
  assign n1090 = ~x1 & ((~x0 & x2 & x3 & ~x4 & x6) | (~x2 & ((x4 & ~x6 & ~x0 & x3) | (x0 & (x3 ? (x4 & x6) : (~x4 & ~x6))))));
  assign n1091 = ~n179 & ~n1092;
  assign n1092 = (x1 | ((x0 | x2 | x5 | (~x3 ^ x4)) & (~x2 | ((~x4 | ~x5 | x0 | ~x3) & (~x0 | x3 | (~x4 ^ x5)))))) & (x0 | ~x1 | (x2 ? (~x3 | (x4 & x5)) : (x3 | x4)));
  assign n1093 = ~n1096 & (n1094 | ~n1095) & (~n154 | ~n654 | ~n892);
  assign n1094 = (x3 | ~x5 | x7 | ~x0 | x1) & (x0 | ~x1 | ~x3 | (~x5 ^ x7));
  assign n1095 = x2 & x4 & ~x6;
  assign n1096 = ~x0 & x1 & ~x3 & (x2 ? x6 : (x4 & ~x6));
  assign z098 = n1098 | n1101 | (x1 ? (~x0 & ~n1104) : ~n1103);
  assign n1098 = x5 & (x3 ? ~n1099 : ~n1100);
  assign n1099 = (((x2 | x4 | ~x0 | x1) & (x0 | ~x1 | ~x2 | ~x4)) | (x6 ^ x7)) & (x0 | x2 | ((x1 | ~x4 | (~x6 ^ x7)) & (~x6 | ~x7 | ~x1 | x4)));
  assign n1100 = (x1 | ((x2 | x4 | x6 | ~x7) & (~x4 | ((~x6 | ~x7 | x0 | x2) & (~x0 | x7 | (~x2 ^ x6)))))) & (x0 | x2 | x4 | (~x6 ^ x7));
  assign n1101 = ~x5 & ((n230 & n153 & n655) | (~x0 & ~n1102));
  assign n1102 = (x2 | ~x3 | x4 | ~x6 | x7) & (x6 | ((~x1 | x3 | x7 | (x2 ^ ~x4)) & (~x3 | ~x7 | (~x2 ^ ~x4))));
  assign n1103 = x3 ? ((x2 | ((~x4 | x5 | ~x7) & (~x0 | (x4 ? ~x7 : (x5 | x7))))) & (x0 | ((x4 | ~x5 | ~x7) & (~x2 | (x4 ? (~x5 | x7) : ~x7))))) : ((x2 | ((x4 | x5 | ~x7) & (x0 | ~x4 | x7))) & (~x2 | ((x4 | ~x5 | x7) & (x0 | ((x5 | x7) & (~x4 | ~x5 | ~x7))))) & (x5 | ((~x4 | x7) & (~x0 | x4 | ~x7))));
  assign n1104 = (~x7 & ((~x3 & (x4 | x5)) | (x2 & (~x3 | (x4 & x5))))) | (x3 & x7) | (~x2 & ~x4 & (x7 | (x3 & ~x5)));
  assign z099 = n1106 | ~n1110 | (n207 & ~n1109);
  assign n1106 = ~x0 & (x4 ? ~n1107 : ~n1108);
  assign n1107 = x1 ? (x5 | ((x2 | x3 | x6 | ~x7) & (~x2 | (x3 ? (x6 | ~x7) : (~x6 | x7))))) : ((x2 | x3 | ~x5 | ~x6 | ~x7) & (~x3 | ((x6 | x7 | x2 | x5) & (~x2 | ~x6 | (~x5 ^ x7)))));
  assign n1108 = x1 ? ((x2 | ~x3 | ~x5 | ~x6 | x7) & (~x2 | x3 | x5 | x6 | ~x7)) : (~x2 | x5 | (x3 ? (x6 | x7) : (~x6 | ~x7)));
  assign n1109 = (x3 | ((~x4 | x6 | (x2 ? (x5 | x7) : (~x5 | ~x7))) & (x2 | ~x6 | ((x5 | x7) & (x4 | ~x5 | ~x7))))) & (x5 | x6 | x7 | x2 | ~x3 | x4);
  assign n1110 = n1113 & (x2 ? (x0 | n1112) : n1111);
  assign n1111 = (x1 | ((x0 | ((~x5 | ~x6 | x3 | x4) & (~x3 | (x4 ? (~x5 | ~x6) : (x5 | x6))))) & (x5 | x6 | x3 | ~x4) & (~x0 | ((x3 | ((x5 | x6) & (~x4 | ~x5 | ~x6))) & (~x4 | x5 | x6) & (~x5 | ~x6 | ~x3 | x4))))) & (x0 | ~x1 | ((x3 | ((~x5 | x6) & (~x4 | x5 | ~x6))) & (x4 | ((~x5 | x6) & (~x3 | x5 | ~x6)))));
  assign n1112 = (~x1 | ~x6 | (x3 ? (~x4 | ~x5) : (x4 | x5))) & (x6 | ((x1 | ~x3 | ~x5) & (x3 | (x1 ? (~x4 ^ x5) : (x4 | x5)))));
  assign n1113 = (x0 | ((x1 | ~x2 | x3 | ~x5) & (~x3 | ((x1 | x2 | x4 | ~x5) & (~x1 | x5 | (~x2 ^ x4)))))) & (x1 | ~x5 | ((~x2 | x3 | x4) & (~x3 | ~x4 | ~x0 | x2)));
  assign z100 = n1115 | n1117 | n1120 | ~n1121 | (~x1 & ~n1119);
  assign n1115 = ~n164 & ~n1116;
  assign n1116 = ((~x4 ^ x5) | ((~x2 | x3 | ~x0 | x1) & (x0 | x2 | (x1 ^ ~x3)))) & (x1 | ((~x3 | x4 | x5 | x0 | ~x2) & (x2 | ((~x0 | (x3 ? (x4 | x5) : (~x4 | ~x5))) & (x0 | x3 | x4 | x5))))) & (x0 | ~x1 | ((~x4 | ~x5 | x2 | ~x3) & (~x2 | x5 | (x3 ^ x4))));
  assign n1117 = x5 & ((n230 & n655 & n404) | (n140 & ~n1118));
  assign n1118 = (x0 | ~x1 | x2 | (~x3 & x4)) & (x1 | ((~x0 | ((x3 | x4) & (x2 | ~x3 | ~x4))) & (~x2 | x3 | x4) & (x0 | ~x4 | (x2 ^ x3))));
  assign n1119 = ((x2 ^ ~x4) | ((x0 | ~x6 | (x3 ^ x5)) & (x5 | x6 | ~x0 | x3))) & (x0 | ~x2 | x3 | ~x4 | x6) & (x2 | ~x6 | ((x4 | ~x5 | x0 | x3) & (~x0 | ~x3 | (~x4 ^ x5))));
  assign n1120 = n152 & (x3 ? (x2 ? (x4 ? (x5 & x6) : ~x6) : (~x5 & (x4 ^ x6))) : ((x5 & x6 & x2 & ~x4) | (~x2 & (x4 ? (x5 & x6) : (~x5 & ~x6)))));
  assign n1121 = (n1123 | ~n1124) & (x0 | n1122) & (~x0 | ~n177 | ~n431);
  assign n1122 = (x1 | ~x3 | ((~x6 | ~x7 | ~x2 | ~x4) & (x6 | x7 | x2 | x4))) & (~x4 | x6 | x7 | ~x1 | ~x2 | x3);
  assign n1123 = (x1 | x2 | x3 | x4) & (~x1 | ~x4 | (~x2 & x3));
  assign n1124 = x7 & x6 & ~x0 & ~x5;
  assign z101 = n1126 | n1129 | (x1 ? (~x0 & ~n1133) : ~n1132);
  assign n1126 = ~x4 & ((~x3 & ~n1127) | (n147 & ~n1128));
  assign n1127 = x5 ? (((x6 ^ x7) | (x0 ? (x1 | ~x2) : (~x1 | x2))) & (x0 | ~x2 | (x1 ? (~x6 | x7) : (x6 | ~x7)))) : ((~x0 | x1 | x2 | x6 | x7) & (x0 | ((x1 | ~x7 | (x2 ^ x6)) & (~x1 | x2 | ~x6 | x7))));
  assign n1128 = (~x1 | ~x2 | ~x5 | ~x6 | ~x7) & (x2 | (((~x5 ^ x6) | (~x1 ^ ~x7)) & (x6 | ~x7 | x1 | x5)));
  assign n1129 = x4 & (x3 ? ~n1130 : ~n1131);
  assign n1130 = (x1 | ((x5 | x6 | x7 | x0 | ~x2) & (x2 | ((~x5 | ~x6 | x7) & (~x0 | ~x7 | (~x5 ^ x6)))))) & (x0 | ~x1 | ((~x2 | x5 | (~x6 ^ x7)) & (x6 | x7 | x2 | ~x5)));
  assign n1131 = (x5 | ~x6 | x7 | ~x0 | x1 | x2) & (x0 | ~x7 | (~x1 ^ x6) | (x2 ^ x5));
  assign n1132 = (x2 | ((~x5 | ((~x0 | (x3 ? (x4 | x7) : ~x7)) & (x3 | ~x4 | ~x7) & (x0 | x4 | (~x3 ^ ~x7)))) & (~x0 | x5 | ((x4 | ~x7) & (~x3 | ~x4 | x7))))) & (x0 | ~x4 | x5 | (~x3 ^ ~x7)) & (~x2 | (x7 ? ((~x4 | x5 | ~x0 | x3) & (x0 | ~x3 | (~x4 & x5))) : ((x3 | x4 | x5) & (x0 | (x3 ? (x4 | ~x5) : ~x4)))));
  assign n1133 = (~x2 | (x3 ? (~x5 | x7) : (x5 | ~x7))) & (x2 | ((x3 | ~x4 | ~x5 | x7) & (~x3 | ((x5 | x7) & (~x4 | ~x5 | ~x7))))) & (~x3 | x4 | x5 | x7);
  assign z102 = n1135 | ~n1140 | (x0 ? (~x1 & ~n1139) : ~n1138);
  assign n1135 = ~x3 & ((~x1 & ~n1136) | (n152 & ~n1137));
  assign n1136 = x5 ? ((x0 | ~x6 | (x2 ? x7 : (~x4 | ~x7))) & (~x0 | ~x2 | ~x4 | x6 | x7)) : ((x2 | ((~x0 | (x4 ? (~x6 | ~x7) : (x6 | x7))) & (~x6 | x7 | x0 | x4))) & (x0 | ~x7 | ((~x2 | ~x4 | ~x6) & (x4 | x6))));
  assign n1137 = (x2 & (~x5 ^ x7)) | (~x2 & (x5 ^ x7)) | (x4 & ~x6) | (x6 & (~x4 | (~x5 & ~x7)));
  assign n1138 = ((~x3 ^ ~x6) | (x2 ? (~x5 | (x1 & ~x4)) : (~x4 | x5))) & (x1 | x2 | ~x3 | x5 | ~x6) & (x4 | ((x2 | ~x3 | x5 | x6) & (~x2 | ((x3 | x5 | ~x6) & (~x5 | x6 | ~x1 | ~x3)))));
  assign n1139 = (x3 | ((~x5 | ~x6 | x2 | x4) & (~x2 | ((x5 | ~x6) & (x4 | ~x5 | x6))))) & (x2 | ~x3 | (x4 ? x6 : x5));
  assign n1140 = (~n147 | n1142) & (n1141 | (x4 ? (x5 | x7) : (~x5 | ~x7)));
  assign n1141 = (x3 | ~x6 | x0 | x2) & (x1 | ((~x3 | x6 | x0 | ~x2) & (~x0 | x2 | (x3 ^ x6))));
  assign n1142 = x7 ? ((x2 | ~x4 | x5 | x6) & (~x2 | ((x4 | x5 | ~x6) & (~x5 | x6 | x1 | ~x4)))) : ((~x1 | x4 | ~x6 | (~x2 ^ ~x5)) & (x2 | ~x5 | x6 | (x1 & ~x4)));
  assign z103 = n1144 | ~n1147 | n1150 | n1153 | (x5 & ~n1146);
  assign n1144 = ~n164 & ~n1145;
  assign n1145 = (~x3 | ~x4 | x5 | ~x0 | x1 | x2) & (x0 | (x3 ? (x4 | ((~x2 | x5) & (~x1 | (~x2 & x5)))) : ((x1 | ~x4) & ((x2 & ~x5) | (x1 & ~x4)))));
  assign n1146 = (~x3 | ((~x0 | x1 | x2 | ~x4 | x6) & (x0 | ~x1 | (x2 ? (~x4 | x6) : (x4 | ~x6))))) & (~x0 | x1 | x3 | (x2 ? (x4 | x6) : (~x4 | ~x6)));
  assign n1147 = (n179 | n1149) & (~n613 | n1148);
  assign n1148 = (~x2 | x3 | x6) & (x2 | ~x3 | x4 | ~x6);
  assign n1149 = (x1 | (x0 ? (x2 | x3 | (x4 & x5)) : (~x3 | (~x4 & ~x5)))) & (x0 | ((x2 | ~x3 | ~x4) & (~x1 | x3 | x4 | (~x2 & x5))));
  assign n1150 = ~x7 & ((x5 & ~n1151) | (~x3 & ~x5 & n171 & ~n1152));
  assign n1151 = (x0 | ~x1 | x2 | x3 | x4) & (~x0 | x1 | ((x2 | ~x3 | x4 | ~x6) & (~x2 | x3 | ~x4 | x6)));
  assign n1152 = x1 ? (~x4 | ~x6) : (x4 | x6);
  assign n1153 = x7 & n147 & ~n1154;
  assign n1154 = (x1 | x2 | x4 | x5) & (~x1 | x6 | (x2 ? (~x4 | x5) : (x4 | ~x5)));
  assign z104 = n1157 | n1159 | n1160 | (~x1 & ~n1156) | ~n1161;
  assign n1156 = (x7 | ((x0 | ((x4 | ~x5) & (~x2 | ~x4 | x5))) & (x2 | ((x3 | x4 | ~x5) & (~x4 | x5 | (~x0 & ~x3)))))) & (~x0 | x3 | ~x4 | ~x7 | (~x2 ^ x5));
  assign n1157 = ~x5 & ((x4 & ~n179 & n428) | (~x3 & ~n1158));
  assign n1158 = (x0 | ~x1 | ~x2 | ~x4 | x6 | ~x7) & (x1 | x2 | ~x6 | ((x4 | x7) & (~x0 | ~x4 | ~x7)));
  assign n1159 = n152 & ((x2 & x3 & x4 & x5 & x7) | (~x7 & ((~x3 & ~x4 & x5) | (~x2 & (x4 ^ x5)))));
  assign n1160 = ~n733 & ((x3 & ((~x2 & x7 & x0 & ~x1) | (~x0 & ~x7 & (~x1 | ~x2)))) | (~x0 & ~x3 & ~x7 & (x1 | x2)));
  assign n1161 = ~n1162 & (~n190 | ~n752) & (~n139 | ~n265 | ~n979);
  assign n1162 = ~x0 & ~x7 & ((~x1 & ~x2 & ~x3 & x4) | (x3 & ~x4 & x1 & x2));
  assign z105 = n1164 | n1167 | n1168 | n1169 | (~x0 & ~n1166);
  assign n1164 = ~x3 & ((n190 & n196) | (~x5 & ~n1165));
  assign n1165 = (x1 | (x0 ? (x2 | (x4 ? (~x6 | ~x7) : (x6 | x7))) : (~x2 | ~x6 | (x4 ^ x7)))) & (x0 | ((x2 | x4 | x6 | ~x7) & (~x1 | ~x2 | ~x4 | ~x6 | x7)));
  assign n1166 = (~x2 | ((~x4 | (x1 ? (x3 ? (~x5 | ~x6) : (x5 | x6)) : (x3 | ~x5))) & (x1 | x4 | x5 | (~x3 & x6)))) & (x1 | ((x5 | x6 | ~x3 | x4) & (x2 | ((~x5 | ~x6) & (~x4 | x5 | x6)))));
  assign n1167 = ~n198 & ((~x1 & (x0 ? (~x4 & (x2 ^ x3)) : (~x2 & x4))) | (~x0 & ((~x2 & ~x3 & ~x4) | (x1 & x2 & x3 & x4))));
  assign n1168 = n207 & (x2 ? (~x3 & ((~x4 & x5 & x6) | (~x5 & (x4 | ~x6)))) : ((x4 & x5) | (x3 & ~x4 & ~x5 & ~x6)));
  assign n1169 = n177 & n1170 & (x0 ? n264 : n265);
  assign n1170 = x5 & x3 & ~x4;
  assign z106 = n1172 | n1175 | ~n1176 | n1179 | (~x4 & ~n1178);
  assign n1172 = ~x3 & ((~x1 & ~n1173) | (~x5 & n152 & ~n1174));
  assign n1173 = (x6 | ((~x0 | x7 | (x2 ? (~x4 | ~x5) : (x4 | x5))) & (~x2 | x4 | x5 | ~x7))) & (~x4 | x5 | ~x6 | ((x2 | ~x7) & (x0 | ~x2 | x7)));
  assign n1174 = x2 ? (x4 ? (~x6 | x7) : (x6 | ~x7)) : (x4 ? (~x6 | ~x7) : (x6 | x7));
  assign n1175 = ~x1 & (x2 ? ((~x0 & x3 & x4) | (~x3 & ((~x4 & x5) | (x0 & x4 & ~x5)))) : (x3 ? (~x4 & ~x5) : (x4 & x5)));
  assign n1176 = ~n1177 & (x3 | ~x4 | ~n154 | ~n171);
  assign n1177 = ~x0 & x1 & (x2 ? (x3 ? x4 : (~x4 & x5)) : (x3 ? (~x4 & ~x5) : (x4 & x5)));
  assign n1178 = (~x3 | ~x5 | ((~x0 | x1 | x2 | x6) & (x0 | (x1 ? (x2 | x6) : (~x2 | ~x6))))) & (~x2 | x3 | x5 | (x0 & x1) | ~x6);
  assign n1179 = n1170 & ((~x2 & x6 & ~x7 & x0 & ~x1) | (~x0 & (~x2 ^ x7) & (x1 ^ ~x6)));
  assign z107 = x3 ? (~n1187 | (~x4 & ~n1186)) : ~n1181;
  assign n1181 = ~n1182 & ~n1184 & (x7 ? (~n139 | n1185) : n1183);
  assign n1182 = ~x0 & x1 & ((x4 & ~x5 & ~x6) | (x5 & x6 & ~x2 & ~x4));
  assign n1183 = (x1 | ((x2 | ~x4 | x5 | ~x6) & (x6 | ((~x2 | x4 | x5) & (~x0 | ((x4 | x5) & (~x2 | ~x4 | ~x5))))))) & (x0 | x5 | ((~x4 | ~x6) & (~x1 | x4 | x6)));
  assign n1184 = ~x1 & ((x4 & ~x5 & (~x6 | (x0 & x2))) | (~x0 & ~x4 & x5 & x6));
  assign n1185 = x0 ? (x1 | ~x6) : (x1 ? (~x2 | ~x6) : x6);
  assign n1186 = (x1 | ((x6 | x7 | x0 | ~x5) & (x2 | ((x5 | x6 | ~x7) & (~x6 | x7 | ~x0 | ~x5))))) & (x0 | ((x5 | x6 | ~x7) & (~x6 | x7 | ~x1 | ~x5)));
  assign n1187 = (x4 | (x5 ? (x6 | n771) : (~x6 | n788))) & ~n1188 & (~x4 | ~x5 | n788);
  assign n1188 = x7 & x6 & ~x5 & ~x0 & x4;
  assign z108 = (~n590 & ~n1192) | (~x6 & ~n1190) | n1193 | (x6 & ~n1194);
  assign n1190 = (x3 | n1191) & (~n231 | (x1 ? (~x5 | ~x7) : (x5 | x7)));
  assign n1191 = (x1 | ((x4 | x5 | x7 | x0 | ~x2) & (~x0 | ~x5 | (x2 ? (~x4 | x7) : (x4 | ~x7))))) & (x0 | ~x1 | x4 | ((~x5 | ~x7) & (x2 | x5 | x7)));
  assign n1192 = (x0 & (x1 | x4)) | (x1 & (x2 ? (x3 & x4) : (~x3 & ~x4))) | (~x4 & (x7 | (~x1 & (~x0 | (x2 & x3)))));
  assign n1193 = ~n591 & ((~x0 & ~x7) | (~x1 & ((~x3 & ~x7) | (x0 & (x2 ^ x3)))));
  assign n1194 = n782 & (~n186 | ~n187 | ~n250);
  assign z109 = n1197 | ~n1199 | (~n293 & ~n1196) | (~x1 & ~n1198);
  assign n1196 = (x0 | (x6 ? x4 : ((x2 | x3 | ~x4) & (x1 | (~x4 & (x2 | x3)))))) & (x1 | ((x2 | x4 | ~x6) & (x3 | ((x4 | ~x6) & (~x2 | ~x4 | x6)))));
  assign n1197 = n152 & ((~x2 & ((~x5 & x6 & ~x7) | (~x4 & x5 & x7))) | (~x4 & ~x5 & ~x6 & ~x7) | (x4 & (x5 ? (~x6 & x7) : (x6 & ~x7))));
  assign n1198 = (x6 | ((~x0 | x2 | (x4 ? ~x7 : (x5 | x7))) & (x0 | ~x2 | x4 | x7))) & (x0 | ((~x4 | (x5 ? ~x7 : (~x6 | x7))) & (~x6 | ((~x5 | ~x7) & (~x2 | x5 | x7)))));
  assign n1199 = (~n448 | ~n763) & (x0 | (~n1202 & (n1200 | ~n1201)));
  assign n1200 = (~x2 | ~x3 | x5 | x6) & (x2 | x3 | ~x5 | ~x6);
  assign n1201 = x1 & x4 & x7;
  assign n1202 = ~x7 & ~x6 & ~x4 & x3 & ~x1 & ~x2;
  assign z110 = n1204 | ~n1207 | (~n179 & ~n1206);
  assign n1204 = ~x6 & ((~x5 & ~n1205) | (n186 & n250 & x5 & x7));
  assign n1205 = (x1 | ((x2 | (x0 ? (x3 | x7) : (~x3 | x4))) & (x0 | x3 | (x7 ? x4 : ~x2)))) & (x0 | ~x1 | ~x4 | ((~x3 | ~x7) & (~x2 | (~x3 & ~x7))));
  assign n1206 = (~x4 | ((x1 | ((~x0 | (x2 ? (x3 | x5) : ~x5)) & (x2 | x5 | (x0 & ~x3)))) & (x0 | ~x1 | ~x5 | (~x2 & ~x3)))) & (x0 | x4 | (x5 ? x1 : (~x1 & (~x2 | ~x3))));
  assign n1207 = (x5 | ~x6 | x7 | n1208) & (~x5 | ((x6 | ~x7 | n1208) & (x0 | ~x6 | n1209)));
  assign n1208 = (x0 | (~x4 & (~x1 | ~x2))) & (x1 | x4 | (x2 & (~x0 | x3)));
  assign n1209 = (x2 | (x1 ? (x4 | ~x7) : (~x4 | x7))) & (~x1 | x4 | x7 | (~x2 & ~x3));
  assign z111 = ~n1213 | (~x1 & (x2 ? ~n1212 : ~n1211));
  assign n1211 = x6 ? ((~x3 | x4 | (x0 ? (x5 | x7) : ~x7)) & (x0 | ((x3 | ~x5 | ~x7) & (~x4 | x5 | x7)))) : ((~x3 | ((x0 | x4 | ~x5 | x7) & (x5 | ~x7 | ~x0 | ~x4))) & (x3 | ~x4 | ~x5 | ~x7) & (~x0 | ((x4 | ~x5 | ~x7) & (x3 | ~x4 | x5 | x7))));
  assign n1212 = (x4 | ((~x0 | x3 | x5 | x6 | x7) & (x0 | ((x6 | x7 | x3 | ~x5) & (~x7 | ((~x5 | ~x6) & (~x3 | (~x5 & ~x6)))))))) & (x0 | ~x4 | x5 | x7 | (~x3 & ~x6));
  assign n1213 = (n188 | n1216) & (n293 | n1215) & (~n152 | n1214);
  assign n1214 = (x2 | ((~x3 | ~x4 | ~x5 | ~x6 | ~x7) & (x6 | x7 | x3 | x5))) & (x6 | x7 | ~x4 | x5) & (~x2 | ((x6 | x7 | ~x3 | ~x4) & (~x7 | ((x4 | ~x5 | x6) & (x3 | (x4 ? (x5 | ~x6) : ~x5))))));
  assign n1215 = (x0 | (x2 ? (x1 ? (x3 | x6) : ((~x4 | ~x6) & (~x3 | x4 | x6))) : ((x3 | x4 | x6) & (~x1 | (x6 ? ~x4 : ~x3))))) & (x1 | ((x3 | (~x0 & x2) | (~x4 ^ x6)) & (x4 | ~x6 | ~x0 | x2)));
  assign n1216 = (x0 | ~x2 | (~x1 ^ ~x6)) & (x1 | x2 | ((~x3 | x6) & (~x0 | x3 | ~x6)));
  assign z112 = ~n1220 | (x5 & (x2 ? ~n1219 : ~n1218));
  assign n1218 = (x4 | ~x6 | ((x0 | ~x1 | ~x3) & (x1 | x7 | (~x0 & ~x3)))) & (x6 | ~x7 | ((x1 | ~x4) & (x0 | (~x4 & (x1 | x3)))));
  assign n1219 = (x1 | x3 | ((x0 | ~x6 | x7) & (x6 | ~x7 | ~x0 | x4))) & (x0 | (x4 ? (~x6 | x7) : (x6 | ~x7 | (~x1 & ~x3))));
  assign n1220 = (n179 | n1221) & (x5 | (x3 ? n1223 : n1222));
  assign n1221 = (x1 | ((x5 | (x0 ? (x2 ? (x3 | ~x4) : ~x3) : (~x2 | (x3 ^ x4)))) & (x2 | ~x5 | (x4 ? ~x3 : (x0 & x3))))) & (x0 | (x3 ? ((x2 | ~x4 | ~x5) & (~x1 | x4 | (~x2 ^ ~x5))) : (~x5 | (x2 ^ x4))));
  assign n1222 = (x1 | ((~x0 | (x2 ? (x4 | x7) : ~x7)) & (x2 | (x4 ? (~x6 | x7) : (x6 | ~x7))) & (x0 | ((x4 | ~x6 | x7) & (~x2 | ~x4 | ~x7))))) & (x0 | ((~x1 | x4 | (~x2 ^ x7)) & (~x4 | (x2 ? (x6 | ~x7) : x7))));
  assign n1223 = (x2 | ((~x6 | x7 | x0 | ~x4) & (x6 | ((x1 | ~x4 | ~x7) & (x0 | ((~x4 | ~x7) & (x1 | x4 | x7))))))) & (x0 | ~x2 | ((x4 | (~x6 ^ x7)) & (~x6 | ~x7 | ~x1 | ~x4)));
  assign z113 = ~n1231 | (x3 ? (~n1226 | (~x1 & ~n1225)) : ~n1228);
  assign n1225 = x0 ? (x2 | ~x4 | (x5 ? (x6 | x7) : ~x6)) : (x4 | ((~x5 | ~x6 | x7) & (x6 | (x5 & (~x2 | ~x7)))));
  assign n1226 = (~x0 | x1 | x2 | n600) & (x0 | ((~x4 | n600) & (~x1 | (n1227 & (~x2 | n600)))));
  assign n1227 = (x2 | x4 | x5 | x6 | x7) & (~x4 | ((x5 | ~x6 | ~x7) & (x6 | x7 | ~x2 | ~x5)));
  assign n1228 = (x1 | n1229) & (~n1019 | n1230);
  assign n1229 = x0 ? (x2 | ~x4 | ((x6 | ~x7) & (~x5 | ~x6 | x7))) : (x4 | ((~x6 | ~x7) & (~x2 | (x5 ? (x6 | x7) : ~x6))));
  assign n1230 = (x2 | x4 | ~x7) & (~x2 | ~x4 | ~x5 | x7);
  assign n1231 = (n420 | n1233) & (n293 | n1232);
  assign n1232 = x0 ? (x1 | ((x3 | ((x4 | ~x6) & (~x2 | ~x4 | x6))) & (x4 | x6 | x2 | ~x3))) : (x4 ? ((x1 & x2) | (~x3 ^ x6)) : ((~x1 | ((~x2 | x3 | ~x6) & (~x3 | x6))) & (x1 | x2 | x3 | x6)));
  assign n1233 = (x1 | x4 | (x0 ? x3 : (x2 | ~x3))) & (x0 | x3 | (~x1 & ~x4));
  assign z114 = n1236 | n1237 | ~n1238 | (~x1 & ~n1235) | ~n1239;
  assign n1235 = (x3 & ((~x4 & x7) | (x2 & (x0 | (x4 & ~x7))))) | (x0 & ((x4 & ~x7) | (~x2 & ~x3 & x7))) | (~x5 & ~x7) | (x7 & (x5 | (~x0 & ~x4)));
  assign n1236 = n152 & ((x4 & n142 & n154) | (~x2 & n885));
  assign n1237 = (x4 ? n871 : n187) & (~n771 | (n141 & n142));
  assign n1238 = (~n753 | ~n892) & (~n153 | ~n894);
  assign n1239 = (n527 | n1240) & (~n233 | n1241);
  assign n1240 = (~x5 | ~x6 | ~x7 | x0 | x1 | x4) & (x5 | x6 | ((~x4 | x7 | ~x0 | x1) & (x0 | ~x7 | (~x1 ^ ~x4))));
  assign n1241 = (x1 | x2 | x3 | x5 | x6 | ~x7) & (~x5 | ~x6 | (x1 ? (~x2 | x7) : (~x7 | (~x2 ^ ~x3))));
  assign z115 = ~n1245 | (~x1 & (x7 ? ~n1243 : ~n1244));
  assign n1243 = (~x4 | ((x5 | ((x0 | x6 | (~x2 & ~x3)) & (~x0 | ~x2 | x3 | ~x6))) & (~x0 | x2 | ~x5 | (~x3 ^ x6)))) & (x0 | x4 | ((~x3 | ~x5 | x6) & (~x2 | ((~x5 | x6) & (~x3 | x5 | ~x6)))));
  assign n1244 = (x0 | ~x2 | x4 | ~x5 | ~x6) & (~x0 | ((x3 | x4 | x5 | ~x6) & (x2 | (x4 ? (x5 ^ x6) : (x5 | ~x6)))));
  assign n1245 = (x1 | n1020) & (~n152 | (n1246 & (~x6 | n1247)));
  assign n1246 = x5 ? (x4 ? (~x6 | (~x2 & ~x3) | ~x7) : (x6 | x7)) : (x7 ? ((x3 | ~x4 | x6) & (x2 | (~x4 ^ x6))) : ((~x3 | x4 | ~x6) & (~x2 | ((x4 | ~x6) & (~x3 | ~x4 | x6)))));
  assign n1247 = (~x4 | x7) & (~x2 | x4 | ~x7) & (x2 | x3 | (~x4 & x7));
  assign z116 = n1249 | (x5 ? (~n1253 | (n207 & ~n1254)) : ~n1252);
  assign n1249 = ~x0 & (x3 ? ~n1250 : (~x5 & ~n1251));
  assign n1250 = (x6 | (x1 ? ((x2 | x4 | x5 | ~x7) & (~x2 | ~x4 | ~x5 | x7)) : (x5 | (x2 ? (x4 | ~x7) : (~x4 | x7))))) & (x1 | x5 | ~x6 | (~x4 ^ ~x7));
  assign n1251 = (x1 | x7 | (~x4 ^ x6)) & (~x7 | (x4 ^ x6) | (~x1 ^ x2));
  assign n1252 = x0 ? (x1 | (x2 & x3) | (~x4 ^ x7)) : ((~x1 | ((~x4 | x7) & (~x2 | x4 | ~x7))) & (~x4 | ((~x2 | ~x3 | x7) & (x1 | x2 | x3 | ~x7))));
  assign n1253 = (x1 | x2 | x3 | ~x4 | ~x7) & (x0 | (x4 ^ x7));
  assign n1254 = x7 ? ((x4 | x6 | ~x2 | x3) & (x2 | ~x3 | ~x4 | ~x6)) : ((x2 & x3) | (~x4 ^ x6));
  assign z117 = ~n1263 | n1261 | n1260 | n1256 | n1259;
  assign n1256 = ~x0 & (n1258 | (x7 & ~n1257));
  assign n1257 = x2 ? (~x3 | ~x4 | (x1 ? (~x5 | x6) : (x5 | ~x6))) : (x5 | (x3 & x4) | (~x1 ^ ~x6));
  assign n1258 = x5 & ~x7 & ((~x3 & x6 & x1 & ~x2) | (~x1 & (x2 ? (x3 & x6) : (~x3 & ~x6))));
  assign n1259 = ~x0 & ((~x1 & x2 & ~x3 & ~x5 & x6) | (x5 & ((x1 & (x2 ? (~x3 & ~x6) : (x3 & x6))) | (~x1 & ~x2 & x3 & ~x6))));
  assign n1260 = ~x0 & ((~x1 & ~x2 & ~x5 & x6) | (x5 & (x1 ? (~x2 ^ x6) : (x2 & ~x6))));
  assign n1261 = ~n1262 & x2 & ~x4;
  assign n1262 = (~x0 | x1 | x3 | ~x5 | ~x6) & (x0 | ~x3 | (x1 ? (~x5 | x6) : (x5 | ~x6)));
  assign n1263 = n1265 & (x2 | x6 | ~n207 | n1264);
  assign n1264 = x7 ? ((x3 & x4) | ~x5) : x5;
  assign n1265 = ~x0 | x1 | ((x2 | ~x5 | ~x6) & (x5 | x6 | ~x2 | x3));
  assign z118 = n1272 | ~n1274 | (~x0 & ~n1267) | (x2 & ~n1271);
  assign n1267 = (~x6 | (x7 ? n1268 : n1269)) & (~x3 | n1270) & (x6 | (x7 ? n1269 : n1268));
  assign n1268 = x1 ? (x2 | (x3 & (x4 | x5))) : (~x2 | ~x3 | (~x4 & ~x5));
  assign n1269 = (x1 | x2 | x3) & (~x1 | ~x2 | ~x3 | ~x4 | ~x5);
  assign n1270 = (x1 | x2 | x4 | x5 | x6 | ~x7) & (~x1 | x7 | ((x2 | x4 | ~x5 | x6) & (x5 | ~x6 | ~x2 | ~x4)));
  assign n1271 = (x0 | (x1 ? (x6 | (x4 & (x3 | ~x5) & (~x3 | x5))) : (~x6 | (x3 ? (x4 | x5) : ~x5)))) & (~x0 | x1 | x3 | x4 | ~x6);
  assign n1272 = ~n1273 & (x2 ? (~x3 & ~x5) : (x3 & x5));
  assign n1273 = (x1 | ~x4 | ~x6) & (x0 | (x1 ? (~x4 | x6) : ~x6));
  assign n1274 = ((x3 & x4) | ~n1276) & (x5 | (~n1276 & (~x3 | ~n303 | n1275)));
  assign n1275 = x1 ? (~x4 | x6) : ~x6;
  assign n1276 = x0 & ~x1 & ~x2 & (x6 ^ x7);
  assign z119 = n1280 | ~n1282 | (x3 & (~n1278 | ~n1279));
  assign n1278 = (x1 | ((x2 | ((x0 | x4 | ~x5 | x7) & (~x0 | ~x4 | (~x5 ^ x7)))) & (x0 | ~x2 | x4 | (x5 ^ x7)))) & (x0 | ~x1 | ~x7 | (x2 ? (~x4 | ~x5) : (x4 | x5)));
  assign n1279 = (x1 | ~x7 | (x0 ? (x2 | x4) : (~x2 | ~x4))) & (x0 | x7 | ((x2 | ~x4) & (~x1 | ~x2 | x4)));
  assign n1280 = ~x6 & ((n655 & n871 & n190) | (n147 & ~n1281));
  assign n1281 = (x1 | x2 | x4 | x5 | ~x7) & (~x1 | ((x2 | x4 | ~x5 | ~x7) & (~x2 | ~x4 | x5 | x7)));
  assign n1282 = ~n1283 & (~n190 | ~n939) & (~n147 | ~n762 | n1284);
  assign n1283 = ~x3 & ((~x0 & (x2 ^ x7)) | (~x1 & (x2 ? (~x4 & ~x7) : x7)));
  assign n1284 = (~x1 | ~x2 | ~x4 | ~x7) & (x1 | x2 | x4 | x7);
  assign z120 = ~n1286 | (~x0 & ~n1289) | (n233 & ~n1290);
  assign n1286 = ~n1287 & (~n261 | ~n1050) & ~n1288;
  assign n1287 = ~x1 & ((~x2 & ((~x3 & x4 & x5) | (x0 & x3 & (~x4 | ~x5)))) | (~x0 & ((~x4 & ~x5) ? (x2 & x3) : ~x3)));
  assign n1288 = ~x0 & x1 & (x3 ? (~x4 & (x2 | ~x5)) : x4);
  assign n1289 = (~x4 | x5 | x6 | ~x1 | ~x2 | ~x3) & (x2 | x4 | (~x3 ^ x6) | (~x1 ^ ~x5));
  assign n1290 = (~x5 | ~x6 | x7 | ~x1 | x2 | ~x3) & (x1 | x3 | x5 | ~x7 | (~x2 ^ ~x6));
  assign z122 = z121;
  assign z123 = z121;
  assign z124 = z121;
  assign z125 = z121;
  assign z126 = z121;
  assign z127 = z121;
  assign z128 = z121;
endmodule


