// Benchmark "X_17" written by ABC on Wed Jun 07 02:57:10 2023

module X_17 ( 
    x0, x1, x2, x3,
    z0, z1, z2, z3, z4, z5, z6, z7  );
  input  x0, x1, x2, x3;
  output z0, z1, z2, z3, z4, z5, z6, z7;
  assign z0 = 1'b0;
  assign z1 = 1'b0;
  assign z2 = 1'b0;
  assign z3 = 1'b0;
  assign z4 = x0;
  assign z5 = x1;
  assign z6 = x2;
  assign z7 = x3;
endmodule


