// Benchmark "32_32_mod" written by ABC on Thu Dec 01 00:28:07 2022

module const_32_32_mod ( 
    x0, x1, x2, x3, x4, x5, x6,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63, z64  );
  input  x0, x1, x2, x3, x4, x5, x6;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63, z64;
  wire n74, n75, n76, n77, n79, n80, n81, n83, n84, n86, n87, n88, n89, n90,
    n91, n92, n94, n95, n96, n97, n99, n100, n101, n103, n104, n106, n107,
    n109, n110, n111, n113, n114, n115, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n127, n128, n130, n131, n132, n134, n135, n136, n138,
    n139, n140, n141, n142, n144, n145, n146, n147, n148, n149, n151, n152,
    n153, n154, n156, n157, n159, n160, n161, n162, n164, n165, n166, n167,
    n168, n170, n171, n173, n174, n175, n176, n177, n178, n179, n181, n182,
    n183, n185, n186, n187, n189, n190, n191, n193, n194, n195, n196, n198,
    n199, n200, n202, n203, n204, n205, n207, n208, n209, n210, n211, n213,
    n214, n215, n216, n217, n218, n219, n220, n221, n223, n224, n225, n226,
    n227, n228, n230, n231, n232, n233, n234, n236, n237, n238, n239, n241,
    n242, n243, n244, n245, n246, n248, n249, n250, n251, n253, n254, n255,
    n256, n258, n259, n260, n261, n262, n263, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n275, n276, n277, n279, n280, n281, n283, n284,
    n285, n286, n287, n288, n290, n291, n292, n293, n295, n296, n297, n298,
    n300, n301, n302, n303, n305, n306, n307, n309, n310, n311, n312, n313,
    n314, n316, n317, n319, n320, n321, n323, n324, n325, n327, n328, n329,
    n331, n332, n333, n334, n335, n337, n338, n339, n341, n342, n343, n344,
    n345, n346, n348, n349, n350;
  assign z58 = 1'b0;
  assign z00 = (~n74 & n75) | (~x5 & ~x6 & n76 & n77);
  assign n74 = (~x2 | ((~x3 | ~x4 | x5 | ~x6) & (x3 | x4 | ~x5 | x6))) & (x2 | x3 | ~x4 | ~x5 | ~x6);
  assign n75 = ~x0 & x1;
  assign n76 = ~x2 & x0 & ~x1;
  assign n77 = x3 & ~x4;
  assign z01 = ~n81 | (~x1 & (~n79 | ~n80));
  assign n79 = (~x5 | (((~x3 ^ x6) | (x0 ? (x2 | x4) : (~x2 | ~x4))) & (x0 | x2 | x3 | x4 | x6))) & (x4 | x5 | (x0 ? (x2 ? (x3 | x6) : (~x3 | ~x6)) : ((x3 | ~x6) & (x2 | ~x3 | x6))));
  assign n80 = (~x4 | ((x2 | (x0 ? (x3 ^ x5) : (x3 | ~x5))) & (x0 | ~x3 | x5))) & (x0 | ~x2 | (x3 ? x5 : (x4 | ~x5)));
  assign n81 = ~n75 | ((x2 | (x3 ? (x5 | ~x6) : (x4 | ~x5))) & (x3 | (x4 ? (x5 | x6) : (~x5 | ~x6))) & (~x3 | (x5 ? (~x4 & (~x2 | x6)) : x4)));
  assign z02 = (~x1 & ~n83) | (~x0 & x1 & ~n84);
  assign n83 = (x2 | (x4 ? ((~x3 | (~x5 & x6)) & (~x5 | x6)) : ((~x0 | (~x6 & (x3 | x5))) & (~x6 | (x3 & x5))))) & (x0 | ((~x2 | ((~x3 | ~x4 | ~x6) & (x4 | ~x5 | x6))) & (~x4 | (x5 ^ x6)))) & (x3 | x4 | x5 | ~x6);
  assign n84 = (x2 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (~x4 | ((x3 | x5 | ~x6) & (~x2 | ~x5 | x6))) & (x4 | ((~x2 | (x5 ^ x6)) & (~x3 | x5 | x6)));
  assign z03 = n87 | n88 | n89 | n91 | (~x0 & ~n86);
  assign n86 = x4 ? ((x1 | ((~x5 | ~x6 | ~x2 | x3) & (x5 | x6 | x2 | ~x3))) & (~x2 | ((~x5 | ~x6 | ~x1 | ~x3) & (x3 | x5 | x6)))) : ((~x1 | ((x2 | (x3 ? ~x5 : (x5 | x6))) & (~x2 | ~x3 | x5 | ~x6))) & (~x5 | ~x6 | x2 | x3));
  assign n87 = ~x1 & (((~x5 ^ x6) & (x0 ? (~x2 & ~x3) : (x2 & x3))) | (~x0 & ~x3 & (x2 ? (~x5 & x6) : (x5 & ~x6))) | (x0 & ~x2 & x3 & x5 & ~x6));
  assign n88 = ~x0 & x1 & ((x2 & ~x5 & (x3 ^ x6)) | (~x2 & ~x3 & x5 & ~x6));
  assign n89 = ~n90 & ((~x0 & ~x2 & x3 & (~x1 | x4)) | (x0 & ~x1 & x2 & ~x3 & ~x4));
  assign n90 = x5 ^ ~x6;
  assign n91 = n77 & n92 & n76;
  assign n92 = x5 & x6;
  assign z04 = ~n95 | (n94 & ~n97) | (~x2 & ~n96);
  assign n94 = ~x0 & x2;
  assign n95 = x0 ? (x1 | ((x2 | (x3 ? (x4 | ~x6) : x6)) & (x3 | x4 | x6))) : ((~x6 | (x1 ? ((~x3 | x4) & (~x2 | x3 | ~x4)) : (x3 | x4))) & (x1 | ~x3 | x6 | (~x2 & x4)));
  assign n96 = (x1 | ((~x0 | ~x6 | (x3 ? (~x4 | x5) : (x4 | ~x5))) & (~x4 | ~x5 | x6 | (x0 & ~x3)))) & (x0 | ((x3 | ((~x4 | x5 | ~x6) & (~x1 | x4 | (x5 ^ x6)))) & (~x5 | x6 | ~x3 | ~x4)));
  assign n97 = (~x1 | ~x5 | (x3 ? (~x4 | x6) : (x4 | ~x6))) & (x3 | x5 | ((x4 | x6) & (x1 | ~x4 | ~x6)));
  assign z05 = ~n101 | n99 | (~x0 & ~x5 & ~n100);
  assign n99 = ~x0 & ~x2 & ((~x1 & (x3 ? (x4 & x5) : (x4 ^ x5))) | (x1 & ~x3 & ~x4 & ~x5));
  assign n100 = (x1 | x2 | ~x6 | (~x3 ^ ~x4)) & (~x1 | ~x2 | ~x3 | ~x4 | x6);
  assign n101 = (x1 | (x0 ? (x2 | (~x3 ^ x4)) : (~x2 | (x3 ^ x4)))) & (x0 | ~x1 | ~x3 | (x2 & x4));
  assign z06 = ~n104 | (~x0 & ~n103);
  assign n103 = (x5 | ((~x3 | ~x4 | (x1 ? (x2 ^ x6) : (x2 | ~x6))) & (x1 | x3 | x4 | (~x2 ^ x6)))) & (x1 | x3 | ~x5 | x6 | (x2 ^ x4));
  assign n104 = (x2 | ((x1 | ((~x0 | x5 | (x3 & ~x4)) & (~x4 | ~x5 | (x0 & x3)))) & (x0 | ((~x1 | ((x4 | ~x5) & (x3 | ~x4 | x5))) & (~x3 | x4 | x5))))) & (x0 | ~x2 | (x1 ? ((x4 | x5) & (~x3 | ~x4 | ~x5)) : (~x4 | x5)));
  assign z07 = x2 ? ~n107 : ~n106;
  assign n106 = (~x0 & ((~x1 & ~x4 & (~x5 | (~x3 & ~x6))) | (x3 & x4 & (~x5 ^ x6)) | (~x3 & ~x5 & x6))) | (~x4 & ((~x1 & ~x5 & (~x3 | x6)) | (x0 & x3 & x5))) | (x0 & (x1 | (~x3 & x5 & x6))) | (x1 & ((x5 & x6) | (x4 & (x3 | ~x5))));
  assign n107 = (x0 | (x5 ? (x4 ? (x1 & (~x3 | x6)) : ~x1) : ((~x1 | (x3 ? ~x4 : x6)) & (x1 | (x3 ? (x4 | x6) : ~x6)) & (x3 | (~x4 ^ x6))))) & (x4 | x5 | x6 | ~x0 | x1 | x3);
  assign z08 = ~n111 | (~x1 & ~n109) | (~x0 & x1 & ~n110);
  assign n109 = x5 ? (((~x4 ^ ~x6) | (x0 ? (x2 | x3) : (~x2 | ~x3))) & (x0 | x2 | x4 | ~x6)) : (((~x0 ^ x2) | (x3 ? (x4 | ~x6) : (~x4 | x6))) & (x3 | ~x6 | (x0 ? (~x2 | x4) : (x2 | ~x4))));
  assign n110 = (~x6 | ((~x2 | x3 | (~x4 ^ x5)) & (x2 | ~x3 | ~x4 | x5))) & (x2 | ~x3 | x6 | (~x4 ^ ~x5));
  assign n111 = (x0 | (x2 ? ((~x1 | ((x4 | x6) & (~x3 | ~x4 | ~x6))) & (x3 | x4 | x6) & (x1 | ~x4 | (~x3 ^ x6))) : (x1 ? ((x4 | ~x6) & (x3 | ~x4 | x6)) : (~x3 | (x4 ^ x6))))) & (~x3 | ~x4 | x6 | ~x0 | x1 | x2);
  assign z09 = ~n115 | (n75 & ~n113) | (~x1 & ~n114);
  assign n113 = x6 ? ((x3 ^ x5) | (x2 ^ x4)) : ((~x2 | x3 | ~x5) & (x2 | ~x3 | x4 | x5));
  assign n114 = x2 ? ((x0 | ((~x4 | (x3 ? (~x5 ^ x6) : (x5 | x6))) & (~x5 | ~x6 | x3 | x4))) & (x4 | ~x5 | x6 | ~x0 | x3)) : (x5 ? (x6 | ((~x3 | x4) & (x0 | x3 | ~x4))) : (x0 ? (x3 ? ~x6 : (x4 | x6)) : (x4 | ~x6)));
  assign n115 = ((~x3 ^ ~x5) | ((x1 | x2 | ~x4) & (x0 | ~x1 | ~x2 | x4))) & (x0 | ((~x1 | x2 | (x3 ? (~x4 | x5) : ~x5)) & (x1 | ~x2 | ~x3 | x4 | x5)));
  assign z10 = n118 | n119 | n120 | n122 | (~x3 & ~n117);
  assign n117 = (x4 | (x0 ? (x1 | (x2 ? (x5 | ~x6) : (~x5 | x6))) : (~x2 | ((~x5 | x6) & (~x1 | x5 | ~x6))))) & (x0 | ~x4 | ((x1 | ~x5 | x6) & (x2 | x5 | ~x6)));
  assign n118 = ~x1 & ((~x0 & ((~x2 & ~x3 & ~x4 & x6) | (x3 & (x2 ? (x4 ^ x6) : (x4 & x6))))) | (~x2 & ((x3 & ~x4 & ~x6) | (x4 & x6 & x0 & ~x3))));
  assign n119 = ~x0 & x1 & ((x2 & (x3 ? (~x4 & x6) : (x4 & ~x6))) | (~x2 & x3 & ~x4 & ~x6));
  assign n120 = ~n121 & ((~x2 & (~x3 ^ x4) & (x0 ^ x1)) | (~x0 & ~x1 & x2 & ~x3 & x4));
  assign n121 = x5 ^ x6;
  assign n122 = n123 & n75 & (x2 ? n125 : n124);
  assign n123 = x3 & x4;
  assign n124 = ~x5 & x6;
  assign n125 = x5 & ~x6;
  assign z11 = ~n128 | (n127 & (x0 ? (x2 & (~x5 | ~x6)) : (~x2 & (x5 | x6))));
  assign n127 = ~x4 & ~x1 & ~x3;
  assign n128 = (x0 & (x1 | x2)) | (~x0 & ~x1 & ~x2 & ~x3 & ~x4);
  assign z16 = ~n132 | (~x1 & ~n130) | (~x0 & x1 & ~n131);
  assign n130 = (x3 | (x0 ? ((x4 | ~x5 | x6) & (x5 | ~x6 | x2 | ~x4)) : (~x2 | (x4 ? (~x5 | x6) : (x5 ^ x6))))) & (x0 | ~x2 | ~x3 | x4 | x5 | ~x6);
  assign n131 = (x2 | ((x5 | ~x6 | ~x3 | x4) & (~x5 | x6 | x3 | ~x4))) & (~x3 | ~x4 | (x5 ^ x6));
  assign n132 = (x0 | ((x3 | ((~x4 | x5) & (~x1 | (x5 & (~x2 | ~x4))))) & (~x3 | x4 | ~x5) & (x1 | ((~x3 | ~x5) & (x2 | x4 | (~x3 & ~x5)))))) & (x1 | ((x2 | ((~x3 | x4 | ~x5) & (~x0 | ~x4 | (~x3 ^ x5)))) & (x4 | x5 | ~x0 | x3)));
  assign z17 = ~n136 | (x2 ? ~n134 : ~n135);
  assign n134 = (x0 | (x1 ? (x3 ? (~x4 | x6) : (x4 | ~x6)) : (x5 | (x3 ? (x4 | x6) : (~x4 | ~x6))))) & (x1 | x3 | x4 | ~x5 | x6);
  assign n135 = ((x5 ^ x6) | ((x0 | ~x1 | ~x3 | x4) & (x3 | ~x4 | ~x0 | x1))) & (x0 | ~x4 | ((~x1 | (x3 ? (~x5 | x6) : (x5 | ~x6))) & (~x5 | ~x6 | x1 | ~x3))) & (x1 | x4 | x5 | ~x6 | (~x0 & x3));
  assign n136 = (x1 | ((x2 | (x0 ? (x3 ? ~x4 : (x4 | ~x5)) : (~x4 | x5))) & (x0 | ((~x3 | (~x4 ^ x5)) & (x4 | x5 | ~x2 | x3))))) & (x0 | ((~x1 | x4 | (x2 ? (~x3 | x5) : x3)) & (~x4 | ((x3 | ~x5) & (x2 | ~x3 | x5)))));
  assign z18 = n140 | ~n142 | (~x0 & (~n138 | ~n139));
  assign n138 = (~x4 | (x1 ? ((~x2 | ~x3 | x5 | ~x6) & (x2 | x3 | ~x5 | x6)) : (x2 | ~x3 | (~x5 ^ x6)))) & (x1 | x4 | ((~x5 | ~x6 | x2 | x3) & (~x2 | ~x3 | (x5 ^ x6))));
  assign n139 = x1 ? ((~x2 | (x3 ? (~x4 ^ x6) : (x4 | x6))) & (x4 | ~x6 | x2 | x3)) : (~x6 | (x2 ? (~x3 | ~x4) : (~x3 ^ x4)));
  assign n140 = ~x4 & n141 & (x2 ? (~x3 & n124) : (x3 & ~n121));
  assign n141 = x0 & ~x1;
  assign n142 = (x1 | ((~x0 | x2 | (x3 ? (~x4 | ~x6) : x6)) & (x3 | x6 | x0 | ~x2))) & (x0 | ~x1 | (x2 ? (x3 | ~x6) : (~x3 | x6)));
  assign z19 = n145 | ~n146 | (~x3 & ~n144);
  assign n144 = (x4 | ((x0 | ((x1 | x2 | x5 | ~x6) & (~x1 | ~x2 | x6))) & (~x0 | x1 | ~x5 | x6))) & (x0 | ~x1 | ~x4 | (x2 ? (~x5 | ~x6) : (x5 | x6)));
  assign n145 = ~x1 & ~x5 & ((~x4 & (x0 ? (x2 ^ x3) : (x2 & x3))) | (x3 & x4 & ~x0 & ~x2));
  assign n146 = ~n148 & ~n147 & (x0 | ~x3 | ~x6 | n149);
  assign n147 = ~x0 & (x1 ? (x2 ? (x3 & ~x4) : (~x3 ^ x4)) : (x2 ? (~x3 & x4) : (x3 & ~x4)));
  assign n148 = x4 & ~x3 & ~x2 & x0 & ~x1;
  assign n149 = (~x1 | (x2 ? (~x4 | x5) : (x4 | ~x5))) & (x1 | ~x2 | ~x4 | ~x5);
  assign z20 = n152 | n153 | (x3 ? (~x0 & ~n154) : ~n151);
  assign n151 = (x4 | (((~x2 ^ x6) | (x0 ? (x1 | ~x5) : x5)) & (x0 | ~x1 | x2 | ~x6))) & (x0 | ((~x2 | ((~x4 | ~x5 | x6) & (~x1 | ((~x5 | x6) & (~x4 | x5 | ~x6))))) & (~x1 | x2 | ~x4 | x5 | x6)));
  assign n152 = ~x1 & ((~x2 & ((x0 & (~x4 ^ x5)) | (x4 & (x3 ^ x5)) | (~x0 & ((x4 & ~x5) | (x3 & ~x4 & x5))))) | (~x0 & x2 & ~x4 & (x3 ^ x5)));
  assign n153 = x5 & ~x4 & x3 & x2 & ~x0 & x1;
  assign n154 = (~x4 | ((~x2 | ((x5 | ~x6) & (x1 | ~x5 | x6))) & (~x5 | ~x6 | ~x1 | x2))) & (~x1 | x2 | x4 | (~x5 ^ x6));
  assign z21 = (~x1 & ((~x2 & x6) | (x0 & x2 & n156))) | ~n157 | (~x0 & x1 & ~x2 & ~x6);
  assign n156 = x6 & ~x5 & ~x3 & ~x4;
  assign n157 = x0 | ~x2 | ((~x1 | (~x3 ^ ~x6)) & (~x3 | x4 | ~x6) & (x1 | (x3 ? (~x4 | x6) : ~x6)));
  assign z22 = ~n161 | (~x1 & (~n159 | ~n160));
  assign n159 = (~x0 | x3 | ((x5 | ~x6 | x2 | ~x4) & (~x2 | x4 | ~x5 | x6))) & (~x4 | x5 | ~x6 | x0 | x2 | ~x3);
  assign n160 = x2 ? ((x3 | x4 | x5) & (x0 | (x3 & x4))) : ((~x3 | ~x4 | ~x5) & (~x0 | (~x3 & (~x4 | ~x5))));
  assign n161 = ~n162 & (x0 | ~x1 | x2 | ~n124 | ~n77);
  assign n162 = ~x0 & x1 & (x2 ? ~x3 : (x3 & (x4 | x5)));
  assign z23 = n166 | n167 | ~n168 | (~x1 & (~n164 | ~n165));
  assign n164 = (x3 | ((~x0 | x6 | (x2 ? (x4 | ~x5) : (~x4 | x5))) & (x0 | ~x2 | ~x4 | x5 | ~x6))) & (~x4 | x5 | x6 | x0 | x2 | ~x3);
  assign n165 = x0 ? (x2 | (~x3 ^ ~x4)) : (~x3 | x4);
  assign n166 = ~x0 & x5 & (x1 ? (x2 ? (x3 & x4) : (~x3 & ~x4)) : (~x3 & x4));
  assign n167 = x3 & ~x5 & n75 & (x2 ? (x4 & x6) : (~x4 & ~x6));
  assign n168 = x3 | ((x0 | ~x1 | (~x2 & ~x4)) & (~x0 | x1 | ~x2 | x4 | x5));
  assign z24 = (~x1 & ~n170) | (~x0 & x1 & ~n171);
  assign n170 = (~x5 & (x4 ? (x6 & (x0 | x2 | x3)) : ((~x2 & ~x3) | (~x0 & (~x2 | (~x3 & ~x6)))))) | (x5 & ((~x0 & ~x2 & (x4 | ~x6)) | (~x3 & x4) | (x0 & x2 & x6))) | (x3 & ((x0 & (x2 | (x4 & ~x6))) | (x2 & x4 & ~x6))) | (x0 & x2 & x4);
  assign n171 = (x3 | (x2 ? ~x4 : (x4 | x5))) & (~x2 | (x4 ? (x5 | x6) : (~x5 | ~x6))) & (x2 | (x4 ? (~x5 & (~x3 | ~x6)) : (x5 | x6)));
  assign z25 = n173 | ~n175 | n178 | n179 | (~x2 & ~n174);
  assign n173 = ~n90 & ((x0 & ~x1 & x2 & ~x3 & ~x4) | (~x0 & ((~x1 & (x2 ? (x3 & x4) : ~x4)) | (x1 & x2 & x3 & ~x4))));
  assign n174 = ((x3 ^ x5) | ((x0 | ~x1 | x4 | ~x6) & (~x0 | x1 | ~x4 | x6))) & (~x4 | ~x5 | ~x6 | x0 | ~x1 | x3);
  assign n175 = ~n176 & ~n177 & (x3 | ~n92 | ~n76);
  assign n176 = ~x0 & x2 & x5 & (x1 ? (~x3 & x4) : ~x4);
  assign n177 = ~x2 & (x3 ^ ~x5) & (x0 ? (~x1 & ~x4) : (x1 & x4));
  assign n178 = ~x0 & ~x5 & ~x6 & ((~x2 & x3) | (~x1 & x2 & ~x3));
  assign n179 = n94 & ((~x1 & ~x3 & x4 & x5 & x6) | (x1 & ~x4 & ~x6 & (~x3 ^ ~x5)));
  assign z26 = ~n183 | (x3 ? ~n182 : ~n181);
  assign n181 = (x0 | (x1 ? (((~x2 ^ x6) | (~x4 ^ x5)) & (x2 | x4 | x5 | x6)) : (x2 ? (~x6 | (x4 ^ x5)) : (x6 | (~x4 ^ x5))))) & (~x0 | x1 | x2 | x4 | x5 | ~x6);
  assign n182 = ((~x5 ^ x6) | ((x2 | ~x4 | ~x0 | x1) & (x0 | x4 | (x1 ^ x2)))) & (x0 | ~x4 | ((x1 | x2 | (x5 ^ x6)) & (~x5 | ~x6 | ~x1 | ~x2)));
  assign n183 = (x1 | (x4 ? ((x0 | (x2 ? x6 : (x3 | ~x6))) & (x3 | x6 | ~x0 | x2)) : ((~x0 | (x2 ? (x3 | x6) : (~x3 | ~x6))) & (~x3 | ~x6 | x0 | ~x2)))) & (x0 | ((~x1 | x2 | ~x3 | x4 | x6) & (~x4 | ((~x2 | ~x3 | x6) & (~x1 | ~x6 | (~x2 ^ x3))))));
  assign z27 = ~n187 | (x3 ? ~n185 : ~n186);
  assign n185 = (x6 | ((x0 | ((~x1 | x5 | (x2 & ~x4)) & (x4 | ~x5 | x1 | ~x2))) & (~x0 | x1 | x2 | x4 | ~x5))) & (~x4 | ~x5 | ~x6 | x0 | ~x1 | ~x2);
  assign n186 = (x1 | ((x2 | ((~x0 | ~x5 | (~x4 ^ x6)) & (x5 | ~x6 | x0 | ~x4))) & (x0 | ~x2 | ((~x5 | ~x6) & (x4 | x5 | x6))))) & (x0 | ~x1 | ~x6 | (x2 ? x5 : (~x4 | ~x5)));
  assign n187 = (x1 | ((x2 | ((~x0 | x5 | (x3 & x4)) & (~x3 | ~x5 | (x0 & ~x4)))) & (x0 | ((~x3 | ~x4 | ~x5) & (~x2 | x5 | (~x3 & ~x4)))))) & (x0 | ~x1 | ~x5 | (x2 ? (~x3 ^ x4) : (x3 | x4)));
  assign z28 = ~n191 | (~x1 & ~n189) | (~x0 & x1 & ~n190);
  assign n189 = ((~x3 ^ x4) | ((~x5 | ~x6 | ~x0 | x2) & (x0 | ~x2 | x5 | x6))) & (x0 | ((x2 | ((x4 | ~x5 | x6) & (x3 | x5 | ~x6))) & (~x5 | ~x6 | ~x2 | x4))) & (~x0 | x2 | ~x4 | x5 | x6);
  assign n190 = ((x3 ^ x6) | (x2 ? (~x4 | ~x5) : (x4 | x5))) & (x5 | ~x6 | ~x2 | x3) & (x2 | ~x3 | ~x4 | ~x5 | x6);
  assign n191 = x0 ? (x1 | x4 | (x2 ? (x3 | x5) : (~x3 ^ x5))) : (x1 ? (x2 ? (x4 | ~x5) : (~x4 | x5)) : (~x4 | ((~x2 | ~x3 | x5) & (~x5 | (x2 & x3)))));
  assign z29 = n195 | ~n196 | (~x1 & (~n193 | ~n194));
  assign n193 = (x0 | ~x2 | x3 | ~x4 | ~x5) & (x4 | ((x2 | ((~x3 | ~x5 | ~x6) & (~x0 | ((~x5 | ~x6) & (~x3 | x5 | x6))))) & (x0 | ~x2 | x3 | x5 | x6)));
  assign n194 = (x3 | (x0 ? ((x4 | x6) & (x2 | ~x4 | ~x6)) : (x4 | ~x6))) & (x0 | ((~x2 | x4 | ~x6) & (~x3 | x6 | (x2 & ~x4))));
  assign n195 = ~n90 & ((~x0 & ((~x3 & x4 & ~x1 & ~x2) | (x1 & ~x4 & (~x2 | ~x3)))) | (x0 & ~x1 & ~x2 & x3 & x4));
  assign n196 = ~n75 | ((~x2 | ((~x4 | x5) & (~x3 | x4 | x6))) & (~x4 | ((x2 | (x6 ? ~x5 : x3)) & (~x3 | x5) & (x3 | ~x5 | ~x6))));
  assign z30 = n199 | ~n200 | (~x0 & ~n198);
  assign n198 = (~x4 | ((~x1 | ((~x5 | ~x6 | ~x2 | ~x3) & (x2 | x3 | x5 | x6))) & (x5 | ~x6 | ~x2 | x3))) & (x1 | x4 | ((x2 | ~x6 | (x3 ^ x5)) & (~x2 | ~x3 | ~x5 | x6)));
  assign n199 = ~x2 & (x4 ? ((~x0 & (x3 | (~x1 & ~x5))) | (~x1 & x3 & ~x5)) : (((~x3 | x5) & (x0 ^ x1)) | (~x1 & ~x3 & x5)));
  assign n200 = (~x3 | ((~x4 | ~x5 | x6 | ~n76) & (x4 | x5 | ~n94))) & (x3 | ~x4 | ~x5 | ~n94);
  assign z31 = n203 | n204 | (x5 ? ~n205 : ~n202);
  assign n202 = (x0 | ((~x4 | ((~x2 | x3 | ~x6) & (~x1 | ((x3 | ~x6) & (x2 | ~x3 | x6))))) & (x1 | x2 | x4 | (~x3 ^ x6)))) & (x3 | x4 | x6 | ~x0 | x1 | ~x2);
  assign n203 = ~x1 & (x0 ? (~x2 & (x3 ? (~x4 & x5) : ~x5)) : (x3 ? (x4 & ~x5) : ((x4 & x5) | (x2 & ~x4 & ~x5))));
  assign n204 = ~x0 & x1 & (x3 ? (~x4 & x5) : ((~x4 & ~x5) | (~x2 & x4 & x5)));
  assign n205 = ((~x3 ^ ~x6) | ((x0 | (x1 ? (~x2 | ~x4) : x4)) & (~x0 | x1 | x2 | ~x4))) & (x3 | x4 | x6 | x0 | x2);
  assign z32 = n207 | ~n210 | (~x5 & ~n208) | (~n121 & ~n209);
  assign n207 = ~x0 & (x1 ? ((x4 & ~x5 & x6) | (x5 & ~x6 & x2 & ~x4)) : ((x4 & x5 & ~x6) | (~x2 & (x4 ^ x6))));
  assign n208 = (x0 | ((x1 | ~x2 | x3 | ~x6) & (~x1 | ~x3 | x4 | x6))) & (x1 | x3 | ~x6 | ((~x2 | x4) & (~x0 | x2 | ~x4)));
  assign n209 = (~x0 | x1 | x2 | ~x4) & (x0 | (x1 ? ((~x2 | ~x3 | ~x4) & (x3 | x4)) : (~x2 | x4)));
  assign n210 = ~x5 | ((x4 | x6 | ~n76) & (~n75 | n211));
  assign n211 = (x2 | ~x3 | x4 | x6) & (~x2 | x3 | ~x4 | ~x6);
  assign z33 = ~n215 | ~n219 | ((~x6 | (~x2 & ~n213)) & (~n214 | (~n213 & (x2 | x6))));
  assign n213 = (~x0 | x1 | x3 | x4 | ~x5) & (x0 | ((~x1 | ~x3 | (~x4 ^ x5)) & (x1 | x3 | x4 | x5)));
  assign n214 = (x0 | ((~x1 | x3 | ~x5 | (~x2 ^ x4)) & (x1 | ~x2 | ~x3 | ~x4 | x5))) & (~x3 | x4 | x5 | ~x0 | x1 | x2);
  assign n215 = ~n217 & ~n218 & (~x2 | ~n75 | ~n216);
  assign n216 = x5 & x6 & (x3 ^ x4);
  assign n217 = ~x0 & x1 & x3 & (x2 ? (x4 & x5) : (~x4 & ~x5));
  assign n218 = ~x6 & ~x5 & ~x3 & ~x2 & x0 & ~x1;
  assign n219 = ~n220 & ~n221;
  assign n220 = ~x1 & ((~x5 & (x0 ? (x2 ? (~x3 & ~x4) : (x3 & x4)) : (x2 & (x3 ^ x4)))) | (~x3 & x5 & ~x0 & ~x2));
  assign n221 = ~x0 & ((~x2 & ((x1 & (x3 ? (x5 & ~x6) : (~x5 & x6))) | (x5 & x6 & ~x1 & x3))) | (~x1 & x2 & ~x3 & x5 & x6));
  assign z34 = n224 | n225 | ~n226 | (~x1 & ~n223);
  assign n223 = (~x3 | ((x0 | ~x6 | (x2 ? (x4 ^ x5) : (~x4 | x5))) & (~x0 | x2 | x4 | x5 | x6))) & (~x2 | x3 | x6 | ((x4 | ~x5) & (x0 | ~x4 | x5)));
  assign n224 = ~x3 & ((~x2 & (~x5 ^ x6) & (x0 ^ x1)) | (~x0 & x2 & ((~x5 & x6) | (x1 & x5 & ~x6))));
  assign n225 = ~x0 & x3 & ~x6 & ((~x2 & x5) | (~x1 & x2 & ~x5));
  assign n226 = n228 & (~n75 | ~n227 | (x3 ? (x4 | ~x6) : (~x4 | x6)));
  assign n227 = ~x2 & x5;
  assign n228 = (~x0 | x1 | x2 | ~x3 | ~x5) & (x0 | ((x3 | ~x5 | x1 | x2) & (~x1 | ~x2 | ~x3 | x5)));
  assign z35 = n231 | n232 | (~x2 & ~n230) | (~n233 & n234);
  assign n230 = ((x3 ^ x6) | ((x4 | ~x5 | ~x0 | x1) & (~x4 | x5 | x0 | ~x1))) & (x1 | ~x3 | x4 | (x0 ? (x5 | x6) : (~x5 ^ x6)));
  assign n231 = ~x0 & ((~x3 & x6 & ((~x2 & x4) | (~x1 & (~x2 | x4)))) | (x4 & ~x6 & ~x1 & x3));
  assign n232 = (x3 ^ ~x6) & ((x0 & ~x1 & ~x2 & x4) | (~x0 & ((x2 & ~x4) | (x1 & (x2 | ~x4)))));
  assign n233 = x0 ^ ~x5;
  assign n234 = x6 & ~x4 & ~x3 & ~x1 & x2;
  assign z36 = n237 | ~n238 | (~x2 & ~n236);
  assign n236 = (x1 | ((~x0 | ((x3 | x4 | x5 | x6) & (~x5 | ~x6 | ~x3 | ~x4))) & (~x4 | x5 | ~x6 | x0 | x3))) & (x0 | ~x1 | ((~x5 | x6 | ~x3 | ~x4) & (x3 | x5 | (~x4 ^ x6))));
  assign n237 = ~x1 & ((~x0 & (x2 ? (x3 & ~x4) : (x4 & x5))) | (~x4 & ~x5 & x2 & ~x3) | (~x2 & (x3 ? (~x4 & ~x5) : (x4 & x5))));
  assign n238 = (~x2 | ((~x4 | ~n75) & (x3 | x4 | ~x5 | n239))) & (~n75 | ((x2 | x4 | ~x5) & (~x3 | ~x4 | x5)));
  assign n239 = (x1 | x6) & (x0 | ~x1 | ~x6);
  assign z37 = n242 | n243 | ~n245 | (~x0 & ~n241);
  assign n241 = x2 ? (~x4 | ~x5 | ~x6 | (x1 & ~x3)) : ((~x5 | ~x6 | x3 | x4) & (x5 | x6 | ((x3 | ~x4) & (~x1 | (x3 & ~x4)))));
  assign n242 = ~x0 & x3 & ((~x2 & ~x4 & ~x5) | (~x1 & (x2 ? (~x4 & x5) : ~x5)));
  assign n243 = ~n90 & (x0 ? (~x1 & ~n244) : (x1 ? ~n244 : (x2 & ~x3)));
  assign n244 = x2 ? (x3 | x4) : (~x3 | ~x4);
  assign n245 = x3 ? (x4 | n246) : ((~x4 | n246) & (x6 | ~n76 | x4 | x5));
  assign n246 = (x0 | ~x1 | ~x2 | ~x5) & (~x0 | x1 | x2 | x5);
  assign z38 = n249 | n250 | n251 | (~x2 & ~n248);
  assign n248 = (x1 | ((x4 | ((~x0 | ~x6 | (~x3 ^ x5)) & (~x5 | x6 | x0 | x3))) & (~x4 | x5 | ~x6 | x0 | ~x3))) & (x0 | ~x4 | ((x3 | (x5 ^ x6)) & (~x1 | ~x3 | ~x5 | x6)));
  assign n249 = ~x1 & (x0 ? ((~x3 & ~x4 & ~x6) | (~x2 & x4 & (x3 ^ x6))) : ((x3 & ~x4 & x6) | (x2 & ~x3 & ~x6)));
  assign n250 = ~x0 & x1 & (x3 ? (~x4 & x6) : ((~x4 & ~x6) | (x2 & x4 & x6)));
  assign n251 = x4 & x5 & n94 & ((x3 & ~x6) | (~x1 & ~x3 & x6));
  assign z39 = n254 | (x2 ? (~x0 & ~n256) : (~n253 | ~n255));
  assign n253 = (x0 | ((x1 | ~x3 | x4 | ~x5 | ~x6) & (x5 | ((~x1 | (x3 ? (~x4 | ~x6) : x4)) & (x4 | x6 | x1 | ~x3))))) & (x1 | x3 | ~x4 | ~x5 | (~x0 & x6));
  assign n254 = ~x0 & x2 & ((x4 & (x1 ? (x5 ^ x6) : (x5 & x6))) | (~x1 & ~x4 & ~x5 & ~x6));
  assign n255 = (x1 | (x0 ? (x4 ? x5 : (~x5 | ~x6)) : (x4 | (~x5 ^ x6)))) & (x0 | ~x4 | ~x5 | (~x1 & ~x6));
  assign n256 = x1 ? (x3 | ((~x4 | ~x5 | ~x6) & (x5 | x6))) : (~x3 | ((x5 | ~x6) & (~x4 | ~x5 | x6)));
  assign z40 = ~n260 | (~x0 & (~n258 | ~n259));
  assign n258 = (~x3 | (((~x1 ^ ~x2) | (x4 ? (~x5 | ~x6) : (x5 | x6))) & (x1 | ~x2 | x4 | ~x5 | ~x6))) & (x1 | x2 | x3 | x4 | ~x5 | ~x6);
  assign n259 = x1 ? (x6 | (x2 ? (x3 | ~x4) : (~x3 | x4))) : (x2 ? (x3 ? (~x4 | ~x6) : x4) : (x3 | ~x4));
  assign n260 = ~n261 & ~n262 & ~n263 & (~n92 | ~n76 | ~n77);
  assign n261 = ~x6 & ((~x0 & x5 & (x1 ? (~x2 & ~x3) : (x2 & x3))) | (x0 & ~x1 & ~x2 & ~x3 & ~x5));
  assign n262 = x0 & ~x1 & ~x2 & (x3 ? x4 : (~x4 & x6));
  assign n263 = ~x0 & x1 & ~x5 & x6 & (x2 ^ x3);
  assign z41 = (~x0 & (~n265 | ~n267)) | ~n268 | (~n121 & ~n266);
  assign n265 = ((~x3 ^ x5) | ((~x1 | x2 | ~x4 | x6) & (x1 | ~x2 | (~x4 ^ ~x6)))) & (x4 | ~x6 | ((~x3 | (x1 ? (x2 ^ ~x5) : (x2 | x5))) & (x1 | ~x2 | x3 | x5)));
  assign n266 = (x0 | ((~x1 | x3 | (x2 ^ x4)) & (x1 | x2 | ~x3 | ~x4))) & (~x0 | x1 | x2 | ~x3 | x4);
  assign n267 = (~x3 | ((~x1 | x2 | (x4 ^ x5)) & (x4 | ~x5 | x1 | ~x2))) & (x1 | ~x2 | x3 | ~x4 | x5);
  assign n268 = ~n270 & ~n271 & ~n273 & (n269 | n272);
  assign n269 = x3 ? (~x5 | x6) : (x5 | ~x6);
  assign n270 = ~x5 & ~x4 & ~x3 & x2 & x0 & ~x1;
  assign n271 = ~x0 & ((~x1 & ~x2 & ~x3 & (x4 ^ x6)) | (x1 & x2 & x3 & x4 & x6));
  assign n272 = (x0 | ~x1 | ~x2 | x4) & (x2 | ~x4 | ~x0 | x1);
  assign n273 = ~x6 & ~x4 & ~x3 & ~x2 & x0 & ~x1;
  assign z42 = ~n277 | (~x1 & ~n275) | (~x0 & x1 & ~n276);
  assign n275 = (x0 | (x6 ? (x3 ? (~x4 | x5) : (~x5 | (x2 & ~x4))) : ((~x3 | x4 | ~x5) & (~x2 | (x3 ? ~x5 : (x4 | x5)))))) & (x2 | ((~x0 | ((x3 | ~x5 | x6) & (~x4 | (x3 ? (x5 ^ x6) : (x5 | ~x6))))) & (x3 | ~x4 | ~x5 | x6) & (x5 | ~x6 | ~x3 | x4)));
  assign n276 = x3 ? (x2 ? (x4 ? (~x5 | ~x6) : (x5 | x6)) : (~x5 | (~x4 ^ x6))) : ((x4 | ((x5 | ~x6) & (~x2 | ~x5 | x6))) & (x5 | x6 | (x2 & ~x4)));
  assign n277 = (x3 | ((x1 | ((x4 | (x0 ? (~x2 ^ x6) : (~x2 | ~x6))) & (~x4 | x6 | x0 | ~x2))) & (x0 | ~x1 | ~x2 | ~x4 | ~x6))) & (x0 | ~x1 | ~x3 | x4 | (x2 ^ x6));
  assign z43 = ~n281 | (~x2 & ~n279) | (~x0 & x2 & ~n280);
  assign n279 = (x0 | ((x5 | x6 | ~x3 | x4) & (~x6 | ((~x1 | ~x3 | ~x4 | x5) & ((x3 & ~x5) | (x1 ^ ~x4)))))) & (x1 | ((~x4 | x6 | ((~x3 | x5) & (~x0 | (~x3 & x5)))) & (~x0 | ~x3 | x4 | ~x5 | ~x6)));
  assign n280 = (~x1 | x3 | (x4 ? (x5 | ~x6) : x6)) & (~x3 | ((x4 | (~x5 ^ x6)) & (x1 | ~x5 | x6)));
  assign n281 = (x1 | (x2 ? (x3 | x5 | (x0 & x4)) : (x0 ? (x3 ? (x4 | x5) : ~x5) : (x4 | ~x5)))) & (x0 | ~x1 | ~x4 | ~x5 | (~x2 ^ ~x3));
  assign z44 = n284 | n287 | n288 | (~x1 & (~n283 | ~n286));
  assign n283 = (x2 | (((~x4 ^ x5) | (~x0 ^ ~x6)) & (~x0 | ~x3 | x4 | x5 | x6))) & (x0 | x3 | (x4 ? ((x5 | x6) & (~x2 | ~x5 | ~x6)) : (~x5 | x6)));
  assign n284 = ~n285 & (x4 ^ ~x5);
  assign n285 = (~x0 | x1 | x2 | x3 | x6) & (x0 | ((~x1 | (x2 ? (~x3 | x6) : (x3 | ~x6))) & (~x3 | ~x6 | x1 | ~x2)));
  assign n286 = (x0 | ~x4 | (x2 ? (~x3 | x6) : ~x6)) & (~x0 | ~x2 | x3 | x4 | x6);
  assign n287 = ~x0 & x1 & ((~x2 & x4 & ~x6) | (~x4 & x6 & (x2 | x3)));
  assign n288 = n125 & x4 & ~x3 & x2 & ~x0 & x1;
  assign z45 = n291 | ~n293 | (~x0 & (~n290 | ~n292));
  assign n290 = x2 ? ((~x1 | (~x3 & ~x4) | (~x5 ^ x6)) & (~x5 | ~x6 | x1 | ~x3)) : ((x3 | (x1 ? (x5 ^ x6) : ((x5 | ~x6) & (~x4 | ~x5 | x6)))) & (x1 | x4 | ((x5 | ~x6) & (~x3 | ~x5 | x6))));
  assign n291 = ~n244 & ((~x1 & (x0 ? (~x5 & ~x6) : x5)) | (~x0 & ~x5 & (x1 | x6)));
  assign n292 = (~x1 | x2 | ~x3 | x4 | x5) & (x1 | ~x2 | x3 | ~x4 | ~x5);
  assign n293 = (~n141 | ~n227 | (x3 & x4)) & (~n92 | ~n76 | ~x3 | ~x4);
  assign z46 = n296 | ~n298 | (x1 ? (~x0 & ~n297) : ~n295);
  assign n295 = (x4 | ((x5 | ~x6 | ~x2 | x3) & (~x5 | ((x0 | (x2 ? (~x3 | ~x6) : x3)) & (~x0 | x2 | ~x3 | ~x6))))) & (x0 | ~x3 | x5 | (x2 ? x6 : (~x4 | ~x6)));
  assign n296 = ~x0 & ((~x1 & x6 & (x2 ? (x3 & x4) : (x3 ^ x4))) | (x1 & ~x2 & x3 & x4 & ~x6));
  assign n297 = (~x2 | x3 | x4 | x5 | ~x6) & (x2 | ~x5 | x6 | (x3 ^ ~x4));
  assign n298 = x6 ? ((x2 | ((x0 | ~x1 | x3) & (~x3 | ~x4 | ~x0 | x1))) & (x0 | ~x1 | (x3 ? ~x2 : ~x4))) : ((x1 | (x0 ? (x2 | (x3 & x4)) : (~x2 | x3))) & (x3 | x4 | x0 | ~x2));
  assign z47 = n301 | ~n302 | (~x0 & ~n300);
  assign n300 = (x5 | ((~x2 | ((x4 | x6 | ~x1 | x3) & (x1 | (x6 ? x4 : ~x3)))) & (x6 | ((~x3 | ~x4) & (~x1 | x2 | (~x3 & ~x4)))))) & (~x5 | ~x6 | ~x1 | x4) & (x2 | ((~x3 | ((x4 | ~x5 | ~x6) & (~x1 | ~x4 | x6))) & (~x1 | ~x6 | (~x5 & (x3 | x4)))));
  assign n301 = ~n90 & ((~x1 & ((~x3 & (x0 ? (x2 ^ x4) : (x2 & x4))) | (~x2 & ((x3 & ~x4) | (~x0 & (x3 | ~x4)))))) | (x2 & x3 & x4 & ~x0 & x1));
  assign n302 = x4 ? (~x6 | n303) : (x6 | (n303 & (~x3 | x5 | ~n76)));
  assign n303 = (~x0 | x1 | x2 | x3 | ~x5) & (x0 | ~x1 | (x2 ? ~x5 : (x3 | x5)));
  assign z48 = ~n307 | (~x2 & ~n305) | (~x0 & x2 & ~n306);
  assign n305 = x0 ? (x1 | ((x3 | ~x6 | (x4 ^ x5)) & (x6 | ((~x4 | x5) & (~x3 | x4 | ~x5))))) : (((~x4 ^ x6) | (x1 ? (x3 | x5) : (~x3 | ~x5))) & (x3 | x4 | ~x5 | x6) & (x5 | ((~x3 | ~x4 | ~x6) & (x1 | ((~x4 | ~x6) & (~x3 | x4 | x6))))));
  assign n306 = ((~x4 ^ x6) | (x1 ? (x3 | ~x5) : (~x3 | x5))) & (~x4 | ~x5 | ~x6 | (x1 & ~x3)) & (x4 | x5 | x6 | (~x1 & x3));
  assign n307 = (x1 | (x0 ? ((x4 | x6 | ~x2 | x3) & (x2 | ~x3 | ~x4 | ~x6)) : (~x2 | x3 | (~x4 ^ x6)))) & (x0 | ~x1 | ((~x3 | (x2 ? (~x4 ^ x6) : (x4 | x6))) & (~x4 | ~x6 | x2 | x3)));
  assign z49 = n310 | n311 | n312 | ~n313 | (~x0 & ~n309);
  assign n309 = x1 ? ((x2 | x3 | x4 | ~x5 | x6) & (~x2 | ((~x3 | ~x6 | (x4 ^ x5)) & (x3 | x4 | x5 | x6)))) : ((x2 | ((x3 | x4 | x5 | ~x6) & (~x3 | x6 | (x4 ^ x5)))) & (~x2 | x3 | ~x4 | ~x5 | ~x6));
  assign n310 = ~n121 & ((x0 & ~x1 & ~x2 & ~x3 & ~x4) | (~x0 & ((~x1 & (x2 ? (x3 & ~x4) : (~x3 & x4))) | (x3 & x4 & x1 & ~x2))));
  assign n311 = ~x1 & ((~x3 & ((x4 & ~x5 & ~x0 & x2) | (x0 & (x2 ? (~x4 & ~x5) : (x4 & x5))))) | (~x0 & x3 & x5 & (~x2 ^ x4)));
  assign n312 = ~n90 & ((x0 & ~x1 & ~x2 & x3 & ~x4) | (~x0 & ~x3 & (x1 ? x4 : (x2 & ~x4))));
  assign n313 = ~n314 & (~n123 | ~n124 | ~n76);
  assign n314 = ~x0 & x1 & ((~x2 & x3 & ~x4 & ~x5) | (x2 & (x3 ? (x4 & ~x5) : (~x4 & x5))));
  assign z50 = ~n317 | (x3 ? ~n316 : ~n181);
  assign n316 = ((~x5 ^ x6) | ((x2 | ~x4 | ~x0 | x1) & (x0 | x4 | (x1 ^ x2)))) & (x0 | ~x4 | (x5 ^ x6) | (x1 ^ x2));
  assign n317 = (x1 | (x4 ? ((x0 | (x2 ? x6 : (x3 | ~x6))) & (x3 | x6 | ~x0 | x2)) : ((~x0 | (x2 ? (x3 | x6) : (~x3 | ~x6))) & (~x3 | ~x6 | x0 | ~x2)))) & (x0 | ~x1 | ((x2 | ~x3 | (x4 ^ x6)) & (~x4 | ~x6 | ~x2 | x3)));
  assign z51 = ~n321 | (~x1 & ~n319) | (~x0 & x1 & ~n320);
  assign n319 = (~x5 | (((~x3 ^ x6) | (x0 ? (x2 | x4) : ~x2)) & (~x0 | x2 | x3 | ~x4 | x6))) & (x0 | x3 | x5 | (x2 ? (x4 | x6) : (~x4 | ~x6)));
  assign n320 = (x2 | ((~x3 | x5 | x6) & (~x5 | ~x6 | x3 | ~x4))) & (x5 | ((~x3 | ~x4 | x6) & (~x2 | x3 | ~x6)));
  assign n321 = (x1 | ((x2 | ((~x0 | x5 | (x3 & x4)) & (~x3 | ~x5 | (x0 & ~x4)))) & (x0 | ~x2 | x5 | (~x3 & ~x4)))) & (x0 | ~x1 | ~x5 | (~x2 ^ (~x3 & ~x4)));
  assign z52 = ~n325 | (~x1 & ~n323) | (~x0 & x1 & ~n324);
  assign n323 = x0 ? (x2 | ((~x3 | ((x5 | x6) & (x4 | ~x5 | ~x6))) & (~x4 | ((x5 | x6) & (x3 | ~x5 | ~x6))))) : (x2 ? ((~x3 | ((~x5 | ~x6) & (x4 | x5 | x6))) & (x3 | ~x4 | x5 | x6) & (x4 | ~x5 | ~x6)) : ((x4 | ~x5 | x6) & (x3 | x5 | ~x6)));
  assign n324 = (x3 | ((~x2 | (~x5 ^ x6)) & (x5 | x6 | x2 | x4))) & (x2 | ~x3 | (x4 ? (~x5 | x6) : (x5 | ~x6)));
  assign n325 = (x1 | ((x3 | (x0 ? (x4 | (~x2 ^ x5)) : (~x4 | ~x5))) & (x0 | ~x4 | (x2 ? (~x3 | x5) : ~x5)))) & (x0 | ~x1 | (x2 ? (~x3 | ~x5) : (~x4 | x5)));
  assign z53 = ~n329 | (~x2 & ~n327) | (~x0 & x2 & ~n328);
  assign n327 = (x1 | ((~x5 | (x0 ? (x3 ? (~x4 | x6) : (x4 | ~x6)) : (x3 ? (x4 | ~x6) : (~x4 | x6)))) & (~x4 | x5 | ~x6 | (x0 ^ x3)))) & (x0 | ~x1 | ((x3 | ~x6 | (x4 ^ x5)) & (x6 | ((x4 | ~x5) & (~x3 | ~x4 | x5)))));
  assign n328 = (~x1 | x3 | x4 | ~x5 | x6) & (x1 | ((~x4 | ~x5 | ~x6) & (x3 | (x4 ? ~x5 : (x5 | x6)))));
  assign n329 = (x1 | ((x2 | (x0 ? (~x6 | (~x3 ^ x4)) : (~x3 | x6))) & (x4 | (x0 ? (x3 | x6) : (~x6 | (~x2 & x3)))))) & (x0 | ((~x4 | x6 | ~x2 | ~x3) & (~x1 | (x2 ? (~x3 ^ x6) : (~x4 | (~x3 ^ ~x6))))));
  assign z54 = ~n333 | n331 | (~x0 & x6 & ~n332);
  assign n331 = ~x1 & ((~x2 & ((~x5 & (x0 ? (~x3 ^ x4) : (~x3 & x4))) | (~x4 & x5 & ~x0 & ~x3))) | (~x0 & x2 & (x3 ? (~x4 & ~x5) : (x4 & x5))));
  assign n332 = x2 ? (x1 ? (x3 ? (~x4 | x5) : (x4 | ~x5)) : (~x4 | (x3 ^ x5))) : (x4 | (x1 ? (~x3 | x5) : (x3 ^ x5)));
  assign n333 = n266 & ~n335 & (~n334 | ~n76);
  assign n334 = ~x6 & x5 & ~x3 & ~x4;
  assign n335 = ~x0 & x1 & x3 & (x2 ? (x4 & x5) : (x4 ^ x5));
  assign z55 = ~n339 | (~x1 & ~n337) | (~x0 & x1 & ~n338);
  assign n337 = x3 ? (~x5 | ((x0 | ~x6 | (x2 ^ x4)) & (~x0 | x2 | x4 | x6))) : ((x4 | ((x0 | ~x2 | x5 | x6) & (x2 | (x0 ? (x5 ^ x6) : (x5 | ~x6))))) & (x0 | ~x4 | ((~x5 | x6) & (~x2 | x5 | ~x6))));
  assign n338 = (~x6 | ((x2 | ~x3 | x4 | x5) & (~x2 | (x3 ? (~x4 | x5) : (x4 | ~x5))))) & (~x4 | x6 | ((x2 | ~x3 | x5) & (x3 | ~x5)));
  assign n339 = x0 ? (x1 | x2 | (x3 ? (x4 ^ x5) : (~x4 | x5))) : ((~x1 | (~x3 ^ ~x5)) & (~x2 | x4 | (x5 ? ~x3 : ~x1)));
  assign z56 = n342 | ~n345 | ~n346 | (~x0 & (~n341 | ~n344));
  assign n341 = (x1 | ((x6 | ((~x2 | (x3 ? (~x4 | x5) : (x4 | ~x5))) & (x4 | x5 | x2 | ~x3))) & (x2 | ~x5 | ~x6 | (~x3 ^ x4)))) & (x4 | x5 | ~x6 | ~x1 | x2 | ~x3);
  assign n342 = ~n343 & (x3 ^ ~x5);
  assign n343 = (~x0 | x1 | x2 | x4 | ~x6) & (x0 | ((~x1 | x6 | (~x2 ^ ~x4)) & (~x4 | ~x6 | x1 | ~x2)));
  assign n344 = (x1 | ((x2 | (x3 ? (~x4 | x5) : (x4 | ~x5))) & (~x4 | ~x5 | ~x2 | x3))) & ((x3 ^ x5) | (x1 ? (x2 | ~x4) : (~x2 | x4)));
  assign n345 = ~x0 | x1 | x3 | (x2 ? (x4 | x5) : ~x5);
  assign n346 = (~x3 | x5 | x6 | ~x0 | x1 | x2) & (x0 | ~x1 | ~x2 | (x3 ? x5 : (~x5 | ~x6)));
  assign z57 = ~n350 | (~x2 & ~n348) | (~x0 & x2 & ~n349);
  assign n348 = ((~x0 ^ x1) | ((x3 | x4 | x5 | ~x6) & (~x5 | x6 | ~x3 | ~x4))) & (~x4 | ((x0 | x3 | ((~x5 | ~x6) & (x1 | x5 | x6))) & (~x0 | x1 | ~x3 | x5 | ~x6))) & (x4 | ~x5 | x6 | x0 | x3);
  assign n349 = (x3 | x5 | ((x4 | x6) & (x1 | ~x4 | ~x6))) & (~x1 | ((x3 | x4 | ~x5 | ~x6) & (~x3 | ~x4 | x5 | x6)));
  assign n350 = (x1 | ((x3 | ((~x0 | x6 | (~x2 ^ x4)) & (x4 | ~x6 | x0 | ~x2))) & (x2 | ~x3 | ((x4 | ~x6) & (x0 | ~x4 | x6))))) & (x0 | ((~x4 | ((~x2 | ~x3 | ~x6) & (~x1 | (x2 ? ~x6 : (x3 | x6))))) & (~x3 | x4 | (~x2 ^ x6))));
  assign z12 = z11;
  assign z13 = z11;
  assign z14 = z11;
  assign z15 = z11;
  assign z59 = z58;
  assign z60 = z58;
  assign z61 = z58;
  assign z62 = z58;
  assign z63 = z58;
  assign z64 = z58;
endmodule


