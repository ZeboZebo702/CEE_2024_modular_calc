module x_100_mod_997_reg(
    input [100:1] X,
    output [10:1] R
    );


assign R = X % 997;

endmodule
