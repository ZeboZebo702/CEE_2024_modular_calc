// Benchmark "32_32_mod" written by ABC on Thu Dec 01 00:27:41 2022

module const_32_32_mod ( 
    x0, x1, x2, x3, x4, x5, x6,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63, z64  );
  input  x0, x1, x2, x3, x4, x5, x6;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63, z64;
  wire n74, n75, n76, n77, n78, n80, n81, n82, n83, n84, n85, n86, n88, n89,
    n90, n91, n92, n93, n94, n95, n96, n98, n99, n100, n101, n102, n103,
    n104, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
    n118, n119, n120, n121, n122, n124, n125, n126, n127, n128, n129, n131,
    n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143, n144,
    n145, n147, n148, n149, n150, n151, n152, n153, n154, n156, n157, n158,
    n159, n160, n161, n162, n163, n165, n166, n167, n169, n170, n171, n172,
    n173, n174, n175, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n188, n189, n190, n191, n192, n193, n194, n195, n196, n198, n199,
    n200, n201, n202, n203, n204, n205, n206, n207, n208, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n221, n222, n223, n224, n225,
    n226, n228, n229, n230, n231, n232, n233, n234, n236, n237, n238, n239,
    n240, n241, n242, n243, n244, n245, n246, n248, n249, n250, n251, n252,
    n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
    n266, n268, n269, n270, n271, n272, n273, n274, n275, n277, n278, n279,
    n280, n281, n282, n283, n284, n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n298, n299, n300, n301, n302, n303, n304, n306,
    n307, n308, n309, n310, n311, n313, n314, n315, n316, n317, n318, n319,
    n320, n321, n322, n324, n325, n326, n327, n328, n329, n330, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n343, n344, n345, n346,
    n347, n348, n349, n350, n352, n353, n354, n355, n356, n357, n358, n360,
    n361, n362, n363, n364, n365, n366, n367, n369, n370, n371, n372, n373,
    n374, n375, n377, n378, n379, n380, n381, n382, n384, n385, n386, n387,
    n388, n389, n391, n392, n393, n394, n395, n396, n397, n398, n399, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n413, n414,
    n415, n416, n417, n418, n420, n421, n422, n423, n424, n425, n427, n428,
    n429, n430, n431, n432, n433, n434, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n447, n448, n449, n450, n451, n452, n453, n454,
    n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n467, n468,
    n469, n470, n471, n472, n474, n475, n476, n477, n478, n479, n480, n481,
    n482, n484, n485, n487, n488, n489, n490, n491, n492, n494, n495, n496,
    n497, n498, n499, n500, n502, n503, n504, n505, n506, n507, n508, n510,
    n511, n512, n513, n514, n516, n517, n518, n519, n520, n521, n522, n524,
    n525, n526, n527, n528, n529, n530, n531, n533, n534, n535, n536, n537,
    n538;
  assign z58 = 1'b0;
  assign z00 = (~n74 & n75) | (n76 & n77 & n78);
  assign n74 = (~x2 | ((~x3 | ~x4 | x5 | ~x6) & (x3 | x4 | ~x5 | x6))) & (~x4 | ~x5 | ~x6 | x2 | x3);
  assign n75 = ~x0 & x1;
  assign n76 = ~x2 & x0 & ~x1;
  assign n77 = x3 & ~x4;
  assign n78 = ~x5 & ~x6;
  assign z01 = ~n83 | (~x1 & ~n80);
  assign n80 = (n81 | (~x3 ^ x6)) & (x4 | n82);
  assign n81 = (x0 | (x2 ? (~x4 | ~x5) : (x4 | x5))) & (~x0 | x2 | x4 | ~x5);
  assign n82 = (x5 | ((~x0 | (x2 ? (x3 | x6) : (~x3 | ~x6))) & (x0 | ~x2 | x3 | ~x6))) & (x0 | x2 | x3 | ~x5 | x6);
  assign n83 = x1 ? (x0 | (n85 & n86)) : n84;
  assign n84 = (~x4 | ((x2 | (x0 ? (x3 ^ x5) : (x3 | ~x5))) & (x0 | ~x3 | x5))) & (x0 | ~x2 | (x3 ? x5 : (x4 | ~x5)));
  assign n85 = (~x3 | (x4 ^ x5)) & (x2 | x3 | x4 | ~x5);
  assign n86 = (~x2 | x4 | ~x5 | (~x3 ^ x6)) & (~x4 | x5 | ((x3 | x6) & (x2 | ~x3 | ~x6)));
  assign z02 = n88 | (n75 & ~n96);
  assign n88 = ~x1 & (n90 | ~n91 | (x6 & ~n89));
  assign n89 = (x0 | ((x4 | ~x5 | x2 | x3) & (~x2 | ~x3 | ~x4 | x5))) & (~x2 | x3 | x4 | x5) & (~x3 | ~x4 | ~x5 | ~x0 | x2);
  assign n90 = ~x2 & (x4 ? ((x5 & ~x6) | (~x0 & (x5 | ~x6))) : (x6 & (x0 | ~x5)));
  assign n91 = ~n95 & ((~n92 & ~n93) | ~n78 | ~n94);
  assign n92 = x3 & x4;
  assign n93 = ~x3 & ~x4;
  assign n94 = x0 & ~x2;
  assign n95 = ~x0 & x2 & (x4 ? (~x5 ^ x6) : (x5 & ~x6));
  assign n96 = (x2 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (~x4 | ((x3 | x5 | ~x6) & (~x2 | ~x5 | x6))) & (x4 | ((~x2 | (x5 ^ x6)) & (~x3 | x5 | x6)));
  assign z03 = ~n100 | (~x0 & (x3 ? ~n99 : ~n98));
  assign n98 = x2 ? (~x4 | ((x5 | x6) & (x1 | ~x5 | ~x6))) : (x4 | ((~x5 | ~x6) & (~x1 | x5 | x6)));
  assign n99 = (~x1 | (x2 ? (~x6 | (x4 ^ x5)) : (x4 | ~x5))) & (x1 | x2 | ~x4 | x5 | x6);
  assign n100 = n103 & (x1 ? (x0 | n102) : n101);
  assign n101 = ((x5 ^ x6) | (x0 ? (x2 | x3) : (~x2 | ~x3))) & (x0 | x3 | (x2 ? (x5 | ~x6) : (~x5 | x6))) & (~x0 | x2 | ~x3 | ~x5 | x6);
  assign n102 = (~x2 | x5 | (x3 ^ ~x6)) & (x2 | x3 | ~x5 | x6);
  assign n103 = x5 ? (x6 ? (~n76 | ~n77) : n104) : (~x6 | n104);
  assign n104 = (x0 | x2 | ~x3 | (x1 & ~x4)) & (~x0 | x1 | ~x2 | x3 | x4);
  assign z04 = n107 | n109 | n112 | (~x0 & ~n106);
  assign n106 = (~x6 | (x1 ? ((~x3 | x4) & (~x2 | x3 | ~x4)) : (x3 | x4))) & (x1 | ~x3 | x6 | (~x2 & x4));
  assign n107 = n108 & ((~x3 & ~x4 & ~x6) | (~x2 & (x3 ? (~x4 & x6) : ~x6)));
  assign n108 = x0 & ~x1;
  assign n109 = ~x2 & ((n93 & ~n111) | (x4 & ~n110));
  assign n110 = x5 ? (x6 | ((x1 | ~x3) & (x0 | (x1 & ~x3)))) : (~x6 | (x0 ? (x1 | ~x3) : x3));
  assign n111 = (x0 | ~x1 | (x5 ^ x6)) & (~x0 | x1 | ~x5 | ~x6);
  assign n112 = n114 & (n115 | (x4 & n113 & n116));
  assign n113 = x5 & ~x6;
  assign n114 = ~x0 & x2;
  assign n115 = ~x3 & ((~x4 & ((~x5 & ~x6) | (x1 & x5 & x6))) | (~x5 & x6 & ~x1 & x4));
  assign n116 = x1 & x3;
  assign z05 = ~n122 | (n118 & ~n119) | (~n120 & n121);
  assign n118 = ~x0 & ~x2;
  assign n119 = (x1 | (x3 ? (~x4 | ~x5) : (~x4 ^ x5))) & (~x1 | x3 | x4 | x5);
  assign n120 = (x1 | x2 | ~x6 | (x3 ^ x4)) & (~x1 | ~x2 | ~x3 | ~x4 | x6);
  assign n121 = ~x0 & ~x5;
  assign n122 = (x1 | (x0 ? (x2 | (~x3 ^ x4)) : (~x2 | (x3 ^ x4)))) & (x0 | ~x1 | ~x3 | (x2 & x4));
  assign z06 = n124 | (n114 & ~n129) | (~x2 & ~n128);
  assign n124 = ~x0 & (x5 ? (n125 & n127) : ~n126);
  assign n125 = ~x1 & ~x3;
  assign n126 = (~x3 | ~x4 | (x1 ? (~x2 ^ ~x6) : (x2 | ~x6))) & (x1 | x3 | x4 | (~x2 ^ x6));
  assign n127 = ~x6 & (x2 ^ ~x4);
  assign n128 = (x1 | ((~x0 | x5 | (x3 & ~x4)) & (~x4 | ~x5 | (x0 & x3)))) & (x0 | ((~x3 | x4 | x5) & (~x1 | ((x4 | ~x5) & (x3 | ~x4 | x5)))));
  assign n129 = x1 ? ((~x3 | ~x4 | ~x5) & (x4 | x5)) : (~x4 | x5);
  assign z07 = (x2 | n131 | n133 | ~n134) & (~x2 | ~n137);
  assign n131 = ~x0 & ~n132;
  assign n132 = x1 ? (x6 | ((x4 | ~x5) & (x3 | (x4 & ~x5)))) : ((~x4 | (x3 ? (~x5 ^ x6) : (x5 | x6))) & (~x5 | ~x6 | x3 | x4));
  assign n133 = ~x1 & ((~x4 & x5 & ~x0 & x3) | (x4 & (x0 ^ (~x3 & x5))));
  assign n134 = x0 ? (x1 | x6 | (~n135 & ~n136)) : (~x1 | ~n136);
  assign n135 = ~x3 & x5;
  assign n136 = ~x5 & x3 & ~x4;
  assign n137 = (~x0 | x4 | ~n78 | ~n125) & (x0 | n138);
  assign n138 = x4 ? (x1 ? ((x5 & x6) | (~x3 & (x5 | x6))) : (x3 & ~x5)) : ((~x1 & (x5 | (~x3 & ~x6))) | (x3 & ~x5 & (x1 | x6)));
  assign z08 = ~n142 | (~x1 & (x2 ? ~n141 : ~n140));
  assign n140 = (~x6 | (x0 ? (x3 ? (x4 | x5) : (~x4 | ~x5)) : ((x4 | ~x5) & (x3 | ~x4 | x5)))) & (~x0 | x3 | x6 | (~x4 ^ x5));
  assign n141 = (x5 | ((x0 | (x3 ? (x4 | ~x6) : (~x4 | x6))) & (~x0 | x3 | x4 | ~x6))) & (x0 | ~x3 | ~x5 | (x4 ^ x6));
  assign n142 = ~n145 & (~n75 | n143) & (x0 | n144);
  assign n143 = (~x6 | ((~x2 | x3 | (~x4 ^ x5)) & (x2 | ~x3 | ~x4 | x5))) & (x2 | ~x3 | x6 | (x4 ^ x5));
  assign n144 = x2 ? ((~x1 | ((~x3 | ~x4 | ~x6) & (x4 | x6))) & (x1 | ~x4 | (~x3 ^ x6)) & (x3 | x4 | x6)) : (x1 ? ((x4 | ~x6) & (x3 | ~x4 | x6)) : (~x3 | (x4 ^ x6)));
  assign n145 = n76 & ~x6 & x3 & x4;
  assign z09 = n148 | ~n151 | (n75 & ~n147);
  assign n147 = x6 ? ((~x3 ^ ~x5) | (~x2 ^ ~x4)) : ((~x2 | x3 | ~x5) & (x2 | ~x3 | x4 | x5));
  assign n148 = ~x1 & (x4 ? ~n150 : ~n149);
  assign n149 = (x3 | ((~x0 | x6 | (~x2 ^ ~x5)) & (x0 | ~x2 | ~x5 | ~x6))) & (x2 | ((~x3 | (~x5 ^ x6)) & (x0 | x5 | ~x6)));
  assign n150 = (x2 | ((x5 | ~x6 | ~x0 | ~x3) & (~x5 | x6 | x0 | x3))) & (x0 | ~x2 | (x3 ? (~x5 ^ x6) : (x5 | x6)));
  assign n151 = (n152 | n153) & (x0 | n154);
  assign n152 = x3 ^ x5;
  assign n153 = (x1 | x2 | ~x4) & (x0 | ~x1 | ~x2 | x4);
  assign n154 = (~x1 | x2 | (x3 ? (~x4 | x5) : ~x5)) & (x1 | ~x2 | ~x3 | x4 | x5);
  assign z10 = n156 | n160 | ~n161 | (~x1 & ~n159);
  assign n156 = ~x3 & ((n75 & ~n158) | (~x1 & ~n157));
  assign n157 = x0 ? (x4 | (x2 ? (x5 | ~x6) : (~x5 | x6))) : ((~x4 | ((~x5 | x6) & (x2 | x5 | ~x6))) & (~x2 | ~x5 | x6));
  assign n158 = (~x2 | x4 | (~x5 ^ x6)) & (x2 | ~x4 | x5 | ~x6);
  assign n159 = (x0 | ((x4 | ~x6 | x2 | x3) & (~x3 | (x2 ? (~x4 ^ x6) : (~x4 | ~x6))))) & (x2 | ((~x3 | x4 | x6) & (~x4 | ~x6 | ~x0 | x3)));
  assign n160 = n75 & ((~x2 & x3 & ~x4 & ~x6) | (x2 & (x3 ? (~x4 & x6) : (x4 & ~x6))));
  assign n161 = x5 ? ((~x6 | n162) & (~x2 | x6 | ~n163)) : ((x6 | n162) & (x2 | ~x6 | ~n163));
  assign n162 = (x2 | (x3 ^ x4) | (~x0 ^ x1)) & (x0 | x1 | ~x2 | x3 | ~x4);
  assign n163 = x4 & x3 & ~x0 & x1;
  assign z11 = ~n165 | (~x4 & n125 & (~n166 | ~n167));
  assign n165 = (x0 & (x1 | x2)) | (~x0 & ~x1 & ~x2 & ~x3 & ~x4);
  assign n166 = x0 ? (~x2 | x5) : (x2 | ~x5);
  assign n167 = (x0 | x2 | x5 | ~x6) & (~x0 | ~x2 | ~x5 | x6);
  assign z16 = ~n172 | (~x1 & ~n169);
  assign n169 = (x3 | n170) & (x0 | ~x2 | ~x3 | ~n171);
  assign n170 = x0 ? ((x4 | ~x5 | x6) & (x5 | ~x6 | x2 | ~x4)) : (~x2 | (x4 ? (~x5 | x6) : (x5 ^ x6)));
  assign n171 = x6 & ~x4 & ~x5;
  assign n172 = (x1 | n174) & (~n75 | (n173 & n175));
  assign n173 = (x2 | ((x5 | ~x6 | ~x3 | x4) & (~x5 | x6 | x3 | ~x4))) & (~x3 | ~x4 | (x5 ^ x6));
  assign n174 = (x2 | ((~x0 | ~x4 | (~x3 ^ x5)) & (x4 | ((~x3 | ~x5) & (x0 | (~x3 & ~x5)))))) & (x0 | (x3 ? ~x5 : (~x4 | x5))) & (~x0 | x3 | x4 | x5);
  assign n175 = x3 ? (x4 | ~x5) : (x5 & (~x2 | ~x4));
  assign z17 = n180 | n186 | (x2 ? ~n177 : ~n185);
  assign n177 = x0 ? (~n178 | ~n125) : n179;
  assign n178 = ~x6 & ~x4 & x5;
  assign n179 = x1 ? (x3 ? (~x4 | x6) : (x4 | ~x6)) : ((~x3 | x4 | x5 | x6) & (x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))));
  assign n180 = ~x2 & (n182 | n184 | (~x1 & ~n181));
  assign n181 = (x5 | ((~x0 | (x3 ? (x4 | ~x6) : (~x4 | x6))) & (x0 | x3 | x4 | ~x6))) & (x0 | ~x3 | ~x4 | ~x5 | ~x6);
  assign n182 = ~n183 & (x3 ? (~x6 & n75) : (x6 & n108));
  assign n183 = x4 ^ x5;
  assign n184 = x6 & n75 & (x3 ? (~x4 & x5) : (x4 & ~x5));
  assign n185 = (x1 | (x0 ? (x3 ? ~x4 : (x4 | ~x5)) : ((~x4 | x5) & (~x3 | x4 | ~x5)))) & (x0 | (x3 ? (~x4 | x5) : (x4 ? ~x5 : ~x1)));
  assign n186 = n114 & (x3 ? (x1 ? (~x4 & ~x5) : (x4 ^ x5)) : ((x4 & x5) | (~x1 & ~x4 & ~x5)));
  assign z18 = ~n192 | (~x0 & (~n188 | ~n191));
  assign n188 = (~x4 | n189) & (x1 | x4 | n190);
  assign n189 = x1 ? ((~x2 | ~x3 | x5 | ~x6) & (x2 | x3 | ~x5 | x6)) : (x2 | ~x3 | (~x5 ^ x6));
  assign n190 = (~x2 | ~x3 | (x5 ^ x6)) & (x2 | x3 | ~x5 | ~x6);
  assign n191 = x1 ? ((x4 | ~x6 | x2 | x3) & (~x2 | (x3 ? (~x4 ^ x6) : (x4 | x6)))) : (~x6 | (x2 ? (~x3 | ~x4) : (~x3 ^ x4)));
  assign n192 = ~n194 & n195 & (x4 | ~n108 | n193);
  assign n193 = (~x2 | x3 | x5 | ~x6) & (x2 | ~x3 | (x5 ^ x6));
  assign n194 = ~x0 & ((x1 & (x2 ? (~x3 & x6) : (x3 & ~x6))) | (~x1 & x2 & ~x3 & ~x6));
  assign n195 = ~n196 & (~x6 | ~n76 | ~x3 | ~x4);
  assign n196 = ~x6 & ~x3 & ~x2 & x0 & ~x1;
  assign z19 = ~n204 | n198 | (~x1 & ~x5 & ~n203);
  assign n198 = ~x3 & (n200 | (~x4 & ~n199));
  assign n199 = (x0 | ((x5 | ~x6 | x1 | x2) & (~x1 | ~x2 | x6))) & (~x5 | x6 | ~x0 | x1);
  assign n200 = n202 & (x2 ? n201 : n78);
  assign n201 = x5 & x6;
  assign n202 = x4 & ~x0 & x1;
  assign n203 = (x0 | x2 | ~x3 | ~x4) & (x4 | (x0 ? (~x2 ^ x3) : (~x2 | ~x3)));
  assign n204 = ~n206 & ~n207 & (~x6 | ~n205 | n208);
  assign n205 = ~x0 & x3;
  assign n206 = ~x0 & (x1 ? (x2 ? (x3 & ~x4) : (~x3 ^ x4)) : (x2 ? (~x3 & x4) : (x3 & ~x4)));
  assign n207 = x4 & ~x3 & ~x2 & x0 & ~x1;
  assign n208 = (~x1 | (x2 ? (~x4 | x5) : (x4 | ~x5))) & (x1 | ~x2 | ~x4 | ~x5);
  assign z20 = ~n216 | (~x3 & ~n210) | (~x1 & ~n215);
  assign n210 = (~n212 | n214) & (x4 | n211 | n213);
  assign n211 = x2 ^ ~x6;
  assign n212 = ~x0 & x4;
  assign n213 = x0 ^ (~x1 & x5);
  assign n214 = (~x2 | ~x5 | x6) & (~x1 | x5 | (~x2 ^ ~x6));
  assign n215 = (x2 | ((~x0 | (x4 ^ x5)) & (~x4 | (~x3 ^ x5)) & (x0 | ((~x4 | x5) & (~x3 | x4 | ~x5))))) & (x0 | ~x2 | x4 | (~x3 ^ x5));
  assign n216 = ~x3 | ((~n217 | ~n218) & (x0 | n219));
  assign n217 = ~x4 & x5;
  assign n218 = x2 & ~x0 & x1;
  assign n219 = (~x4 | ((~x2 | ((x5 | ~x6) & (x1 | ~x5 | x6))) & (~x5 | ~x6 | ~x1 | x2))) & (~x1 | x2 | x4 | (~x5 ^ x6));
  assign z21 = n226 | ~n222 | (~x0 & ~x1 & n221);
  assign n221 = x2 & x3 & (x4 ^ x6);
  assign n222 = ~n225 & (~n93 | ~n224 | ~x0 | ~n223);
  assign n223 = ~x5 & x6;
  assign n224 = ~x1 & x2;
  assign n225 = ~x2 & ((~x1 & x6) | (~x0 & x1 & ~x6));
  assign n226 = ~x0 & x2 & (x1 ? (~x3 ^ x6) : (~x3 & x6));
  assign z22 = n232 | n233 | (~x1 & (~n228 | ~n231));
  assign n228 = (x0 | x2 | ~x3 | ~n229) & (~x0 | x3 | n230);
  assign n229 = x6 & x4 & ~x5;
  assign n230 = (x2 | ~x4 | x5 | ~x6) & (~x2 | x4 | ~x5 | x6);
  assign n231 = x2 ? ((x3 | x4 | x5) & (x0 | (x3 & x4))) : ((~x3 | ~x4 | ~x5) & (~x0 | (~x3 & (~x4 | ~x5))));
  assign n232 = n75 & (x2 ? ~x3 : (n92 | (x3 & n217)));
  assign n233 = n234 & n223 & n77;
  assign n234 = ~x2 & ~x0 & x1;
  assign z23 = n240 | ~n242 | (~x1 & (~n236 | ~n239));
  assign n236 = (x3 | n238) & (x0 | x2 | ~x3 | ~n237);
  assign n237 = ~x6 & x4 & ~x5;
  assign n238 = (~x0 | x6 | (x2 ? (x4 | ~x5) : (~x4 | x5))) & (x0 | ~x2 | ~x4 | x5 | ~x6);
  assign n239 = x0 ? (x2 | (x3 ^ x4)) : (~x3 | x4);
  assign n240 = ~n241 & ~x0 & x5;
  assign n241 = x1 ? (x2 ? (~x3 | ~x4) : (x3 | x4)) : (x3 | ~x4);
  assign n242 = ~n244 & ~n246 & (~x0 | ~n224 | ~n243);
  assign n243 = ~x5 & ~x3 & ~x4;
  assign n244 = n75 & n245 & (x2 ? (x4 & x6) : (~x4 & ~x6));
  assign n245 = x3 & ~x5;
  assign n246 = ~x0 & x1 & ~x3 & (x2 | x4);
  assign z24 = (~x1 & ~n249) | (~x0 & (x1 ? ~n252 : ~n248));
  assign n248 = (x5 | ((~x2 | x3 | x4 | ~x6) & (x2 | ~x4 | (x3 & x6)))) & (~x5 | ~x6 | x2 | x4);
  assign n249 = x0 ? (x2 ? (~n93 | n251) : n250) : (~x2 | n250);
  assign n250 = (~x3 | (x4 & (~x5 | ~x6))) & (x4 | ~x5) & (x3 | ~x4 | x5 | x6);
  assign n251 = x5 & x6;
  assign n252 = (x3 | (x2 ? ~x4 : (x4 | x5))) & (~x2 | (x4 ? (x5 | x6) : (~x5 | ~x6))) & (x2 | (x4 ? (~x5 & (~x3 | ~x6)) : (x5 | x6)));
  assign z25 = n256 | ~n260 | (~n254 & ~n255);
  assign n254 = x5 ^ ~x6;
  assign n255 = (~x0 | x1 | ~x2 | x3 | x4) & (x0 | ((~x1 | ~x2 | ~x3 | x4) & (x1 | (x2 ? (~x3 | ~x4) : x4))));
  assign n256 = ~x2 & ((~n152 & ~n258) | (n257 & n259));
  assign n257 = x6 & x4 & x5;
  assign n258 = (x0 | ~x1 | x4 | ~x6) & (~x0 | x1 | ~x4 | x6);
  assign n259 = ~x3 & ~x0 & x1;
  assign n260 = ~n261 & ~n262 & n264 & (~n76 | ~n263);
  assign n261 = x5 & n114 & (x1 ? (~x3 & x4) : ~x4);
  assign n262 = ~x2 & ~n152 & (x0 ? (~x1 & ~x4) : (x1 & x4));
  assign n263 = x6 & ~x3 & x5;
  assign n264 = (~n114 | n266) & (x6 | ~n121 | n265);
  assign n265 = (x2 | ~x3) & (x1 | ~x2 | x3);
  assign n266 = (~x4 | ~x5 | ~x6 | x1 | x3) & (~x1 | x4 | x6 | (x3 ^ ~x5));
  assign z26 = n275 | n273 | n268 | n270;
  assign n268 = ~x3 & ((n76 & n171) | (~x0 & ~n269));
  assign n269 = x1 ? (((~x2 ^ x6) | (~x4 ^ x5)) & (x2 | x4 | x5 | x6)) : (x2 ? (~x6 | (x4 ^ x5)) : (x6 | (~x4 ^ x5)));
  assign n270 = x3 & (n271 | (n212 & ~n272));
  assign n271 = ~n254 & ((x0 & ~x1 & ~x2 & x4) | (~x0 & ~x4 & (~x1 ^ x2)));
  assign n272 = (~x5 | ~x6 | ~x1 | ~x2) & (x1 | x2 | (x5 ^ x6));
  assign n273 = ~x1 & ~n274;
  assign n274 = x4 ? ((x0 | (x2 ? x6 : (x3 | ~x6))) & (~x0 | x2 | x3 | x6)) : ((~x0 | (x2 ? (x3 | x6) : (~x3 | ~x6))) & (x0 | ~x2 | ~x3 | ~x6));
  assign n275 = n75 & ((~x2 & x3 & ~x4 & ~x6) | (x4 & (x2 ? (~x3 ^ ~x6) : (x3 & x6))));
  assign z27 = n277 | n279 | ~n283 | (~x1 & ~n282);
  assign n277 = x3 & ((~x6 & ~n278) | (n257 & n218));
  assign n278 = (x0 | ((x4 | ~x5 | x1 | ~x2) & (~x1 | x5 | (x2 & ~x4)))) & (~x0 | x1 | x2 | x4 | ~x5);
  assign n279 = ~x3 & (n281 | (~x1 & ~n280));
  assign n280 = (x2 | ((x5 | ~x6 | x0 | ~x4) & (~x0 | ~x5 | (~x4 ^ x6)))) & (x0 | ~x2 | ((~x5 | ~x6) & (x4 | x5 | x6)));
  assign n281 = x6 & n75 & (x2 ? ~x5 : (x4 & x5));
  assign n282 = (~x3 | ((x2 | ~x4 | ~x5) & (x0 | (x2 ? ~x4 : ~x5)))) & (~x0 | x2 | x3 | x4 | x5);
  assign n283 = x3 ? (x4 | n284) : ((~n217 | ~n234) & (~x4 | n284));
  assign n284 = (~x0 | x1 | x2 | x5) & (x0 | ~x2 | (~x1 ^ ~x5));
  assign z28 = ~n293 | (~x1 & (n286 | n287 | n290));
  assign n286 = n118 & ((~x4 & x5 & ~x6) | (~x3 & ~x5 & x6));
  assign n287 = ~n288 & ~n289;
  assign n288 = x0 ? (x2 | ~x3) : (~x2 | x3);
  assign n289 = x4 ? (x5 | x6) : (~x5 | ~x6);
  assign n290 = ~n291 & ((n94 & n292) | (n77 & n114));
  assign n291 = x5 ^ x6;
  assign n292 = ~x3 & x4;
  assign n293 = (x1 | n296) & (~n75 | (n294 & n295));
  assign n294 = x2 ? (x4 | ~x5) : (~x4 | x5);
  assign n295 = ((~x3 ^ ~x6) | (x2 ? (~x4 | ~x5) : (x4 | x5))) & (x5 | ~x6 | ~x2 | x3) & (x2 | ~x3 | ~x4 | ~x5 | x6);
  assign n296 = x5 ? ((~x0 | x2 | x3 | x4) & (x0 | ~x4 | (x2 & x3))) : ((x0 | ~x2 | ~x3 | ~x4) & (~x0 | x4 | (~x2 ^ x3)));
  assign z29 = ~n301 | (~x1 & (~n298 | ~n300));
  assign n298 = (~x5 | n299) & (x4 | x5 | x6 | n288);
  assign n299 = (x2 | x4 | ~x6 | (~x0 & ~x3)) & (x0 | ~x2 | x3 | ~x4);
  assign n300 = (x3 | (x0 ? ((x4 | x6) & (x2 | ~x4 | ~x6)) : (x4 | ~x6))) & (x0 | ((~x2 | x4 | ~x6) & (~x3 | x6 | (x2 & ~x4))));
  assign n301 = ~n303 & ~n304 & (n254 | n302);
  assign n302 = (x0 | ((x3 | ~x4 | x1 | x2) & (~x1 | x4 | (x2 & x3)))) & (~x0 | x1 | x2 | ~x3 | ~x4);
  assign n303 = n75 & (x2 ? (x3 ? (~x4 & ~x6) : (x4 & x6)) : (x4 & (x3 ^ ~x6)));
  assign n304 = n202 & ((~x2 & ~x3 & x5 & x6) | (~x5 & ((x3 & ~x6) | (x2 & (x3 | ~x6)))));
  assign z30 = ~n308 | (~x0 & (x6 ? ~n307 : ~n306));
  assign n306 = (x1 | ~x2 | ~x3 | x4 | ~x5) & (~x1 | x2 | x3 | ~x4 | x5);
  assign n307 = (x1 | x2 | x4 | (x3 ^ x5)) & (~x2 | ~x4 | ((x3 | x5) & (~x1 | ~x3 | ~x5)));
  assign n308 = ~n310 & (~n76 | ~n311) & (x2 | n309);
  assign n309 = (~x4 & ((x3 & ~x5) | (~x0 & ~x1 & (x3 | ~x5)))) | (x1 & (x0 | (~x3 & x4))) | (x4 & ((~x3 & x5) | (x0 & (~x3 | x5))));
  assign n310 = ~x0 & x2 & (x3 ? (~x4 & ~x5) : (x4 & x5));
  assign n311 = ~x6 & x5 & x3 & x4;
  assign z31 = n313 | n317 | n320 | (~x1 & ~n316);
  assign n313 = ~x5 & (x0 ? (n224 & n314) : ~n315);
  assign n314 = ~x6 & ~x3 & ~x4;
  assign n315 = (~x4 | ((~x2 | x3 | ~x6) & (~x1 | ((x3 | ~x6) & (x2 | ~x3 | x6))))) & (x1 | x2 | x4 | (~x3 ^ x6));
  assign n316 = x0 ? (x2 | (x3 ? (x4 | ~x5) : x5)) : (x3 ? (~x4 | x5) : ((~x4 | ~x5) & (~x2 | x4 | x5)));
  assign n317 = n75 & ((~x4 & ~n152) | (n318 & n319));
  assign n318 = ~x2 & ~x3;
  assign n319 = x4 & x5;
  assign n320 = x5 & ((~n321 & ~n322) | (n314 & n234));
  assign n321 = x3 ^ x6;
  assign n322 = (~x0 | x1 | x2 | ~x4) & (x0 | (x1 ? (~x2 | ~x4) : x4));
  assign z32 = ~n327 | (~x5 & ~n325) | (~x0 & ~n324);
  assign n324 = x1 ? ((~x4 | x5 | ~x6) & (~x5 | x6 | ~x2 | x4)) : ((~x4 | ~x5 | x6) & (x2 | (~x4 ^ x6)));
  assign n325 = ~n326 & (~x3 | x4 | x6 | ~n75);
  assign n326 = x6 & n125 & ((x0 & ~x2 & x4) | (x2 & (~x0 | ~x4)));
  assign n327 = n329 & (n291 | n328);
  assign n328 = (~x0 | x1 | x2 | ~x4) & (x0 | (x1 ? ((~x2 | ~x3 | ~x4) & (x3 | x4)) : (~x2 | x4)));
  assign n329 = (~n76 | ~n178) & (~x5 | ~n75 | n330);
  assign n330 = (~x2 | x3 | ~x4 | ~x6) & (x2 | ~x3 | x4 | x6);
  assign z33 = ~n332 | (~x1 & ~n340) | (~x0 & ~n341);
  assign n332 = ~n334 & ~n336 & n338 & (n211 | n333);
  assign n333 = (~x0 | x1 | x3 | x4 | ~x5) & (x0 | ((x1 | x3 | x4 | x5) & (~x1 | ~x3 | (~x4 ^ x5))));
  assign n334 = ~x6 & ((n76 & n136) | (~x0 & ~n335));
  assign n335 = (x1 | ~x2 | ~x3 | ~x4 | x5) & (~x1 | x3 | ~x5 | (x2 ^ ~x4));
  assign n336 = n337 & x2 & n75;
  assign n337 = x5 & x6 & (x3 ^ x4);
  assign n338 = x3 ? (~n75 | n339) : (~n76 | ~n78);
  assign n339 = x2 ? (~x4 | ~x5) : (x4 | x5);
  assign n340 = (x0 | x2 | x3 | ~x5) & (x5 | (x0 ? (x2 ? (x3 | x4) : (~x3 | ~x4)) : (~x2 | (~x3 ^ x4))));
  assign n341 = (x2 | ((~x1 | (x3 ? (~x5 | x6) : (x5 | ~x6))) & (~x5 | ~x6 | x1 | ~x3))) & (x1 | ~x2 | x3 | ~x5 | ~x6);
  assign z34 = n343 | n347 | ~n348 | (~x3 & ~n346);
  assign n343 = ~x1 & ((n212 & ~n345) | (~x4 & ~n344));
  assign n344 = (~x0 | x2 | ~x3 | x5 | x6) & (~x2 | ((x3 | ~x5 | x6) & (x5 | ~x6 | x0 | ~x3)));
  assign n345 = (x2 | ~x3 | x5 | ~x6) & (~x2 | (x3 ? (~x5 | ~x6) : (x5 | x6)));
  assign n346 = (x2 | (x5 ^ x6) | (~x0 ^ x1)) & (x0 | ~x2 | ((x5 | ~x6) & (~x1 | ~x5 | x6)));
  assign n347 = ~x6 & n205 & ((~x2 & x5) | (~x1 & x2 & ~x5));
  assign n348 = n350 & (~n349 | (x3 ? (x4 | ~x6) : (~x4 | x6)));
  assign n349 = x5 & ~x2 & ~x0 & x1;
  assign n350 = (x0 | ((x3 | ~x5 | x1 | x2) & (~x1 | ~x2 | ~x3 | x5))) & (~x0 | x1 | x2 | ~x3 | ~x5);
  assign z35 = ~n355 | (~x2 & (n352 | n353));
  assign n352 = ~n321 & (x4 ? (~x5 & n75) : (x5 & n108));
  assign n353 = n354 & (x0 ? (~x5 & ~x6) : (x5 ^ x6));
  assign n354 = ~x4 & ~x1 & x3;
  assign n355 = ~n357 & ((x0 & (x5 | ~n358)) | (n356 & (~n358 | (~x0 & ~x5))));
  assign n356 = (x3 | ~x6 | ((x2 | ~x4) & (x1 | (x2 & ~x4)))) & (~x4 | x6 | x1 | ~x3);
  assign n357 = ~n321 & ((x0 & ~x1 & ~x2 & x4) | (~x0 & ((x2 & ~x4) | (x1 & (x2 | ~x4)))));
  assign n358 = x6 & ~x4 & ~x3 & ~x1 & x2;
  assign z36 = n360 | n364 | n366 | (~x1 & ~n363);
  assign n360 = ~x2 & ((n75 & ~n362) | (~x1 & ~n361));
  assign n361 = (x0 | x3 | ~x4 | x5 | ~x6) & (~x0 | ((x3 | x4 | x5 | x6) & (~x5 | ~x6 | ~x3 | ~x4)));
  assign n362 = (~x3 | ~x4 | ~x5 | x6) & (x3 | x5 | (x4 ^ ~x6));
  assign n363 = (x0 | (x2 ? (~x3 | x4) : (~x4 | ~x5))) & (~x2 | x3 | x4 | x5) & (x2 | (x3 ? (x4 | x5) : (~x4 | ~x5)));
  assign n364 = n75 & ((~x2 & ~x4 & x5) | (x4 & (x2 | (~x5 & n365))));
  assign n365 = ~x2 & x3;
  assign n366 = n217 & n367 & ((~x1 & ~x6) | (~x0 & x1 & x6));
  assign n367 = x2 & ~x3;
  assign z37 = n369 | n372 | ~n374 | (~n254 & ~n373);
  assign n369 = ~x0 & (n371 | (x4 & ~n370));
  assign n370 = x2 ? (~x5 | ~x6 | (x1 & ~x3)) : (x5 | x6 | (~x1 & x3));
  assign n371 = ~x4 & n318 & ((x5 & x6) | (x1 & ~x5 & ~x6));
  assign n372 = n205 & ((~x2 & ~x4 & ~x5) | (~x1 & (x2 ? (~x4 & x5) : ~x5)));
  assign n373 = x2 ? (x3 | ((x1 | x4) & (x0 | (x1 & x4)))) : (~x3 | ~x4 | (~x0 ^ x1));
  assign n374 = x3 ? (x4 | n375) : (x4 ? n375 : (~n76 | ~n78));
  assign n375 = (~x0 | x1 | x2 | x5) & (x0 | ~x1 | ~x2 | ~x5);
  assign z38 = ~n379 | (~x2 & (n378 | (~x1 & ~n377)));
  assign n377 = (~x6 | (~x0 ^ x4) | (x3 ^ ~x5)) & (x0 | x3 | x6 | (~x4 ^ x5));
  assign n378 = n202 & (x3 ? (x5 & ~x6) : (~x5 ^ x6));
  assign n379 = ~n382 & (x1 ? (x0 | n381) : n380);
  assign n380 = x0 ? ((x3 | x4 | x6) & (x2 | ~x4 | (~x3 ^ x6))) : ((~x2 | x3 | x6) & (~x3 | x4 | ~x6));
  assign n381 = x3 ? (x4 | ~x6) : ((x4 | x6) & (~x2 | ~x4 | ~x6));
  assign n382 = n319 & n114 & ((x3 & ~x6) | (~x1 & ~x3 & x6));
  assign z39 = ~n386 | (~x2 & (n385 | (~x3 & ~n384)));
  assign n384 = (x0 | ~x1 | x4 | x5) & (x1 | ~x4 | ~x5 | (~x0 & x6));
  assign n385 = n205 & (x1 ? (x4 & n223) : (~x4 & ~n291));
  assign n386 = (x2 | n388) & (~n114 | (n387 & n389));
  assign n387 = (x1 | x4 | x5 | x6) & (~x4 | (x1 ? (~x5 ^ x6) : (~x5 | ~x6)));
  assign n388 = (x1 | (x0 ? (x4 ? x5 : (~x5 | ~x6)) : (x4 | (~x5 ^ x6)))) & (x0 | ~x4 | ~x5 | (~x1 & ~x6));
  assign n389 = x1 ? (x3 | ((~x4 | ~x5 | ~x6) & (x5 | x6))) : (~x3 | ((x5 | ~x6) & (~x4 | ~x5 | x6)));
  assign z40 = ~n395 | (~x0 & (~n391 | ~n394));
  assign n391 = (x1 | x2 | x3 | ~n392) & (~x3 | (x1 ? (~x2 | n393) : (x2 ? ~n392 : n393)));
  assign n392 = x6 & ~x4 & x5;
  assign n393 = x4 ? (~x5 | ~x6) : (x5 | x6);
  assign n394 = x1 ? (x6 | (x2 ? (x3 | ~x4) : (~x3 | x4))) : (x2 ? (x3 ? (~x4 | ~x6) : x4) : (x3 | ~x4));
  assign n395 = ~n396 & ~n398 & ~n399 & (x6 | n397);
  assign n396 = n77 & n201 & n76;
  assign n397 = (~x0 | x1 | x2 | x3 | x5) & (x0 | ~x5 | (x1 ? (x2 | x3) : (~x2 | ~x3)));
  assign n398 = ~x2 & n108 & (x3 ? x4 : (~x4 & x6));
  assign n399 = n223 & n75 & (x2 ^ x3);
  assign z41 = n401 | ~n406 | (~n291 & ~n405);
  assign n401 = ~x0 & (n402 | (~x4 & x6 & ~n404));
  assign n402 = ~n403 & (n135 | n245);
  assign n403 = (x1 | ~x2 | (x4 ^ x6)) & (~x1 | x2 | ~x4 | x6);
  assign n404 = (x1 | ~x2 | x3 | x5) & (~x3 | (x1 ? (x2 ^ ~x5) : (x2 | x5)));
  assign n405 = (~x0 | x1 | x2 | ~x3 | x4) & (x0 | ((~x3 | ~x4 | x1 | x2) & (~x1 | x3 | (x2 ^ x4))));
  assign n406 = ~n409 & n411 & (x0 | (n407 & n408));
  assign n407 = (~x3 | ((~x1 | x2 | (x4 ^ x5)) & (x1 | ~x2 | x4 | ~x5))) & (x1 | ~x2 | x3 | ~x4 | x5);
  assign n408 = (x1 | x2 | x3 | (~x4 ^ x6)) & (~x3 | ~x4 | ~x6 | ~x1 | ~x2);
  assign n409 = ~n410 & (x3 ? n113 : n223);
  assign n410 = (~x0 | x1 | x2 | ~x4) & (x0 | ~x1 | ~x2 | x4);
  assign n411 = ~x0 | x1 | (x2 ? ~n243 : ~n314);
  assign z42 = ~n415 | (~x1 & (n414 | (~x0 & ~n413)));
  assign n413 = (x6 | ((~x3 | x4 | ~x5) & (~x2 | (x3 ? ~x5 : (x4 | x5))))) & (x2 | x3 | ~x4 | ~x5) & (~x6 | (x2 & ~x4) | (x3 ^ ~x5));
  assign n414 = n94 & (x3 ? (x4 ? (~x5 ^ x6) : (~x5 & x6)) : ((x5 & ~x6) | (x4 & ~x5 & x6)));
  assign n415 = ~n418 & (~n75 | n416) & (x3 | n417);
  assign n416 = x3 ? (x2 ? (x4 ? (~x5 | ~x6) : (x5 | x6)) : (~x5 | (~x4 ^ x6))) : ((x4 | ((x5 | ~x6) & (~x2 | ~x5 | x6))) & (x5 | x6 | (x2 & ~x4)));
  assign n417 = (x0 | ~x1 | ~x2 | ~x4 | ~x6) & (x1 | ((~x4 | x6 | x0 | ~x2) & (x4 | (x0 ? (~x2 ^ x6) : (~x2 | ~x6)))));
  assign n418 = n75 & n77 & (x2 ^ ~x6);
  assign z43 = ~n422 | (~x2 & (n421 | (~x1 & ~n420)));
  assign n420 = x6 ? ((x0 | ~x4 | (x3 & ~x5)) & (x4 | ~x5 | ~x0 | ~x3)) : (x0 ? (~x4 | (~x3 & x5)) : (~x3 | x5));
  assign n421 = n75 & ((x3 & ~x5 & (x4 ^ ~x6)) | (~x4 & x6 & (~x3 | x5)));
  assign n422 = ~n425 & (~n114 | n423) & (x0 | n424);
  assign n423 = (~x1 | x3 | (x4 ? (x5 | ~x6) : x6)) & (~x3 | ((x4 | (~x5 ^ x6)) & (x1 | ~x5 | x6)));
  assign n424 = (~x5 | (x1 ? (~x4 | (x2 ^ x3)) : (x2 | x4))) & (x1 | ~x2 | x3 | x5);
  assign n425 = n108 & ((x2 & ~x3 & ~x4 & ~x5) | (~x2 & (x3 ? (~x4 & ~x5) : x5)));
  assign z44 = ~n430 | (~x1 & (~n428 | (~x2 & ~n427)));
  assign n427 = x0 ? (~x6 | ((x3 | x4 | ~x5) & (~x4 | x5))) : (x6 | (~x4 ^ x5));
  assign n428 = (n291 | n429) & (x0 | ~n367 | ~n178);
  assign n429 = (x0 | ~x2 | x3 | ~x4) & (~x0 | x2 | ~x3 | x4);
  assign n430 = n433 & (n183 | n431) & (x1 | n432);
  assign n431 = (~x0 | x1 | x2 | x3 | x6) & (x0 | ((~x1 | (x2 ? (~x3 | x6) : (x3 | ~x6))) & (~x3 | ~x6 | x1 | ~x2)));
  assign n432 = (x0 | ~x4 | (x2 ? (~x3 | x6) : ~x6)) & (~x0 | ~x2 | x3 | x4 | x6);
  assign n433 = (~n75 | n434) & (~n113 | ~n292 | ~n218);
  assign n434 = (x2 | ~x4 | x6) & (x4 | ~x6 | (~x2 & ~x3));
  assign z45 = n441 | ~n444 | (~x0 & (~n436 | ~n443));
  assign n436 = ~n440 & n437 & ~n439;
  assign n437 = ~n438 & (x1 | ~x4 | ~n113 | ~n318);
  assign n438 = (x2 ? (x3 & x5) : (~x3 & ~x5)) & (x1 ^ x6);
  assign n439 = x1 & x6 & (x2 ? (x3 & ~x5) : (~x3 & x5));
  assign n440 = ~n254 & (x1 ? (x2 & n292) : (~x2 & n77));
  assign n441 = ~n442 & (x2 ? n93 : n92);
  assign n442 = (x1 | (x0 ? (x5 | x6) : ~x5)) & (x0 | x5 | (~x1 & ~x6));
  assign n443 = (~x1 | x2 | ~x3 | x4 | x5) & (x1 | ~x2 | x3 | ~x4 | ~x5);
  assign n444 = (x3 & x4) ? (~n201 | ~n76) : ~n445;
  assign n445 = x5 & ~x2 & x0 & ~x1;
  assign z46 = ~n450 | (~x1 & ~n447) | (~x0 & ~n449);
  assign n447 = (x4 | n448) & (~x4 | x5 | ~n205 | n211);
  assign n448 = (~x5 | ((x0 | (x2 ? (~x3 | ~x6) : x3)) & (~x0 | x2 | ~x3 | ~x6))) & (~x2 | x5 | ((x3 | ~x6) & (x0 | ~x3 | x6)));
  assign n449 = (~x1 | x2 | ~x3 | ~x4 | x6) & (x1 | ~x6 | (x2 ? (~x3 | ~x4) : (~x3 ^ x4)));
  assign n450 = ~n196 & ~n452 & ~n453 & (~n75 | n451);
  assign n451 = (~x2 | x3 | x4 | x5 | ~x6) & (x2 | ~x5 | x6 | (~x3 ^ x4));
  assign n452 = ~x0 & ((x1 & x6 & (~x2 ^ x3)) | (~x1 & x2 & ~x3 & ~x6));
  assign n453 = ~n454 & ((n75 & n367) | (n365 & n108));
  assign n454 = x4 ^ x6;
  assign z47 = ~n462 | (~x0 & (n456 | ~n458));
  assign n456 = ~n457 & x1 & ~x4;
  assign n457 = (x2 | ~x3 | x5 | x6) & (x3 | (x2 ? (x5 ^ x6) : (x5 | ~x6)));
  assign n458 = n459 & (n289 | (x2 & ~x3) | (~x1 & (x2 | ~x3)));
  assign n459 = (~n237 | ~n460) & (n461 | (~x3 & ~x6));
  assign n460 = x3 & ~x1 & x2;
  assign n461 = (~x1 | x2 | ~x4 | ~x5) & (x1 | ~x2 | x4 | x5);
  assign n462 = n464 & (n254 | n463);
  assign n463 = (x0 | ~x1 | ~x2 | ~x3 | ~x4) & (x1 | ((x3 | (x0 ? (~x2 ^ x4) : (~x2 | ~x4))) & (x2 | ((~x3 | x4) & (x0 | (~x3 & x4))))));
  assign n464 = (n454 | n465) & (~n76 | ~n77 | ~n78);
  assign n465 = (~x0 | x1 | x2 | x3 | ~x5) & (x0 | ~x1 | (x2 ? ~x5 : (x3 | x5)));
  assign z48 = ~n469 | (~x2 & (n468 | (~x0 & ~n467)));
  assign n467 = ((~x4 ^ x6) | (x1 ? (x3 | x5) : (~x3 | ~x5))) & (x3 | x4 | ~x5 | x6) & (x5 | ((~x3 | ~x4 | ~x6) & (x1 | ((~x4 | ~x6) & (~x3 | x4 | x6)))));
  assign n468 = n108 & ((~x3 & x6 & (~x4 ^ x5)) | (~x6 & ((x4 & ~x5) | (x3 & ~x4 & x5))));
  assign n469 = ~n472 & (~n114 | n470) & (x1 | n471);
  assign n470 = ((~x4 ^ x6) | (x1 ? (x3 | ~x5) : (~x3 | x5))) & (~x4 | ~x5 | ~x6 | (x1 & ~x3)) & (x4 | x5 | x6 | (~x1 & x3));
  assign n471 = x0 ? ((~x2 | x3 | x4 | x6) & (~x4 | ~x6 | x2 | ~x3)) : (~x2 | x3 | (~x4 ^ x6));
  assign n472 = n75 & ((~x2 & ~x3 & x4 & x6) | (x3 & (x2 ? (x4 ^ x6) : (~x4 & ~x6))));
  assign z49 = n474 | ~n478 | (~n291 & ~n477);
  assign n474 = ~x0 & (x1 ? ~n476 : ~n475);
  assign n475 = (~x4 | ~x5 | ~x6 | ~x2 | x3) & (x2 | ((x5 | ~x6 | x3 | x4) & (~x3 | x6 | (x4 ^ x5))));
  assign n476 = (x2 | x3 | x4 | ~x5 | x6) & (~x2 | ((~x3 | ~x6 | (x4 ^ x5)) & (x3 | x4 | x5 | x6)));
  assign n477 = (~x0 | x1 | x2 | x3 | x4) & (x0 | ((x1 | (x2 ? (~x3 | x4) : (x3 | ~x4))) & (~x3 | ~x4 | ~x1 | x2)));
  assign n478 = n481 & (n254 | n480) & (x1 | n479);
  assign n479 = (x3 | ((~x0 | (x2 ? (x4 | x5) : (~x4 | ~x5))) & (x0 | ~x2 | ~x4 | x5))) & (x0 | ~x3 | ~x5 | (~x2 ^ ~x4));
  assign n480 = (~x0 | x1 | x2 | ~x3 | x4) & (x0 | x3 | (x1 ? ~x4 : (~x2 | x4)));
  assign n481 = (~n75 | n482) & (~n92 | ~n223 | ~n76);
  assign n482 = (x2 | ~x3 | x4 | x5) & (~x2 | (x3 ? (~x4 | x5) : (x4 | ~x5)));
  assign z50 = n268 | n273 | n485 | (x3 & ~n484);
  assign n484 = ~n271 & (n291 | ~n212 | (~x1 ^ ~x2));
  assign n485 = n75 & ((~x2 & x3 & (~x4 ^ x6)) | (x2 & ~x3 & x4 & x6));
  assign z51 = ~n489 | (~x1 & (n488 | (~x0 & ~n487)));
  assign n487 = (x2 | x3 | ~x4 | x5 | ~x6) & (~x2 | (x3 ? (~x5 | x6) : ((~x5 | ~x6) & (x4 | x5 | x6))));
  assign n488 = x5 & n94 & (x3 ? (~x4 & ~x6) : (~x4 ^ ~x6));
  assign n489 = ~n492 & (~n75 | n490) & (x1 | n491);
  assign n490 = (x2 | ((~x3 | x5 | x6) & (~x5 | ~x6 | x3 | ~x4))) & (x5 | ((~x3 | ~x4 | x6) & (~x2 | x3 | ~x6)));
  assign n491 = (x2 | ((~x0 | x5 | (x3 & x4)) & (~x3 | ~x5 | (x0 & ~x4)))) & (x0 | ~x2 | x5 | (~x3 & ~x4));
  assign n492 = x5 & n75 & (~x2 ^ (x3 | x4));
  assign z52 = ~n497 | (~x1 & (~n495 | (~x0 & ~n494)));
  assign n494 = x2 ? ((~x5 | ~x6 | ~x3 | ~x4) & (x3 | (x4 ? (x5 | x6) : (~x5 | ~x6)))) : ((x4 | ~x5 | x6) & (x3 | x5 | ~x6));
  assign n495 = (n291 | n496) & (~x0 | ~n365 | ~n237);
  assign n496 = (~x0 | x2 | (~x3 ^ x4)) & (x0 | ~x2 | ~x3 | x4);
  assign n497 = (x1 | n499) & (~n75 | (n498 & n500));
  assign n498 = (x3 | ((~x2 | (~x5 ^ x6)) & (x5 | x6 | x2 | x4))) & (x2 | ~x3 | (x4 ? (~x5 | x6) : (x5 | ~x6)));
  assign n499 = (x0 | ~x4 | (x2 ? (~x3 | x5) : ~x5)) & (x3 | (x0 ? (x4 | (~x2 ^ x5)) : (~x4 | ~x5)));
  assign n500 = x2 ? (~x3 | ~x5) : (~x4 | x5);
  assign z53 = ~n505 | (~x2 & (~n503 | (x5 & ~n502)));
  assign n502 = (~x0 | x1 | x3 | x4 | ~x6) & (x0 | ((x4 | ~x6 | x1 | ~x3) & (~x1 | (x3 ? (x4 | x6) : (~x4 | ~x6)))));
  assign n503 = (n254 | n504) & (x0 | ~n237 | ~n116);
  assign n504 = (~x0 | x1 | ~x3 | ~x4) & (x0 | x3 | (x1 ^ ~x4));
  assign n505 = ~n508 & (~n114 | n506) & (x1 | n507);
  assign n506 = (~x1 | x3 | x4 | ~x5 | x6) & (x1 | ((~x4 | ~x5 | ~x6) & (x3 | (x4 ? ~x5 : (x5 | x6)))));
  assign n507 = (~x4 | ((x0 | ~x3 | x6) & (~x0 | x2 | x3 | ~x6))) & (x4 | (x0 ? ((x2 | ~x3 | ~x6) & (x3 | x6)) : (~x6 | (~x2 & x3)))) & (x0 | x2 | ~x3 | x6);
  assign n508 = n75 & (x2 ? (~x3 ^ ~x6) : (x4 & (x3 ^ ~x6)));
  assign z54 = ~n513 | n510 | (~x0 & x6 & ~n512);
  assign n510 = ~x1 & ~n511;
  assign n511 = (x0 | ~x2 | (x3 ? (x4 | x5) : (~x4 | ~x5))) & (x2 | ((x5 | (x0 ? (x3 ^ x4) : (x3 | ~x4))) & (x4 | ~x5 | x0 | x3)));
  assign n512 = x2 ? (x1 ? (x3 ? (~x4 | x5) : (x4 | ~x5)) : (~x4 | (x3 ^ x5))) : (x4 | (x1 ? (~x3 | x5) : (x3 ^ x5)));
  assign n513 = n405 & ~n514 & (~n93 | ~n113 | ~n76);
  assign n514 = x3 & n75 & (x2 ? (x4 & x5) : (x4 ^ x5));
  assign z55 = n516 | ~n520 | (n75 & ~n519);
  assign n516 = ~x1 & (x3 ? (x5 & ~n518) : ~n517);
  assign n517 = (x4 | ((x2 | (x0 ? (x5 ^ x6) : (x5 | ~x6))) & (x0 | ~x2 | x5 | x6))) & (x0 | ~x4 | ((~x5 | x6) & (~x2 | x5 | ~x6)));
  assign n518 = (~x0 | x2 | x4 | x6) & (x0 | ~x6 | (x2 ^ x4));
  assign n519 = (~x6 | ((x2 | ~x3 | x4 | x5) & (~x2 | (x3 ? (~x4 | x5) : (x4 | ~x5))))) & (~x4 | x6 | ((x3 | ~x5) & (x2 | ~x3 | x5)));
  assign n520 = (~x0 | x1 | x2 | n521) & (x0 | (n522 & (~x1 | ~x2 | n521)));
  assign n521 = x3 ? (x4 ^ x5) : (~x4 | x5);
  assign n522 = (~x2 | ~x3 | x4 | ~x5) & (~x1 | ((x3 | x4 | x5) & (x2 | (x3 ^ x5))));
  assign z56 = n524 | n527 | ~n529 | (~n152 & ~n526);
  assign n524 = ~x0 & (x1 ? (n365 & n171) : ~n525);
  assign n525 = (x6 | ((x2 | ~x3 | x4 | x5) & (~x2 | (x3 ? (~x4 | x5) : (x4 | ~x5))))) & (x2 | ~x5 | ~x6 | (~x3 ^ x4));
  assign n526 = (~x0 | x1 | x2 | x4 | ~x6) & (x0 | ((~x1 | x6 | (x2 ^ x4)) & (~x4 | ~x6 | x1 | ~x2)));
  assign n527 = ~x0 & ~n528;
  assign n528 = (x1 | ((x2 | (x3 ? (~x4 | x5) : (x4 | ~x5))) & (~x4 | ~x5 | ~x2 | x3))) & ((x3 ^ x5) | (x1 ? (x2 | ~x4) : (~x2 | x4)));
  assign n529 = n530 & n531 & (~x3 | ~n76 | ~n78);
  assign n530 = ~x0 | x1 | (x2 ? ~n243 : ~n135);
  assign n531 = x0 | ~x1 | ~x2 | (~n245 & ~n263);
  assign z57 = n536 | (x2 ? ~n538 : (~n533 | ~n537));
  assign n533 = ~n535 & (x0 ? (~n125 | ~n171) : n534);
  assign n534 = (~x1 | ~x3 | ~x4 | ~x5 | x6) & (x3 | ((~x4 | ~x5 | ~x6) & (x1 | x6 | (~x4 ^ x5))));
  assign n535 = ~n254 & ((n93 & n75) | (n92 & n108));
  assign n536 = n114 & (n115 | (n237 & n116));
  assign n537 = (~x4 | x6 | (x0 ? (x1 | x3) : (~x1 ^ x3))) & (~x3 | x4 | ~x6 | (x0 & x1));
  assign n538 = (x4 | ((~x0 | x1 | x3 | x6) & (x0 | ((~x3 | x6) & (x1 | x3 | ~x6))))) & (x0 | ~x4 | ~x6 | (~x1 & ~x3));
  assign z12 = z11;
  assign z13 = z11;
  assign z14 = z11;
  assign z15 = z11;
  assign z59 = z58;
  assign z60 = z58;
  assign z61 = z58;
  assign z62 = z58;
  assign z63 = z58;
  assign z64 = z58;
endmodule


