// Benchmark "256_256_mod" written by ABC on Thu Dec 01 02:21:14 2022

module const_256_256_mod ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z000, z001, z002, z003, z004, z005, z006, z007, z008, z009, z010, z011,
    z012, z013, z014, z015, z016, z017, z018, z019, z020, z021, z022, z023,
    z024, z025, z026, z027, z028, z029, z030, z031, z032, z033, z034, z035,
    z036, z037, z038, z039, z040, z041, z042, z043, z044, z045, z046, z047,
    z048, z049, z050, z051, z052, z053, z054, z055, z056, z057, z058, z059,
    z060, z061, z062, z063, z064, z065, z066, z067, z068, z069, z070, z071,
    z072, z073, z074, z075, z076, z077, z078, z079, z080, z081, z082, z083,
    z084, z085, z086, z087, z088, z089, z090, z091, z092, z093, z094, z095,
    z096, z097, z098, z099, z100, z101, z102, z103, z104, z105, z106, z107,
    z108, z109, z110, z111, z112, z113, z114, z115, z116, z117, z118, z119,
    z120, z121, z122, z123, z124, z125, z126, z127, z128, z129, z130, z131,
    z132, z133, z134, z135, z136, z137, z138, z139, z140, z141, z142, z143,
    z144, z145, z146, z147, z148, z149, z150, z151, z152, z153, z154, z155,
    z156, z157, z158, z159, z160, z161, z162, z163, z164, z165, z166, z167,
    z168, z169, z170, z171, z172, z173, z174, z175, z176, z177, z178, z179,
    z180, z181, z182, z183, z184, z185, z186, z187, z188, z189, z190, z191,
    z192, z193, z194, z195, z196, z197, z198, z199, z200, z201, z202, z203,
    z204, z205, z206, z207, z208, z209, z210, z211, z212, z213, z214, z215,
    z216, z217, z218, z219, z220, z221, z222, z223, z224, z225, z226, z227,
    z228, z229, z230, z231, z232, z233, z234, z235, z236, z237, z238, z239,
    z240, z241, z242, z243, z244, z245, z246, z247, z248, z249, z250, z251,
    z252, z253, z254, z255, z256, z257, z258, z259, z260, z261, z262, z263,
    z264, z265, z266, z267, z268, z269, z270, z271, z272, z273, z274, z275,
    z276, z277, z278, z279, z280, z281, z282, z283, z284, z285, z286, z287,
    z288, z289, z290, z291, z292, z293, z294, z295, z296, z297, z298, z299,
    z300, z301, z302, z303, z304, z305, z306, z307, z308, z309, z310, z311,
    z312, z313, z314, z315, z316, z317, z318, z319, z320, z321, z322, z323,
    z324, z325, z326, z327, z328, z329, z330, z331, z332, z333, z334, z335,
    z336, z337, z338, z339, z340, z341, z342, z343, z344, z345, z346, z347,
    z348, z349, z350, z351, z352, z353, z354, z355, z356, z357, z358, z359,
    z360, z361, z362, z363, z364, z365, z366, z367, z368, z369, z370, z371,
    z372, z373, z374, z375, z376, z377, z378, z379, z380, z381, z382, z383,
    z384, z385, z386, z387, z388, z389, z390, z391, z392, z393, z394, z395,
    z396, z397, z398, z399, z400, z401, z402, z403, z404, z405, z406, z407,
    z408, z409, z410, z411, z412, z413, z414, z415, z416, z417, z418, z419,
    z420, z421, z422, z423, z424, z425, z426, z427, z428, z429, z430, z431,
    z432, z433, z434, z435, z436, z437, z438, z439, z440, z441, z442, z443,
    z444, z445, z446, z447, z448, z449, z450, z451, z452, z453, z454, z455,
    z456, z457, z458, z459, z460, z461, z462, z463, z464, z465, z466, z467,
    z468, z469, z470, z471, z472, z473, z474, z475, z476, z477, z478, z479,
    z480, z481, z482, z483, z484, z485, z486, z487, z488, z489, z490, z491,
    z492, z493, z494, z495, z496, z497, z498, z499, z500, z501, z502, z503,
    z504, z505, z506, z507, z508, z509, z510, z511, z512  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z000, z001, z002, z003, z004, z005, z006, z007, z008, z009, z010,
    z011, z012, z013, z014, z015, z016, z017, z018, z019, z020, z021, z022,
    z023, z024, z025, z026, z027, z028, z029, z030, z031, z032, z033, z034,
    z035, z036, z037, z038, z039, z040, z041, z042, z043, z044, z045, z046,
    z047, z048, z049, z050, z051, z052, z053, z054, z055, z056, z057, z058,
    z059, z060, z061, z062, z063, z064, z065, z066, z067, z068, z069, z070,
    z071, z072, z073, z074, z075, z076, z077, z078, z079, z080, z081, z082,
    z083, z084, z085, z086, z087, z088, z089, z090, z091, z092, z093, z094,
    z095, z096, z097, z098, z099, z100, z101, z102, z103, z104, z105, z106,
    z107, z108, z109, z110, z111, z112, z113, z114, z115, z116, z117, z118,
    z119, z120, z121, z122, z123, z124, z125, z126, z127, z128, z129, z130,
    z131, z132, z133, z134, z135, z136, z137, z138, z139, z140, z141, z142,
    z143, z144, z145, z146, z147, z148, z149, z150, z151, z152, z153, z154,
    z155, z156, z157, z158, z159, z160, z161, z162, z163, z164, z165, z166,
    z167, z168, z169, z170, z171, z172, z173, z174, z175, z176, z177, z178,
    z179, z180, z181, z182, z183, z184, z185, z186, z187, z188, z189, z190,
    z191, z192, z193, z194, z195, z196, z197, z198, z199, z200, z201, z202,
    z203, z204, z205, z206, z207, z208, z209, z210, z211, z212, z213, z214,
    z215, z216, z217, z218, z219, z220, z221, z222, z223, z224, z225, z226,
    z227, z228, z229, z230, z231, z232, z233, z234, z235, z236, z237, z238,
    z239, z240, z241, z242, z243, z244, z245, z246, z247, z248, z249, z250,
    z251, z252, z253, z254, z255, z256, z257, z258, z259, z260, z261, z262,
    z263, z264, z265, z266, z267, z268, z269, z270, z271, z272, z273, z274,
    z275, z276, z277, z278, z279, z280, z281, z282, z283, z284, z285, z286,
    z287, z288, z289, z290, z291, z292, z293, z294, z295, z296, z297, z298,
    z299, z300, z301, z302, z303, z304, z305, z306, z307, z308, z309, z310,
    z311, z312, z313, z314, z315, z316, z317, z318, z319, z320, z321, z322,
    z323, z324, z325, z326, z327, z328, z329, z330, z331, z332, z333, z334,
    z335, z336, z337, z338, z339, z340, z341, z342, z343, z344, z345, z346,
    z347, z348, z349, z350, z351, z352, z353, z354, z355, z356, z357, z358,
    z359, z360, z361, z362, z363, z364, z365, z366, z367, z368, z369, z370,
    z371, z372, z373, z374, z375, z376, z377, z378, z379, z380, z381, z382,
    z383, z384, z385, z386, z387, z388, z389, z390, z391, z392, z393, z394,
    z395, z396, z397, z398, z399, z400, z401, z402, z403, z404, z405, z406,
    z407, z408, z409, z410, z411, z412, z413, z414, z415, z416, z417, z418,
    z419, z420, z421, z422, z423, z424, z425, z426, z427, z428, z429, z430,
    z431, z432, z433, z434, z435, z436, z437, z438, z439, z440, z441, z442,
    z443, z444, z445, z446, z447, z448, z449, z450, z451, z452, z453, z454,
    z455, z456, z457, z458, z459, z460, z461, z462, z463, z464, z465, z466,
    z467, z468, z469, z470, z471, z472, z473, z474, z475, z476, z477, z478,
    z479, z480, z481, z482, z483, z484, z485, z486, z487, z488, z489, z490,
    z491, z492, z493, z494, z495, z496, z497, z498, z499, z500, z501, z502,
    z503, z504, z505, z506, z507, z508, z509, z510, z511, z512;
  wire n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n553, n554, n555, n556, n557, n558, n559,
    n560, n561, n562, n563, n564, n565, n566, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
    n585, n586, n587, n588, n590, n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
    n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628, n629, n631, n632, n633, n634,
    n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
    n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
    n659, n660, n661, n662, n663, n664, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n714, n715, n716, n717, n718, n719, n720, n721,
    n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
    n746, n747, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
    n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
    n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
    n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n795, n796,
    n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
    n809, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n832, n833, n834,
    n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
    n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866, n867, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n889, n890, n891, n892, n893, n894, n895, n896, n897,
    n898, n899, n900, n901, n902, n903, n904, n905, n907, n908, n909, n910,
    n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
    n923, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
    n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n948,
    n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
    n961, n962, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
    n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
    n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1047, n1048, n1049, n1050,
    n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076, n1078, n1079, n1080, n1081,
    n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
    n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
    n1123, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
    n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1152, n1153, n1154,
    n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
    n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1211, n1212, n1214, n1215, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
    n1250, n1252, n1253, n1254, n1255, n1256, n1258, n1259, n1260, n1261,
    n1262, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1273,
    n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
    n1284, n1285, n1286, n1287, n1288, n1290, n1291, n1292, n1293, n1294,
    n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1314, n1315,
    n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1367,
    n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
    n1388, n1389, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
    n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
    n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
    n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1450,
    n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
    n1471, n1472, n1473, n1474, n1476, n1477, n1478, n1479, n1480, n1481,
    n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
    n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1502,
    n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
    n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
    n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
    n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
    n1554, n1555, n1556, n1557, n1558, n1559, n1561, n1562, n1563, n1564,
    n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
    n1575, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1588, n1589, n1590, n1591, n1593, n1594, n1595, n1596, n1598,
    n1599, n1600, n1601, n1604, n1605, n1606, n1608, n1609, n1610, n1611,
    n1612, n1613, n1614, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
    n1623, n1624, n1625, n1626, n1627, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
    n1644, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
    n1655, n1656, n1657, n1658, n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
    n1676, n1677, n1678, n1679, n1681, n1682, n1683, n1684, n1685, n1686,
    n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
    n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1727, n1728,
    n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
    n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1752, n1754, n1755, n1756, n1757, n1758, n1759,
    n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
    n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1779, n1780,
    n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
    n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
    n1822, n1823, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
    n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
    n1843, n1844, n1845, n1846, n1847, n1848, n1850, n1851, n1852, n1853,
    n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
    n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1872, n1873, n1874,
    n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
    n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1893, n1894, n1895,
    n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1912, n1913, n1914, n1915, n1916,
    n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
    n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1937,
    n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
    n1958, n1959, n1960, n1961, n1962, n1964, n1965, n1966, n1967, n1968,
    n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
    n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
    n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
    n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
    n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2050, n2051, n2052,
    n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
    n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2072, n2073,
    n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
    n2084, n2085, n2086, n2087, n2088, n2089, n2091, n2092, n2093, n2094,
    n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
    n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
    n2126, n2127, n2128, n2129, n2131, n2132, n2133, n2134, n2135, n2136,
    n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
    n2147, n2148, n2149, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
    n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2167, n2168,
    n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
    n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
    n2189, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
    n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
    n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2239, n2240, n2241,
    n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
    n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
    n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
    n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2288, n2289, n2290, n2291, n2292, n2293,
    n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
    n2304, n2305, n2306, n2307, n2308, n2310, n2311, n2312, n2313, n2314,
    n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
    n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2334, n2335,
    n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
    n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2361, n2362, n2363, n2364, n2365, n2366,
    n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
    n2377, n2378, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
    n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2397, n2398,
    n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
    n2409, n2410, n2411, n2412, n2413, n2414, n2416, n2417, n2418, n2419,
    n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
    n2430, n2431, n2432, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
    n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
    n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2471, n2472,
    n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
    n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
    n2493, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
    n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
    n2514, n2515, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
    n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
    n2535, n2536, n2537, n2538, n2540, n2541, n2542, n2543, n2544, n2545,
    n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
    n2556, n2557, n2558, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
    n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
    n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
    n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
    n2598, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
    n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
    n2630, n2631, n2632, n2633, n2634, n2636, n2637, n2638, n2639, n2640,
    n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
    n2651, n2652, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
    n2662, n2663, n2664, n2665, n2666, n2667, n2669, n2670, n2671, n2672,
    n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
    n2683, n2684, n2685, n2686, n2688, n2689, n2690, n2691, n2692, n2693,
    n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2702, n2703, n2704,
    n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721, n2723, n2724, n2725, n2726,
    n2727, n2728, n2729, n2730, n2731, n2732, n2734, n2735, n2736, n2737,
    n2738, n2739, n2740, n2741, n2742, n2743, n2745, n2746, n2747, n2748,
    n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2757, n2758, n2759,
    n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2770,
    n2771, n2772, n2773, n2774, n2775, n2776, n2778, n2779, n2780, n2781,
    n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2792,
    n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
    n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
    n2813, n2814, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
    n2834, n2835, n2836, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
    n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2854, n2855,
    n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
    n2877, n2879, n2880, n2881, n2882, n2883, n2885, n2886, n2887, n2888,
    n2889, n2890, n2891, n2892, n2894, n2895, n2896, n2897, n2898, n2899,
    n2900, n2901, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2915, n2916, n2918, n2919, n2920, n2921,
    n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
    n2932, n2933, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
    n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
    n2953, n2954, n2955, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
    n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
    n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
    n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2994, n2995,
    n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
    n3006, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
    n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3027,
    n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
    n3038, n3039, n3040, n3041, n3042, n3044, n3045, n3046, n3047, n3048,
    n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
    n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3079, n3080,
    n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
    n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
    n3101, n3102, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
    n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
    n3122, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
    n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3143,
    n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
    n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3162, n3163, n3165,
    n3166, n3167, n3168, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
    n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3185, n3186, n3187,
    n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
    n3198, n3199, n3200, n3201, n3203, n3204, n3205, n3206, n3207, n3208,
    n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
    n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
    n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3239, n3240,
    n3241, n3242, n3243, n3244, n3245, n3246, n3248, n3249, n3250, n3251,
    n3252, n3253, n3254, n3255, n3256, n3257, n3259, n3260, n3261, n3262,
    n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3273,
    n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
    n3284, n3285, n3286, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
    n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
    n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
    n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
    n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
    n3337, n3338, n3339, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
    n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
    n3358, n3359, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
    n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
    n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
    n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3399, n3400,
    n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
    n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
    n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
    n3442, n3443, n3444, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
    n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
    n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3471, n3472, n3473,
    n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
    n3484, n3485, n3486, n3487, n3488, n3490, n3491, n3492, n3493, n3494,
    n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
    n3505, n3506, n3507, n3508, n3509, n3510, n3512, n3513, n3514, n3515,
    n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
    n3526, n3527, n3528, n3529, n3531, n3532, n3533, n3534, n3535, n3536,
    n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
    n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3557,
    n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
    n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
    n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3599,
    n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
    n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
    n3631, n3632, n3633, n3634, n3636, n3637, n3638, n3639, n3640, n3641,
    n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
    n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
    n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3671, n3672, n3673,
    n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
    n3684, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
    n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
    n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
    n3716, n3717, n3718, n3719, n3721, n3722, n3723, n3724, n3725, n3726,
    n3727, n3728, n3729, n3730, n3731, n3733, n3734, n3735, n3736, n3737,
    n3738, n3739, n3740, n3741, n3742, n3743, n3745, n3746, n3747, n3748,
    n3749, n3750, n3751, n3752, n3753, n3754, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765, n3767, n3768, n3769, n3770,
    n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3779, n3780, n3781,
    n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
    n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
    n3803, n3804, n3805, n3806, n3807, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
    n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
    n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
    n3846, n3847, n3848, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
    n3857, n3858, n3859, n3860, n3861, n3862, n3864, n3865, n3866, n3867,
    n3868, n3869, n3870, n3871, n3872, n3873, n3875, n3876, n3877, n3878,
    n3879, n3880, n3881, n3882, n3883, n3884, n3886, n3887, n3888, n3889,
    n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
    n3900, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
    n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
    n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
    n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3942,
    n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
    n3953, n3954, n3955, n3956, n3957, n3958, n3960, n3961, n3962, n3963,
    n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
    n3974, n3975, n3976, n3977, n3978, n3979, n3981, n3982, n3983, n3984,
    n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3994, n3995,
    n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
    n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4015, n4016,
    n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
    n4027, n4028, n4029, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
    n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
    n4048, n4049, n4050, n4051, n4052, n4054, n4055, n4056, n4057, n4058,
    n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
    n4069, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
    n4080, n4081, n4082, n4083, n4084, n4085, n4087, n4088, n4089, n4090,
    n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
    n4101, n4102, n4103, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
    n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
    n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
    n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4142, n4143,
    n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
    n4154, n4155, n4156, n4157, n4159, n4160, n4161, n4162, n4163, n4164,
    n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
    n4175, n4176, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
    n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
    n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
    n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
    n4217, n4218, n4219, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
    n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
    n4238, n4239, n4240, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
    n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
    n4259, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
    n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4278, n4279, n4280,
    n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
    n4291, n4292, n4293, n4294, n4296, n4297, n4298, n4299, n4300, n4301,
    n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
    n4312, n4313, n4314, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
    n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
    n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
    n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
    n4354, n4355, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
    n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
    n4375, n4376, n4377, n4378, n4379, n4380, n4382, n4383, n4384, n4385,
    n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
    n4396, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
    n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
    n4417, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
    n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
    n4438, n4439, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
    n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
    n4459, n4460, n4461, n4462, n4463, n4464, n4466, n4467, n4468, n4469,
    n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
    n4480, n4481, n4482, n4483, n4485, n4486, n4487, n4488, n4489, n4490,
    n4491, n4492, n4493, n4494, n4496, n4497, n4498, n4499, n4500, n4501,
    n4502, n4503, n4504, n4505, n4506, n4507, n4509, n4510, n4511, n4512,
    n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
    n4523, n4524, n4525, n4526, n4527, n4529, n4530, n4531, n4532, n4533,
    n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
    n4544, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
    n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4563, n4564, n4565,
    n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
    n4576, n4577, n4578, n4579, n4581, n4582, n4583, n4584, n4585, n4586,
    n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
    n4598, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
    n4609, n4611, n4612, n4613, n4614, n4616, n4617, n4618, n4619, n4620,
    n4621, n4622, n4623, n4625, n4626, n4627, n4630, n4631, n4632, n4634,
    n4635, n4636, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
    n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
    n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
    n4668, n4669, n4670, n4671, n4672, n4674, n4675, n4676, n4677, n4678,
    n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
    n4689, n4690, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
    n4710, n4711, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
    n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
    n4731, n4732, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
    n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
    n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
    n4763, n4764, n4765, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
    n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
    n4784, n4785, n4786, n4787, n4789, n4790, n4791, n4792, n4793, n4794,
    n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4803, n4804, n4805,
    n4806, n4807, n4808, n4809, n4810, n4811, n4813, n4814, n4816, n4817,
    n4818, n4819, n4820, n4822, n4823, n4824, n4825, n4826, n4828, n4829,
    n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4838, n4839, n4840,
    n4841, n4842, n4843, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
    n4852, n4853, n4854, n4855, n4857, n4858, n4859, n4860, n4861, n4862,
    n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
    n4873, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
    n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4892, n4893, n4894,
    n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
    n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4913, n4914, n4915,
    n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
    n4926, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
    n4937, n4938, n4939, n4940, n4941, n4943, n4944, n4945, n4946, n4947,
    n4948, n4949, n4950, n4951, n4953, n4954, n4955, n4956, n4957, n4958,
    n4959, n4960, n4961, n4962, n4963, n4965, n4966, n4967, n4968, n4969,
    n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
    n4980, n4981, n4982, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
    n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
    n5001, n5002, n5003, n5004, n5006, n5007, n5008, n5009, n5010, n5011,
    n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5022,
    n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
    n5033, n5034, n5035, n5036, n5038, n5039, n5040, n5041, n5042, n5043,
    n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5054,
    n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
    n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5074, n5075,
    n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
    n5086, n5087, n5088, n5089, n5090, n5092, n5093, n5094, n5095, n5096,
    n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
    n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
    n5118, n5119, n5120, n5121, n5123, n5124, n5125, n5126, n5127, n5128,
    n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5139,
    n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
    n5150, n5151, n5152, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
    n5161, n5162, n5163, n5164, n5166, n5167, n5168, n5169, n5170, n5171,
    n5172, n5173, n5174, n5175, n5176, n5178, n5179, n5180, n5181, n5182,
    n5183, n5185, n5186, n5187, n5188, n5189, n5191, n5192, n5193, n5194,
    n5195, n5196, n5197, n5198, n5200, n5201, n5202, n5203, n5204, n5205,
    n5206, n5207, n5208, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
    n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
    n5227, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
    n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5248,
    n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
    n5269, n5270, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
    n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
    n5290, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
    n5301, n5302, n5303, n5304, n5305, n5306, n5308, n5309, n5310, n5311,
    n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
    n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5330, n5331, n5332,
    n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
    n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5351, n5352, n5353,
    n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
    n5364, n5365, n5366, n5367, n5368, n5369, n5371, n5372, n5373, n5374,
    n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
    n5385, n5386, n5387, n5388, n5389, n5390, n5392, n5393, n5394, n5395,
    n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
    n5406, n5407, n5408, n5409, n5410, n5411, n5413, n5414, n5415, n5416,
    n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
    n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5436, n5437,
    n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
    n5448, n5449, n5450, n5451, n5452, n5453, n5455, n5456, n5457, n5458,
    n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
    n5469, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
    n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5488, n5489, n5490,
    n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
    n5501, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
    n5512, n5513, n5514, n5515, n5516, n5518, n5519, n5520, n5521, n5522,
    n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
    n5533, n5534, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
    n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
    n5554, n5555, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
    n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
    n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
    n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
    n5596, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
    n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5617,
    n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
    n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5636, n5637, n5638,
    n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
    n5649, n5650, n5651, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
    n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
    n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
    n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5689, n5690, n5691,
    n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5701, n5702,
    n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
    n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5723,
    n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
    n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5743, n5744,
    n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
    n5755, n5756, n5757, n5758, n5760, n5761, n5762, n5763, n5764, n5765,
    n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5775, n5776,
    n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
    n5787, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5797, n5798,
    n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
    n5809, n5810, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
    n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5828, n5829, n5830,
    n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
    n5841, n5842, n5843, n5844, n5845, n5846, n5848, n5849, n5850, n5851,
    n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
    n5862, n5863, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
    n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
    n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
    n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5903, n5904,
    n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5915,
    n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5926,
    n5927, n5928, n5929, n5930, n5931, n5932, n5934, n5935, n5936, n5937,
    n5939, n5940, n5941, n5942, n5943, n5944, n5946, n5947, n5948, n5949,
    n5950, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5961,
    n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
    n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
    n5983, n5984, n5985, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
    n5994, n5995, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
    n6005, n6006, n6008, n6009, n6010, n6011, n6012, n6013, n6015, n6016,
    n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
    n6027, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
    n6038, n6039, n6040, n6041, n6042, n6043, n6045, n6046, n6047, n6048,
    n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
    n6059, n6060, n6061, n6062, n6063, n6065, n6066, n6067, n6068, n6069,
    n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6080,
    n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
    n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
    n6102, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
    n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6121, n6122, n6123,
    n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
    n6134, n6135, n6136, n6137, n6138, n6139, n6141, n6142, n6143, n6144,
    n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
    n6155, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
    n6166, n6167, n6168, n6169, n6171, n6172, n6173, n6174, n6175, n6176,
    n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
    n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
    n6198, n6199, n6200, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
    n6209, n6210, n6211, n6212, n6214, n6215, n6216, n6217, n6218, n6219,
    n6220, n6222, n6223, n6224, n6225, n6226, n6227, n6229, n6230, n6231,
    n6232, n6233, n6234, n6235, n6236, n6238, n6239, n6240, n6242, n6243,
    n6244, n6245, n6246, n6247, n6249, n6250, n6251, n6252, n6253, n6254,
    n6255, n6256, n6257, n6258, n6259, n6260, n6262, n6263, n6264, n6265,
    n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
    n6276, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
    n6287, n6288, n6289, n6290, n6291, n6292, n6294, n6295, n6296, n6297,
    n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
    n6308, n6309, n6310, n6311, n6313, n6314, n6315, n6316, n6317, n6318,
    n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
    n6329, n6330, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
    n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6348, n6349, n6350,
    n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
    n6361, n6362, n6363, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
    n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6381, n6382,
    n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
    n6393, n6394, n6395, n6396, n6398, n6399, n6400, n6401, n6402, n6403,
    n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
    n6414, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
    n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
    n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
    n6446, n6447, n6448, n6449, n6450, n6452, n6453, n6454, n6455, n6456,
    n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6466, n6467,
    n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
    n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6486, n6487, n6488,
    n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
    n6499, n6500, n6501, n6502, n6504, n6505, n6506, n6507, n6508, n6509,
    n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
    n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
    n6531, n6532, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
    n6542, n6543, n6544, n6545, n6546, n6547, n6549, n6550, n6551, n6552,
    n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
    n6563, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
    n6574, n6575, n6576, n6577, n6578, n6579, n6581, n6582, n6583, n6584,
    n6585, n6586, n6587, n6589, n6590, n6591, n6592, n6593, n6594, n6596,
    n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
    n6607, n6608, n6609, n6610, n6612, n6613, n6614, n6615, n6616, n6617,
    n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6626, n6627, n6628,
    n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
    n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6648, n6649, n6650,
    n6651, n6652, n6653, n6654, n6656, n6657, n6658, n6659, n6660, n6661,
    n6662, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
    n6673, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6684,
    n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6693, n6694, n6695,
    n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
    n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
    n6717, n6718, n6719, n6720, n6722, n6723, n6724, n6725, n6726, n6727,
    n6728, n6729, n6730, n6731, n6732, n6733, n6735, n6736, n6737, n6738,
    n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
    n6749, n6750, n6751, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
    n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6769, n6770,
    n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
    n6781, n6782, n6783, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
    n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6800, n6801, n6802,
    n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
    n6813, n6814, n6815, n6816, n6818, n6819, n6820, n6821, n6822, n6823,
    n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
    n6834, n6835, n6836, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
    n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
    n6855, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
    n6866, n6867, n6868, n6869, n6870, n6872, n6873, n6874, n6875, n6876,
    n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
    n6887, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
    n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6908,
    n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
    n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6928, n6929,
    n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
    n6940, n6941, n6942, n6943, n6945, n6946, n6947, n6948, n6949, n6950,
    n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
    n6961, n6962, n6963, n6964, n6966, n6967, n6969, n6970, n6971, n6972,
    n6973, n6974, n6975, n6976, n6977, n6979, n6980, n6981, n6982, n6983,
    n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
    n6994, n6995, n6996, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
    n7005, n7006, n7007, n7008, n7009, n7010, n7012, n7013, n7014, n7015,
    n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
    n7026, n7027, n7028, n7029, n7031, n7032, n7033, n7034, n7035, n7036,
    n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
    n7047, n7048, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
    n7058, n7059, n7060, n7061, n7062, n7064, n7065, n7066, n7067, n7068,
    n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
    n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
    n7090, n7091, n7092, n7093, n7094, n7095, n7097, n7098, n7099, n7100,
    n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
    n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
    n7122, n7123, n7124, n7125, n7126, n7127, n7129, n7130, n7131, n7132,
    n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
    n7143, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
    n7154, n7155, n7156, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
    n7165, n7166, n7167, n7168, n7169, n7171, n7172, n7173, n7174, n7175,
    n7176, n7177, n7178, n7179, n7181, n7182, n7183, n7184, n7185, n7186,
    n7187, n7188, n7189, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
    n7198, n7199, n7201, n7202, n7203, n7204, n7205, n7207, n7208, n7209,
    n7210, n7211, n7212, n7214, n7215, n7217, n7219, n7220, n7221, n7223,
    n7224, n7225, n7226, n7227, n7229, n7230, n7231, n7232, n7233, n7234,
    n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7244, n7245, n7246,
    n7247, n7248, n7249, n7251, n7252, n7253, n7254, n7255, n7256, n7258,
    n7259, n7260, n7261, n7263, n7264, n7265, n7266, n7268, n7269, n7270,
    n7271, n7272, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
    n7282, n7283, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
    n7293, n7294, n7295, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
    n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
    n7314, n7315, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
    n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
    n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
    n7346, n7347, n7348, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
    n7357, n7358, n7359, n7360, n7361, n7362, n7364, n7365, n7366, n7367,
    n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
    n7378, n7379, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
    n7389, n7390, n7391, n7392, n7393, n7394, n7397, n7398, n7399, n7400,
    n7401, n7402, n7403, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
    n7412, n7413, n7414, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
    n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7433,
    n7434, n7435, n7437, n7438, n7439, n7440, n7441, n7442, n7444, n7445,
    n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
    n7456, n7457, n7458, n7459, n7460, n7462, n7463, n7464, n7465, n7466,
    n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
    n7477, n7478, n7479, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
    n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7498,
    n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
    n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7518, n7519,
    n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
    n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7538, n7539, n7540,
    n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
    n7551, n7552, n7553, n7554, n7555, n7557, n7558, n7559, n7560, n7561,
    n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
    n7572, n7573, n7574, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
    n7583, n7584, n7585, n7586, n7587, n7588, n7590, n7591, n7592, n7593,
    n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
    n7604, n7605, n7606, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
    n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7623, n7624, n7625,
    n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
    n7636, n7637, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
    n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7656, n7657,
    n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
    n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
    n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
    n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7697, n7698, n7699,
    n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
    n7710, n7711, n7712, n7713, n7715, n7716, n7717, n7718, n7719, n7720,
    n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7731,
    n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
    n7742, n7743, n7744, n7745, n7746, n7747, n7749, n7750, n7751, n7752,
    n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7762, n7763,
    n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
    n7774, n7775, n7776, n7777, n7778, n7779, n7781, n7782, n7783, n7784,
    n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
    n7795, n7796, n7797, n7798, n7799, n7801, n7802, n7803, n7804, n7805,
    n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
    n7816, n7817, n7818, n7819, n7821, n7822, n7823, n7824, n7825, n7826,
    n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
    n7837, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
    n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
    n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
    n7869, n7870, n7871, n7872, n7873, n7874, n7876, n7877, n7878, n7879,
    n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
    n7890, n7891, n7892, n7893, n7895, n7896, n7897, n7898, n7899, n7900,
    n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
    n7911, n7912, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
    n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
    n7932, n7933, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
    n7943, n7944, n7945, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
    n7954, n7955, n7956, n7957, n7958, n7959, n7961, n7962, n7963, n7964,
    n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
    n7975, n7976, n7977, n7978, n7980, n7981, n7982, n7983, n7984, n7985,
    n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
    n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
    n8007, n8008, n8009, n8010, n8011, n8012, n8014, n8015, n8016, n8017,
    n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
    n8028, n8029, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
    n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8048, n8049,
    n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
    n8060, n8061, n8062, n8063, n8064, n8066, n8067, n8068, n8069, n8070,
    n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8081,
    n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
    n8092, n8093, n8094, n8095, n8096, n8097, n8099, n8100, n8101, n8102,
    n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
    n8113, n8114, n8115, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
    n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8132, n8133, n8134,
    n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
    n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
    n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8165, n8166,
    n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
    n8177, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
    n8188, n8189, n8190, n8191, n8192, n8193, n8195, n8196, n8197, n8198,
    n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8209,
    n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8220,
    n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
    n8231, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
    n8242, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
    n8253, n8254, n8255, n8256, n8258, n8259, n8260, n8261, n8262, n8263,
    n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8274,
    n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
    n8285, n8286, n8287, n8288, n8289, n8291, n8292, n8293, n8294, n8295,
    n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
    n8306, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
    n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
    n8327, n8328, n8329, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
    n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8348,
    n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
    n8359, n8360, n8361, n8362, n8363, n8364, n8366, n8367, n8368, n8369,
    n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8379, n8380,
    n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
    n8391, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400;
  assign z034 = 1'b0;
  assign z000 = ~x2 & (~n531 | (~x3 & (n523 | n528)));
  assign n523 = n527 & ((~x0 & ~n524) | (n525 & n526));
  assign n524 = x4 ? (~x5 | x7) : (x5 | ~x7);
  assign n525 = x0 & x4;
  assign n526 = x5 & x7;
  assign n527 = ~x1 & ~x6;
  assign n528 = n529 & n530;
  assign n529 = ~x4 & ~x0 & x1;
  assign n530 = x7 & x5 & x6;
  assign n531 = ~n533 & (x1 | n532);
  assign n532 = x0 ? ((~x3 | (x4 & (x5 | x6))) & (x3 | ~x4 | ~x5 | ~x6)) : (x3 | (x5 ? x4 : (~x4 & ~x6)));
  assign n533 = ~x0 & x1 & (x3 ? (~x4 & ~x5) : x4);
  assign z001 = n546 | n542 | n535 | n540;
  assign n535 = ~x1 & ((n536 & ~n537) | (~n538 & n539));
  assign n536 = x0 & x3;
  assign n537 = (~x2 | x4 | ~x5 | x6) & (x2 | ~x4 | x5 | ~x6);
  assign n538 = x2 ? (x5 | x6) : (~x5 | ~x6);
  assign n539 = x4 & ~x0 & ~x3;
  assign n540 = ~x1 & ~n541;
  assign n541 = x2 ? ((x3 | x4) & (~x0 | (x3 & (x4 | x5)))) : (~x3 | (x0 & (~x4 | ~x5)));
  assign n542 = n543 & (~n544 | n545);
  assign n543 = ~x0 & x1;
  assign n544 = x2 ? x3 : (~x3 | ~x4);
  assign n545 = x5 & ~x4 & ~x2 & x3;
  assign n546 = n551 & ((n549 & n550) | (n547 & n548));
  assign n547 = ~x3 & ~x0 & ~x2;
  assign n548 = x7 & x4 & ~x6;
  assign n549 = x3 & x0 & x2;
  assign n550 = ~x7 & ~x4 & x6;
  assign n551 = ~x1 & x5;
  assign z002 = ~n553 | n556 | n562 | (n560 & n561);
  assign n553 = x1 ? n555 : n554;
  assign n554 = (~x2 | ((~x0 | (~x3 ^ ~x4)) & (~x4 | ~x5 | x0 | x3))) & (~x3 | (x0 ? (~x4 | ~x5) : (x4 & (x2 | x5))));
  assign n555 = (x2 | ((x0 | ~x3 | ~x5) & (x4 | x5 | ~x0 | x3))) & (x0 | ~x3 | (x5 ? x4 : (~x2 & ~x4)));
  assign n556 = ~x0 & ((x2 & ~n557) | (n558 & n559));
  assign n557 = (~x1 | x6 | (x3 ? (~x4 | ~x5) : (x4 | x5))) & (x1 | x3 | ~x4 | x5 | ~x6);
  assign n558 = ~x3 & ~x1 & ~x2;
  assign n559 = x6 & x4 & x5;
  assign n560 = ~x2 & x0 & ~x1;
  assign n561 = x6 & ~x5 & x3 & x4;
  assign n562 = x5 & ((~n563 & n564) | (~n565 & n566));
  assign n563 = (~x1 | x2 | x3 | x6 | x7) & (x1 | ~x2 | ~x3 | ~x6 | ~x7);
  assign n564 = x0 & ~x4;
  assign n565 = (~x1 | ~x2 | ~x3 | ~x6 | x7) & (x1 | x2 | x3 | x6 | ~x7);
  assign n566 = ~x0 & x4;
  assign z003 = n574 | ~n578 | (~x3 & ~n568);
  assign n568 = (n571 | ~n572) & (~n569 | ~n570 | n573);
  assign n569 = x6 & ~x7;
  assign n570 = ~x1 & x2;
  assign n571 = (x4 | ((x0 | (x1 ? (~x5 | ~x6) : (x5 | x6))) & (~x0 | ~x1 | ~x5 | x6))) & (x1 | ~x4 | ~x5 | x6);
  assign n572 = ~x2 & x7;
  assign n573 = x0 ? (~x4 | ~x5) : (x4 | x5);
  assign n574 = x0 & ((n576 & n577) | (~x1 & ~n575));
  assign n575 = (x2 | (~x4 ^ ~x6) | (~x3 ^ x5)) & (~x2 | ~x4 | ~x5 | x6);
  assign n576 = ~x3 & x1 & ~x2;
  assign n577 = x6 & ~x4 & x5;
  assign n578 = ~n579 & n584 & (x2 ? n583 : n582);
  assign n579 = ~x0 & ((~x5 & ~n580) | (~x1 & n581));
  assign n580 = x1 ? ((x2 | ~x3 | ~x4 | x6) & (~x2 | x3 | x4 | ~x6)) : (x3 | (x2 ? (~x4 ^ ~x6) : (x4 | ~x6)));
  assign n581 = ~x2 & ~x3 & x5 & (x4 ^ ~x6);
  assign n582 = x3 ? ((x0 | x4 | (~x1 ^ ~x5)) & (x1 | ~x4 | ~x5)) : (x5 | ((~x1 | ~x4) & (~x0 | x1 | x4)));
  assign n583 = (x0 & (~x4 | x5)) | (~x1 & ~x4) | (x1 & x4) | (~x0 & ~x3 & ~x5);
  assign n584 = (n585 | n586) & (~n587 | ~n588);
  assign n585 = (~x2 | ((~x6 | ~x7 | ~x3 | ~x5) & (x6 | x7 | x3 | x5))) & (x2 | ~x3 | x5 | ~x6 | x7);
  assign n586 = x0 ? (x1 | x4) : (~x1 | ~x4);
  assign n587 = x3 & x2 & ~x0 & ~x1;
  assign n588 = ~x7 & ~x6 & ~x4 & ~x5;
  assign z004 = n611 | ~n614 | (x1 ? ~n602 : ~n590);
  assign n590 = ~n591 & ~n595 & (~n600 | ~n601);
  assign n591 = ~x7 & ((n592 & n594) | (x2 & ~n593));
  assign n592 = x6 & x4 & ~x5;
  assign n593 = (~x5 | ((~x0 | (x3 ? (~x4 | ~x6) : (x4 | x6))) & (x0 | ~x3 | x4 | x6))) & (x0 | ~x3 | ~x4 | x5 | x6);
  assign n594 = x3 & x0 & ~x2;
  assign n595 = ~n599 & ((n596 & n597) | (~x2 & n598));
  assign n596 = x2 & ~x3;
  assign n597 = x4 & x6;
  assign n598 = ~x6 & (x3 ^ x4);
  assign n599 = x0 ? (~x5 | ~x7) : (x5 | x7);
  assign n600 = ~x3 & x0 & ~x2;
  assign n601 = x7 & x6 & ~x4 & x5;
  assign n602 = ~n609 & (x0 | (~n603 & (~n607 | ~n608)));
  assign n603 = x7 & (n606 | (~n604 & ~n605));
  assign n604 = x3 ? (~x4 | ~x6) : (x4 | x6);
  assign n605 = x2 ^ x5;
  assign n606 = ~x6 & x5 & x4 & ~x2 & ~x3;
  assign n607 = ~x7 & (x4 ^ ~x5);
  assign n608 = x6 & ~x2 & ~x3;
  assign n609 = n600 & n610;
  assign n610 = ~x7 & ~x6 & x4 & x5;
  assign n611 = ~x2 & (x0 ? ~n612 : ~n613);
  assign n612 = (x3 | ((~x1 | x6 | (~x5 ^ ~x7)) & (~x6 | x7 | x1 | ~x5))) & (x1 | ~x3 | (x5 ? (x6 | x7) : (~x6 | ~x7)));
  assign n613 = (x3 | ((~x1 | (x5 ? (~x6 | ~x7) : (x6 | x7))) & (x6 | ~x7 | x1 | x5))) & (x1 | ~x3 | ~x5 | ~x6 | x7);
  assign n614 = ~n617 & ~n621 & n625 & (n615 | n616);
  assign n615 = x3 ? (x4 | ~x6) : (~x4 | x6);
  assign n616 = (x0 | ((~x1 | (x2 ? (x5 | ~x7) : (~x5 | x7))) & (~x5 | ~x7 | x1 | x2))) & (~x2 | x5 | x7 | ~x0 | x1);
  assign n617 = x2 & ((~n618 & n619) | (~x0 & n620));
  assign n618 = x0 ? (x3 ? (~x5 | ~x6) : (x5 | x6)) : (x5 | (~x3 ^ x6));
  assign n619 = ~x1 & x7;
  assign n620 = x1 & ~x7 & (x3 ? (~x5 & x6) : (x5 & ~x6));
  assign n621 = ~x2 & ((n622 & ~n623) | (n543 & n624));
  assign n622 = x0 & ~x3;
  assign n623 = x1 ? (~x5 | ~x6) : (x5 | x6);
  assign n624 = ~x6 & x3 & x5;
  assign n625 = (n627 | n628) & (~n626 | ~n629);
  assign n626 = ~x0 & ~x1;
  assign n627 = x3 ^ ~x6;
  assign n628 = (~x0 | x1 | ~x2 | x5) & (x0 | (x1 ? (~x2 | x5) : (x2 | ~x5)));
  assign n629 = x2 & (x3 ? (~x5 & x6) : (x5 & ~x6));
  assign z005 = n638 | n642 | ~n648 | (~x3 & ~n631);
  assign n631 = ~n636 & (x6 | (~n633 & (~n632 | ~n635)));
  assign n632 = x1 & ~x2;
  assign n633 = ~x4 & ~n634;
  assign n634 = (x0 | ~x1 | x2 | ~x5 | x7) & (x1 | ((~x5 | x7 | x0 | ~x2) & (~x0 | (x2 ? (~x5 | ~x7) : (x5 | x7)))));
  assign n635 = x7 & x4 & ~x5;
  assign n636 = n569 & ~n637;
  assign n637 = (x0 | ~x2 | ~x5 | (~x1 ^ x4)) & (x1 | x2 | ~x4 | x5);
  assign n638 = ~n640 & (x0 ? (n570 & n639) : ~n641);
  assign n639 = x5 & x3 & ~x4;
  assign n640 = x6 ^ x7;
  assign n641 = (x2 | ((~x1 | x4 | (~x3 ^ ~x5)) & (~x4 | ~x5 | x1 | ~x3))) & (x1 | ~x2 | x3 | x4 | x5);
  assign n642 = ~n643 & (~n644 | n645);
  assign n643 = x6 ^ ~x7;
  assign n644 = (x0 | ~x2 | (x1 ? (x3 | ~x4) : (~x3 | x4))) & (~x0 | ~x1 | x2 | x3 | x4);
  assign n645 = ~x1 & (x0 ? ~n646 : (~x2 & ~n647));
  assign n646 = (x4 | x5 | ~x2 | x3) & (~x4 | ~x5 | x2 | ~x3);
  assign n647 = x3 ? (x4 | x5) : (~x4 | ~x5);
  assign n648 = ~n663 & ~n660 & ~n656 & ~n649 & ~n652;
  assign n649 = ~x2 & (~n651 | (x3 & ~n650));
  assign n650 = (x0 | ~x1 | ~x4 | ~x5 | ~x6) & (x1 | (~x4 ^ x5) | (~x0 ^ ~x6));
  assign n651 = (~x1 | x6 | (x3 ? (x4 | x5) : (~x4 | ~x5))) & (x1 | x3 | x4 | ~x6);
  assign n652 = x2 & (~n655 | (x6 & n653 & ~n654));
  assign n653 = ~x0 & ~x3;
  assign n654 = x1 ? (x4 | x5) : (x4 ^ ~x5);
  assign n655 = (x0 | ~x1 | ~x3 | x4 | x6) & (x1 | ~x4 | (x0 ? (~x3 ^ ~x6) : (~x3 | x6)));
  assign n656 = x3 & ((n657 & n658) | (~n586 & n659));
  assign n657 = x4 & ~x0 & x1;
  assign n658 = ~x7 & x5 & ~x6;
  assign n659 = ~x5 & (x6 ^ ~x7);
  assign n660 = n661 & n662;
  assign n661 = ~x3 & x0 & ~x1;
  assign n662 = x7 & x6 & x4 & x5;
  assign n663 = n662 & n664;
  assign n664 = x3 & x2 & ~x0 & x1;
  assign z006 = ~n666 | (~n685 & n686) | (~x2 & ~n677);
  assign n666 = ~n667 & n673 & (n671 | n672);
  assign n667 = ~x0 & ((x1 & ~n668) | (n669 & n670));
  assign n668 = (~x2 | (~x4 ^ ~x7) | (~x3 & x5)) & (~x3 | ~x7 | ((~x4 | x5) & (x2 | x4 | ~x5)));
  assign n669 = x3 & ~x1 & ~x2;
  assign n670 = ~x7 & x4 & ~x5;
  assign n671 = x4 ^ ~x7;
  assign n672 = (~x1 | x2 | x3 | ~x5) & (x1 | ((~x2 | (~x3 & x5)) & (~x0 | ~x3 | x5)));
  assign n673 = (x2 | n675) & (~n674 | ~n676);
  assign n674 = ~x7 & x4 & x5;
  assign n675 = (~x5 | ~x7 | x1 | ~x4) & (x4 | (x1 ? (x5 | (x3 ^ ~x7)) : (~x5 | x7)));
  assign n676 = ~x3 & ~x1 & x2;
  assign n677 = ~n680 & (~x4 | (~n679 & (x7 | n678)));
  assign n678 = x1 ? (~x6 | ((x3 | x5) & (x0 | ~x3 | ~x5))) : (x6 | ((x3 | x5) & (~x0 | ~x3 | ~x5)));
  assign n679 = ~x3 & ~x5 & x7 & (~x1 ^ ~x6);
  assign n680 = n681 & ((~n682 & n683) | (n626 & n684));
  assign n681 = ~x4 & ~x5;
  assign n682 = x1 ^ ~x6;
  assign n683 = ~x3 & ~x7;
  assign n684 = x7 & x3 & ~x6;
  assign n685 = ((~x4 ^ ~x7) | ((x1 | ~x6) & (x0 | ~x1 | x6))) & (x4 | ~x7 | (x0 ? (x1 | x6) : (~x1 | ~x6)));
  assign n686 = x5 & x2 & ~x3;
  assign z007 = n688 | n695 | ~n703 | (n622 & ~n700);
  assign n688 = ~x0 & (n690 | (x5 & n689 & ~n694));
  assign n689 = ~x1 & ~x3;
  assign n690 = x1 & (x6 ? ~n692 : (n691 & ~n693));
  assign n691 = ~x2 & x5;
  assign n692 = (~x2 | ((x3 | ~x4 | ~x5 | ~x7) & (~x3 | x4 | x5 | x7))) & (x2 | x3 | ~x4 | ~x5 | x7);
  assign n693 = x3 ? (~x4 | ~x7) : (x4 | x7);
  assign n694 = (~x2 | ~x7 | (~x4 ^ ~x6)) & (x2 | ~x4 | ~x6 | x7);
  assign n695 = ~n697 & ((n696 & n699) | (~x1 & ~n698));
  assign n696 = ~x6 & ~x4 & ~x5;
  assign n697 = x2 ^ ~x7;
  assign n698 = (x5 | x6 | x3 | x4) & (~x3 | ((~x0 | ~x4 | ~x5 | x6) & (x5 | ~x6 | x0 | x4)));
  assign n699 = ~x3 & ~x0 & x1;
  assign n700 = (x2 | n701) & (x1 | ~x2 | ~x4 | ~n702);
  assign n701 = (~x4 | ~x5 | ~x6 | x7) & (~x1 | x4 | x5 | x6 | ~x7);
  assign n702 = x6 & (~x5 ^ x7);
  assign n703 = x2 ? (~n709 & (~n704 | ~n712)) : n705;
  assign n704 = x6 & ~x4 & ~x5;
  assign n705 = n708 & (~n706 | n707);
  assign n706 = x5 & ~x6;
  assign n707 = (~x0 | x1 | ~x3 | x4) & (x0 | ~x1 | (~x3 ^ x4));
  assign n708 = (x3 | x5 | ~x6) & (~x5 | ((x0 | (x6 ? ~x3 : x1)) & (x1 | ~x3 | ~x6) & (~x0 | x3 | x6)));
  assign n709 = ~n710 & ~n711;
  assign n710 = x0 & x1;
  assign n711 = (x5 | ((~x4 | x6) & (~x3 | (~x4 & x6)))) & (x3 | x4 | ~x5 | ~x6);
  assign n712 = x3 & x0 & ~x1;
  assign z008 = n715 | ~n721 | ~n735 | (~n714 & ~n734);
  assign n714 = x4 ^ ~x5;
  assign n715 = ~x1 & (n716 | (n719 & n720));
  assign n716 = x6 & ((n600 & n717) | (~x5 & ~n718));
  assign n717 = x7 & x4 & x5;
  assign n718 = (~x0 | ~x4 | (x2 ? (x3 | ~x7) : (~x3 | x7))) & (x0 | ~x2 | ~x3 | x4 | ~x7);
  assign n719 = x5 & ~x6 & (~x3 ^ ~x7);
  assign n720 = ~x4 & ~x0 & x2;
  assign n721 = n722 & (n643 | n729) & (x2 | n725);
  assign n722 = (n524 | n723) & (x1 | n724);
  assign n723 = x1 ? ((x2 | x3 | x6) & (x0 | ((x3 | x6) & (~x2 | ~x3 | ~x6)))) : ((~x3 | ~x6 | x0 | x2) & (x3 | x6 | ~x0 | ~x2));
  assign n724 = (~x4 | x6 | x0 | ~x3) & (~x0 | x4 | (x2 ? (x3 | ~x6) : (~x3 | x6)));
  assign n725 = (~n727 | ~n728) & (x5 | ~n525 | n726);
  assign n726 = x1 ? (x3 | ~x6) : (~x3 | x6);
  assign n727 = x3 & ~x0 & ~x1;
  assign n728 = ~x6 & ~x4 & x5;
  assign n729 = (~n731 | ~n733) & (x1 | (~n730 & n732));
  assign n730 = ~x5 & ~x4 & ~x3 & x0 & ~x2;
  assign n731 = x5 & x3 & x4;
  assign n732 = (x4 | x5 | x0 | x3) & (~x4 | ~x5 | ~x0 | ~x3);
  assign n733 = ~x2 & ~x0 & x1;
  assign n734 = (x0 | ((x3 | ~x6) & (~x1 | x2 | ~x3 | x6))) & (x1 | ((x2 | x3 | ~x6) & (~x0 | ~x2 | ~x3 | x6)));
  assign n735 = ~n736 & ~n739 & ~n741 & (~n746 | ~n747);
  assign n736 = ~n737 & n738;
  assign n737 = (x2 | ~x5 | x6 | ~x7) & (x5 | ~x6 | x7);
  assign n738 = ~x4 & ~x3 & ~x0 & x1;
  assign n739 = ~n740 & (~x0 | (x1 & ~x2) | (~x1 & x2));
  assign n740 = (~x3 | x4 | x5 | x6 | x7) & (x3 | ~x4 | ~x5 | ~x6 | ~x7);
  assign n741 = x1 & ((n743 & n744) | (n742 & n745));
  assign n742 = ~x0 & x2;
  assign n743 = x0 & ~x2;
  assign n744 = x6 & ~x3 & ~x4;
  assign n745 = ~x6 & x3 & x4;
  assign n746 = x2 & ~x0 & x1;
  assign n747 = ~x6 & x5 & x3 & ~x4;
  assign z009 = ~n763 | (x0 ? (n756 | n760) : ~n749);
  assign n749 = ~n751 & (~n750 | n755);
  assign n750 = x5 & ~x7;
  assign n751 = x7 & ((~n752 & ~n753) | (x5 & ~n754));
  assign n752 = x3 ? (x4 | x6) : (~x4 | ~x6);
  assign n753 = x1 ? (x2 | x5) : (~x2 | ~x5);
  assign n754 = (~x1 | x2 | x3 | x4 | x6) & (x1 | ((~x3 | ~x4 | ~x6) & (~x2 | x3 | x4 | x6)));
  assign n755 = (~x1 | ~x2 | ~x3 | ~x4 | x6) & (x1 | (x4 ? (x6 | (x2 & x3)) : ~x6));
  assign n756 = ~x1 & ((~x7 & ~n758) | (n757 & ~n759));
  assign n757 = ~x5 & x7;
  assign n758 = (x2 & (x5 | (x3 & ~x6))) | (~x4 & ~x6) | (x3 & x5) | (x4 & x6) | (~x2 & ~x3 & ~x5);
  assign n759 = (~x2 | (~x4 ^ ~x6)) & (~x3 | ~x4 | ~x6);
  assign n760 = n757 & n632 & (n761 | n762);
  assign n761 = ~x6 & x3 & ~x4;
  assign n762 = ~x3 & (x4 ^ ~x6);
  assign n763 = x4 ? (~n764 & (x1 | n766)) : n767;
  assign n764 = ~n765 & ((~x0 & x1) | (~x2 & ~x3) | (x2 & x3 & x0 & ~x1));
  assign n765 = x5 ^ x7;
  assign n766 = x0 ? (~x5 | ~x7 | (x2 ^ ~x3)) : (x7 | ((~x3 | x5) & (~x2 | (~x3 & x5))));
  assign n767 = ~n768 & ~n769 & (x2 | n770);
  assign n768 = ~x0 & ((~x1 & ~x5 & x7) | (x2 & ((~x5 & x7) | (x1 & x5 & ~x7))));
  assign n769 = ~x7 & x5 & x2 & x0 & ~x1;
  assign n770 = ((~x0 ^ x1) | (x3 ? (~x5 | x7) : (x5 | ~x7))) & (~x0 | ~x1 | x3 | ~x5 | x7);
  assign z010 = n773 | n780 | n786 | (n772 & ~n789);
  assign n772 = ~x1 & x4;
  assign n773 = x1 & (n775 | (n774 & n743 & n779));
  assign n774 = x3 & ~x4;
  assign n775 = ~x0 & ((~n777 & n778) | (~x6 & ~n776));
  assign n776 = x2 ? (~x3 | x7 | (~x4 ^ ~x5)) : (x3 | (~x4 ^ x5));
  assign n777 = (x5 | (x3 ? (~x4 | ~x7) : (~x4 ^ x7))) & (x3 | x4 | ~x5 | x7);
  assign n778 = ~x2 & x6;
  assign n779 = ~x5 & (~x6 | ~x7);
  assign n780 = x3 & (n781 | ~n783 | (~x1 & ~n782));
  assign n781 = ~x1 & (x0 ? (x2 ? (~x5 & ~x6) : (x5 & x6)) : ((~x5 & x6) | (x2 & x5 & ~x6)));
  assign n782 = x0 ? ((~x6 | ~x7 | ~x2 | ~x5) & (x6 | x7 | x2 | x5)) : (x2 | x6 | (~x5 ^ x7));
  assign n783 = x5 | ~n543 | (n784 & n785);
  assign n784 = x2 ^ x6;
  assign n785 = x2 ? (x6 | ~x7) : (~x6 | x7);
  assign n786 = ~x3 & (n788 | (~x2 & ~n787));
  assign n787 = x5 ? (x1 ? (~x6 | ~x7) : (x6 | x7)) : ((~x0 | (x7 ? x6 : ~x1)) & (x1 | (~x6 & ~x7)));
  assign n788 = x2 & ((~x1 & (x0 ? (x5 ^ ~x6) : (x5 & ~x6))) | (~x0 & ~x5 & (x1 | x6)));
  assign n789 = (~n792 | ~n793) & (~x3 | n790 | n791);
  assign n790 = x2 ? (~x6 | x7) : (x6 | ~x7);
  assign n791 = x0 ^ ~x5;
  assign n792 = x5 & (x6 | x7);
  assign n793 = ~x3 & x0 & ~x2;
  assign z011 = n795 | ~n799 | ~n803 | (~n640 & ~n798);
  assign n795 = ~n643 & (~n797 | (x3 & ~n796));
  assign n796 = (~x0 | x4 | (x1 ? (x2 | x5) : (~x2 | ~x5))) & (x0 | x1 | ~x2 | ~x4 | ~x5);
  assign n797 = (~x1 | x2 | (x3 & (x0 | x4))) & (~x0 | x1 | ~x2 | ~x3 | ~x4);
  assign n798 = (x0 | ~x3 | (x1 ? (~x2 | ~x4) : (x2 | x4))) & (x1 | x2 | x3 | (~x0 & ~x4));
  assign n799 = ~n801 & (n544 | n800) & (~n601 | ~n802);
  assign n800 = x0 ? (x1 | x6) : (~x1 | ~x6);
  assign n801 = n742 & ((~x1 & ~x6 & (~x3 | ~x4)) | (x1 & x3 & ~x4 & x6));
  assign n802 = x3 & ~x2 & ~x0 & x1;
  assign n803 = (~n804 | n805) & (~n527 | (~n806 & ~n808));
  assign n804 = ~x1 & ~x2;
  assign n805 = (~x0 | ~x3 | x4 | x6 | x7) & (x0 | ((~x6 | ~x7 | x3 | x4) & (x6 | x7 | ~x3 | ~x4)));
  assign n806 = x3 & ~n807 & (x2 ? ~x5 : (x5 & x7));
  assign n807 = x0 ^ ~x4;
  assign n808 = n547 & n809;
  assign n809 = ~x7 & ~x4 & x5;
  assign z012 = ~n821 | n811 | n818;
  assign n811 = x3 & ((n816 & n817) | (~x4 & ~n812));
  assign n812 = (~n560 | ~n813) & (~x7 | n814 | n815);
  assign n813 = ~x7 & ~x5 & ~x6;
  assign n814 = x0 ? (x1 | x5) : (~x1 | ~x5);
  assign n815 = x2 ^ ~x6;
  assign n816 = ~x2 & ~x0 & ~x1;
  assign n817 = x7 & x6 & x4 & ~x5;
  assign n818 = x3 & (x4 ? (n626 & ~n820) : ~n819);
  assign n819 = (~x1 | x5 | (x0 ? (x2 | x7) : (~x2 | ~x7))) & (~x0 | x1 | ~x5 | (~x2 ^ x7));
  assign n820 = x2 ? (x5 ^ ~x7) : (~x5 ^ ~x7);
  assign n821 = ~n822 & ~n824 & n827 & (x3 | n826);
  assign n822 = ~n823 & (x2 ? (x3 ? (x4 & ~x7) : x7) : (x3 ? (x4 & x7) : ~x7));
  assign n823 = x0 ^ ~x1;
  assign n824 = ~x4 & n825 & ((~x2 & ~x7) | (~x1 & x2 & x7));
  assign n825 = ~x0 & x3;
  assign n826 = (x0 | x1 | (x2 ? ~x7 : (~x4 | x7))) & (~x0 | ~x1 | x2 | x7);
  assign n827 = (~n829 | ~n830) & (~n750 | ~n828 | ~n816);
  assign n828 = ~x3 & ~x4;
  assign n829 = ~x3 & ~x2 & ~x0 & ~x1;
  assign n830 = ~x7 & x6 & ~x4 & ~x5;
  assign z013 = n832 | n834 | ~n840 | (~x3 & ~n839);
  assign n832 = ~x1 & ((n704 & n594) | (~x3 & ~n833));
  assign n833 = (x0 | ~x2 | ~x4 | x5 | ~x6) & (x4 | ((~x0 | x2 | (~x5 & ~x6)) & (x0 | ~x2 | x5 | x6)));
  assign n834 = x6 & ((n837 & n838) | (~n835 & ~n836));
  assign n835 = x3 ^ x7;
  assign n836 = (~x2 | x4 | x5 | ~x0 | x1) & (x0 | ((x1 | x2 | ~x4 | x5) & (~x1 | x4 | ~x5)));
  assign n837 = ~x2 & x0 & x1;
  assign n838 = ~x7 & ~x5 & ~x3 & ~x4;
  assign n839 = (~x0 | x1 | x4 | x5 | x6) & (x0 | ((~x1 | x4 | ~x5 | x6) & (x1 | x5 | (~x4 ^ x6))));
  assign n840 = ~n842 & n844 & (~n841 | ~n843);
  assign n841 = x0 & ~x1;
  assign n842 = ~x0 & ((x1 & (x3 ? x4 : (~x4 & ~x5))) | (x5 & ((x3 & x4) | (~x1 & ~x3 & ~x4))));
  assign n843 = x3 & (x4 | x5);
  assign n844 = (~n837 | ~n846) & (~n845 | ~n829);
  assign n845 = x7 & ~x6 & ~x4 & ~x5;
  assign n846 = ~x6 & ~x5 & ~x3 & ~x4;
  assign z014 = ~n862 | ~n855 | n848 | n853;
  assign n848 = ~x2 & ((~n851 & n852) | (~x3 & ~n849));
  assign n849 = (x1 | n850) & (n671 | n791 | ~x1 | ~x6);
  assign n850 = (~x4 | ((~x6 | ~x7 | x0 | x5) & (x6 | x7 | ~x0 | ~x5))) & (x0 | x4 | x5 | (~x6 ^ x7));
  assign n851 = x1 ? (~x5 | (~x4 ^ x7)) : (x5 | (~x4 ^ ~x7));
  assign n852 = x6 & ~x0 & x3;
  assign n853 = ~x2 & ((n704 & n712) | (~x6 & ~n854));
  assign n854 = (~x4 | (x0 ? (x5 | (x1 ^ ~x3)) : (~x1 | ~x5))) & (x0 | x1 | ~x3 | x4 | x5);
  assign n855 = ~n857 & n858 & (x2 | n856 | ~n841);
  assign n856 = x3 ? (x4 | ~x5) : (~x4 | x5);
  assign n857 = ~x0 & (x1 ? (x4 & ~x5) : ((x4 & x5) | (x2 & ~x4 & ~x5)));
  assign n858 = (~n841 | ~n860) & (x6 | ~n859 | n861);
  assign n859 = x2 & x4;
  assign n860 = x5 & x2 & ~x4;
  assign n861 = (x0 | ~x1 | x3 | ~x5) & (~x0 | x1 | x5);
  assign n862 = ~n864 & (~x1 | n863);
  assign n863 = (~x0 | x2 | x3 | x4 | ~x5) & (x0 | ((~x4 | ~x5 | ~x2 | ~x3) & (x4 | x5 | x2 | x3)));
  assign n864 = n865 & ((n866 & n867) | (~n671 & ~n861));
  assign n865 = x2 & x6;
  assign n866 = x3 & ~x0 & x1;
  assign n867 = x7 & ~x4 & x5;
  assign z015 = ~n884 | ~n883 | n879 | n869 | n875;
  assign n869 = ~x2 & (n870 | (n738 & n874));
  assign n870 = x4 & ((~n871 & n872) | (n779 & n873));
  assign n871 = x3 ? (~x6 | x7) : (x6 | ~x7);
  assign n872 = x5 & x0 & ~x1;
  assign n873 = ~x3 & ~x0 & x1;
  assign n874 = x5 & (~x6 | ~x7);
  assign n875 = n878 & (x0 ? (~x1 & ~n877) : (x1 & n876));
  assign n876 = x3 & ~x5;
  assign n877 = x3 ^ x5;
  assign n878 = ~x2 & ~x6;
  assign n879 = (n706 | n881) & (n880 | (~x1 & ~n882));
  assign n880 = ~x3 & ~x2 & x0 & x1;
  assign n881 = x6 & (~x5 ^ ~x7);
  assign n882 = x0 ^ x2;
  assign n883 = (~x0 | x1 | x2 | x5 | ~x6) & (x0 | ~x2 | (x1 ? (x5 | x6) : ~x5));
  assign n884 = ~x6 | ~n543 | (n887 & (~n885 | ~n886));
  assign n885 = x2 & x3;
  assign n886 = x7 & (x4 ^ x5);
  assign n887 = x7 ? (~x5 | (x2 & x3)) : (x5 | (~x2 & ~x3));
  assign z016 = n903 | n901 | n896 | n889 | n892;
  assign n889 = ~n640 & (~n891 | (n691 & ~n890));
  assign n890 = x0 ? (x1 | ~x4) : (x3 | x4);
  assign n891 = (~x0 & (x2 ? ~x1 : (~x3 & ~x4))) | (x1 & x2 & (x0 | (x3 & x4))) | (x0 & ~x2 & (~x1 | x3));
  assign n892 = ~x6 & ((n894 & n895) | (~x0 & ~n893));
  assign n893 = (~x1 | x2 | x3 | x4 | x5) & (~x2 | ((~x3 | (x1 & (~x4 | ~x5))) & (x1 | (~x4 & ~x5))));
  assign n894 = ~x3 & (~x4 | ~x5);
  assign n895 = ~x2 & x0 & ~x1;
  assign n896 = ~x2 & ((~n897 & n898) | (~n899 & n900));
  assign n897 = (~x1 | ~x3 | x4 | x5 | x6) & (x1 | x3 | ~x4 | ~x5 | ~x6);
  assign n898 = x0 & ~x7;
  assign n899 = x1 ? (~x5 | x6) : (x5 | ~x6);
  assign n900 = x7 & ~x4 & ~x0 & ~x3;
  assign n901 = x6 & n902 & n841 & (~x4 | ~x5);
  assign n902 = ~x2 & x3;
  assign n903 = ~n905 & n742 & ~x7 & n904;
  assign n904 = ~x5 & ~x6;
  assign n905 = x1 ? (~x3 | ~x4) : (x3 | x4);
  assign z017 = ~n915 | n912 | n907 | n910;
  assign n907 = ~x0 & (n908 | (n676 & n830));
  assign n908 = x7 & (x1 ? ~n909 : (n596 & n696));
  assign n909 = (~x2 | ~x3 | ~x4 | x5 | x6) & (x2 | x3 | x4 | ~x5 | ~x6);
  assign n910 = ~x1 & (x0 ? n911 : (n596 & n809));
  assign n911 = ~x2 & x3 & x4 & (x5 ^ ~x7);
  assign n912 = ~x7 & (n914 | (~x0 & ~x3 & ~n913));
  assign n913 = x1 ? (x2 | x4) : (~x2 | ~x4);
  assign n914 = ~x4 & x3 & ~x2 & x0 & ~x1;
  assign n915 = ~n916 & ~n919 & n921 & (n917 | ~n918);
  assign n916 = ~x1 & (x0 ? (x2 ? x7 : (~x3 & ~x7)) : (x2 ? (x3 & ~x7) : x7));
  assign n917 = x0 ? (x2 | x3) : (x2 ^ ~x3);
  assign n918 = x1 & x7;
  assign n919 = ~n920 & x7 & n543;
  assign n920 = x2 ? (~x3 | x4) : (x3 | ~x4);
  assign n921 = (~n746 | ~n923) & (~n902 | ~n922 | ~n845);
  assign n922 = x0 & x1;
  assign n923 = ~x7 & x5 & x3 & x4;
  assign z018 = n940 | n937 | ~n930 | n925 | n929;
  assign n925 = n742 & ((n926 & n927) | (~x1 & ~n928));
  assign n926 = ~x6 & x4 & ~x5;
  assign n927 = x1 & x3;
  assign n928 = (x5 | x6 | x3 | x4) & (~x5 | ~x6 | ~x3 | ~x4);
  assign n929 = ~x1 & ((~x3 & x4 & ~x0 & ~x2) | (x0 & x3 & (x2 ^ ~x4)));
  assign n930 = ~n880 & ~n932 & n933 & (~n664 | ~n931);
  assign n931 = ~x7 & x6 & x4 & ~x5;
  assign n932 = ~x4 & x3 & x2 & ~x0 & x1;
  assign n933 = ~n935 & (~n934 | (~n738 & ~n936));
  assign n934 = ~x2 & ~x5;
  assign n935 = ~x0 & (x1 ? (x2 & ~x3) : (~x2 & x3));
  assign n936 = x4 & x3 & x0 & ~x1;
  assign n937 = ~x2 & (n938 | (x5 & ~n682 & n939));
  assign n938 = x0 & ~n897;
  assign n939 = ~x4 & ~x0 & ~x3;
  assign n940 = ~x2 & (n941 | (n543 & n946));
  assign n941 = x0 & ((n943 & n944) | (n942 & n945));
  assign n942 = ~x7 & ~x5 & x6;
  assign n943 = x7 & x5 & ~x6;
  assign n944 = x4 & ~x1 & ~x3;
  assign n945 = ~x4 & x1 & x3;
  assign n946 = x5 & x6 & (x3 ? (x4 & x7) : (~x4 & ~x7));
  assign z019 = ~n956 | (~x0 & (n948 | n952 | ~n953));
  assign n948 = x1 & ((n949 & n951) | (x4 & ~n950));
  assign n949 = ~x4 & ~x2 & x3;
  assign n950 = (x2 | ~x3 | ~x5 | ~x6 | x7) & (~x2 | ((~x3 | x5 | ~x6 | x7) & (x3 | ~x5 | x6 | ~x7)));
  assign n951 = x7 & ~x5 & ~x6;
  assign n952 = n558 & n845;
  assign n953 = x2 ? n954 : n955;
  assign n954 = (x4 | (~x3 & (x1 | x5 | x6))) & (~x1 | x3 | ~x4 | ~x5 | ~x6) & (~x3 | ((x5 | x6) & (x1 | (x5 & x6))));
  assign n955 = (x1 & (~x3 | (x4 & x5 & x6))) | (~x3 & (x4 | (x5 & x6))) | (~x4 & ~x5 & (~x6 | (~x1 & x3)));
  assign n956 = ~x0 | (~n958 & (x2 | (n957 & n961)));
  assign n957 = x3 ? ((x4 | x5 | x6) & (x1 | (x4 & x5))) : ((~x4 | ~x6) & (~x1 | (~x4 & (~x5 | ~x6))));
  assign n958 = n570 & (n774 | n959 | n960);
  assign n959 = x5 & ~x3 & x4;
  assign n960 = x6 & ~x5 & ~x3 & x4;
  assign n961 = (~x1 | ~x3 | x4 | ~n942) & (x1 | x3 | ~x4 | ~n962);
  assign n962 = ~x6 & (~x5 ^ ~x7);
  assign z020 = n964 | ~n966 | n983 | (~x0 & ~n974);
  assign n964 = ~x6 & (x0 ? ~n965 : (n731 & n570));
  assign n965 = (x1 | ~x2 | x3 | ~x4 | x5) & (~x1 | x2 | x4 | (~x3 ^ x5));
  assign n966 = n970 & (n968 | n969) & (x1 | n967);
  assign n967 = (~x5 | (x0 ? (x4 | (~x2 & x3)) : (~x4 | (x2 ^ ~x3)))) & (~x3 | x5 | (x0 ? (x2 | ~x4) : (~x2 ^ ~x4)));
  assign n968 = x2 ^ ~x5;
  assign n969 = (~x3 | ((x4 | ~x6 | ~x0 | x1) & (x0 | ~x1 | ~x4 | x6))) & (x0 | x1 | x3 | (~x4 ^ ~x6));
  assign n970 = (~x1 | n972) & (~n971 | n973);
  assign n971 = ~x3 & x6;
  assign n972 = (~x0 | x2 | x3 | x4 | x5) & (x0 | (x2 ? (x3 ? (x4 | ~x5) : (~x4 | x5)) : (~x4 | (~x3 ^ x5))));
  assign n973 = (x4 | x5 | x1 | x2) & (~x1 | ((x0 | (x2 ? (x4 | ~x5) : (~x4 | x5))) & (~x4 | ~x5 | ~x0 | x2)));
  assign n974 = x4 ? (n977 & (n975 | n976)) : n980;
  assign n975 = x3 ? (x5 | ~x6) : (~x5 | x6);
  assign n976 = x1 ? (~x2 | x7) : (x2 | ~x7);
  assign n977 = (~n676 | ~n951) & (~n978 | ~n979);
  assign n978 = ~x7 & x5 & x6;
  assign n979 = x3 & x1 & ~x2;
  assign n980 = x7 ? n982 : (n981 | ~n632);
  assign n981 = x3 ? (x5 | x6) : (~x5 | ~x6);
  assign n982 = (x1 | ((~x5 | ~x6 | ~x2 | ~x3) & (x5 | x6 | x2 | x3))) & (~x1 | x2 | x3 | ~x5 | x6);
  assign n983 = x0 & (n984 | (x7 & n570 & ~n987));
  assign n984 = ~x2 & ((x1 & ~n985) | (n527 & ~n986));
  assign n985 = (x3 | ~x4 | ~x5 | x6 | ~x7) & (~x3 | x4 | x5 | ~x6 | x7);
  assign n986 = (~x5 | ~x7 | ~x3 | x4) & (x3 | ~x4 | (~x5 ^ ~x7));
  assign n987 = (~x3 | (x4 ? (~x5 | ~x6) : (x5 | x6))) & (x3 | x4 | x5 | ~x6);
  assign z021 = n997 | ~n1000 | ~n1013 | (~x1 & ~n989);
  assign n989 = ~n994 & (x2 | (~n991 & (~n653 | n990)));
  assign n990 = (x4 | x5 | ~x6 | ~x7) & (x6 | x7 | ~x4 | ~x5);
  assign n991 = n536 & (n993 | (x4 & n992));
  assign n992 = x7 & (x5 ^ ~x6);
  assign n993 = ~x7 & ~x6 & ~x4 & x5;
  assign n994 = n995 & ~n996;
  assign n995 = x0 & x2;
  assign n996 = (~x3 | x4 | x5 | x6 | x7) & (x3 | ((x4 | x5 | ~x6 | x7) & (x6 | ~x7 | ~x4 | ~x5)));
  assign n997 = ~x2 & (x4 ? ~n999 : ~n998);
  assign n998 = ((x0 ? (x3 | x6) : (~x3 | ~x6)) | (~x1 ^ ~x5)) & (~x0 | ((~x5 | ~x6 | x1 | x3) & (x5 | x6 | ~x1 | ~x3))) & (x0 | x3 | (x1 ? (x5 | ~x6) : (~x5 | x6)));
  assign n999 = (~x0 | x1 | x3 | ~x5 | x6) & (x0 | (((~x3 ^ ~x5) | (x1 ^ ~x6)) & (~x1 | x3 | ~x5 | ~x6)));
  assign n1000 = ~n1004 & ~n1007 & (~x2 | (n1001 & n1003));
  assign n1001 = (~n577 | ~n712) & (x0 | n1002);
  assign n1002 = (x1 | ~x3 | ~x4 | x5 | ~x6) & (~x1 | x3 | x4 | ~x5 | x6) & ((~x4 ^ ~x5) | (x1 ? (~x3 | ~x6) : (x3 | x6)));
  assign n1003 = (~x0 | x1 | x3 | x5 | x6) & (((x1 | ~x5) & (x0 | ~x1 | x5)) | (~x3 ^ x6));
  assign n1004 = n934 & ((n626 & n1005) | (x0 & n1006));
  assign n1005 = x3 & ~x6;
  assign n1006 = x6 & (x1 ^ x3);
  assign n1007 = ~n1008 & ((~n1011 & n1012) | (~n1009 & ~n1010));
  assign n1008 = x5 ^ ~x7;
  assign n1009 = (x3 | x6 | ~x1 | x2) & (~x3 | ~x6 | x1 | ~x2);
  assign n1010 = x0 ^ x4;
  assign n1011 = x2 ? (x3 | x6) : (~x3 | ~x6);
  assign n1012 = x4 & ~x0 & x1;
  assign n1013 = (n1014 | n1015) & (n1016 | ~n1017);
  assign n1014 = x4 ? (x5 | x7) : (~x5 | ~x7);
  assign n1015 = (~x0 | x1 | x2 | x3 | x6) & (x0 | ((~x3 | ~x6 | ~x1 | ~x2) & (x1 | (x2 ? (x3 | x6) : (~x3 | ~x6)))));
  assign n1016 = (~x0 | ~x3 | x5 | ~x6 | x7) & (x0 | ((x3 | ~x5 | ~x6 | ~x7) & (~x3 | x6 | (~x5 ^ ~x7))));
  assign n1017 = ~x4 & x1 & ~x2;
  assign z022 = n1031 | ~n1037 | (x0 ? ~n1019 : ~n1023);
  assign n1019 = x1 ? (~n902 | ~n830) : n1020;
  assign n1020 = x4 ? n1022 : (~n596 | (~n943 & ~n1021));
  assign n1021 = ~x5 & (~x6 ^ ~x7);
  assign n1022 = (x2 | x3 | ~x5 | x6 | ~x7) & (~x3 | ((~x5 | ~x6 | x7) & (~x2 | (~x6 ^ x7))));
  assign n1023 = ~n1028 & (x4 | (n1025 & (~x2 | n1024)));
  assign n1024 = (~x1 | x3 | x5 | x6 | ~x7) & (~x3 | ~x5 | ((x6 | ~x7) & (x1 | ~x6 | x7)));
  assign n1025 = (~n978 | ~n669) & (n1026 | n1027);
  assign n1026 = x3 ^ x6;
  assign n1027 = x1 ? (~x5 | x7) : (x5 | (~x2 ^ x7));
  assign n1028 = n1029 & ~n1030;
  assign n1029 = x3 & x4;
  assign n1030 = x6 ? (x7 | ((x2 | x5) & (~x1 | (x2 & x5)))) : (~x7 | ((~x1 | ~x2 | x5) & (~x5 | (x1 & x2))));
  assign n1031 = ~n640 & (n1033 | ~n1034 | (~x1 & ~n1032));
  assign n1032 = (x0 | ~x2 | (x3 ? (~x4 | ~x5) : (~x4 ^ x5))) & (~x0 | x2 | ~x4 | x5);
  assign n1033 = ~x3 & ((~x0 & x1 & x2 & x4) | (~x2 & (x0 ? (x1 ^ ~x4) : (~x1 & x4))));
  assign n1034 = ~n914 & (~n1017 | n1035) & (n647 | n1036);
  assign n1035 = x0 ? (x3 | ~x5) : (~x3 ^ ~x5);
  assign n1036 = x0 ? (x1 | ~x2) : (~x1 | x2);
  assign n1037 = ~n1043 & (n1041 | n1042) & (~x2 | n1038);
  assign n1038 = (x1 | n1039) & (x0 | ~x1 | ~x3 | n1040);
  assign n1039 = x0 ? ((~x3 | x4 | ~x5 | ~x6) & (x3 | ~x4 | x5 | x6)) : (~x4 | (x3 ? (x5 | x6) : (~x5 | ~x6)));
  assign n1040 = x4 ? (~x5 | x6) : (x5 | ~x6);
  assign n1041 = (x2 | (x0 ? (x4 ? (~x6 | x7) : (x6 | ~x7)) : (x4 ? (x6 | ~x7) : (~x6 | x7)))) & (x0 | ~x2 | x4 | x6 | ~x7);
  assign n1042 = x1 ? (x3 | ~x5) : x5;
  assign n1043 = ~x6 & n1044 & (n1045 | (n681 & n922));
  assign n1044 = ~x2 & ~x3;
  assign n1045 = ~x0 & (x1 ? (x4 & ~x5) : (~x4 & x5));
  assign z023 = n1067 | n1064 | n1058 | n1047 | n1055;
  assign n1047 = ~x2 & (~n1052 | (~x0 & (n1048 | n1050)));
  assign n1048 = x6 & ~n1049;
  assign n1049 = (x1 | ~x3 | x4 | x5 | ~x7) & (x7 | ((~x1 | (x3 ? (~x4 | ~x5) : (x4 | x5))) & (x1 | x3 | ~x4 | ~x5)));
  assign n1050 = x7 & n1051 & (x1 ? x4 : (~x4 & x5));
  assign n1051 = ~x3 & ~x6;
  assign n1052 = ~n1054 & (~n661 | ~n662) & (x4 | n1053);
  assign n1053 = (x0 | ~x1 | ~x5 | x6 | x7) & (~x0 | ((~x1 | x5 | x6 | ~x7) & (x1 | ~x6 | x7)));
  assign n1054 = x7 & ~x5 & x4 & x0 & ~x1;
  assign n1055 = ~n1008 & (x0 ? ~n1057 : ~n1056);
  assign n1056 = x2 ? ((x1 | (x3 ? (~x4 | ~x6) : x4)) & (x4 | ~x6 | ~x1 | ~x3)) : (~x4 | (x1 ? (~x3 ^ x6) : (x3 | x6)));
  assign n1057 = (~x1 | x2 | x3 | x4 | ~x6) & (x1 | (x2 ? (x3 | ~x4) : (x4 | x6)));
  assign n1058 = ~n765 & (~n1060 | (~x1 & ~n1059));
  assign n1059 = x0 ? ((~x2 | x3 | x4 | ~x6) & (x2 | ~x4 | x6)) : (x2 | ~x6 | (~x3 ^ ~x4));
  assign n1060 = ~n1061 & (~n873 | n1063) & (~x0 | n1062);
  assign n1061 = ~x0 & ((~x1 & x2 & ~x3 & x4) | (x1 & x3 & (x2 ^ ~x4)));
  assign n1062 = (x1 | ~x2 | ~x3 | x4) & (x3 | ~x4 | ~x1 | x2);
  assign n1063 = (x4 | x6) & (~x2 | ~x4 | ~x6);
  assign n1064 = ~n671 & (x0 ? ~n1065 : ~n1066);
  assign n1065 = (x1 | ~x2 | ~x3 | x5 | ~x6) & (~x1 | x2 | x3 | ~x5 | x6);
  assign n1066 = (x1 | x2 | (x3 ? x6 : (x5 | ~x6))) & (~x1 | ~x2 | x3 | ~x5 | ~x6);
  assign n1067 = x2 & (n1075 | (~x1 & (n1068 | ~n1069)));
  assign n1068 = ~x0 & x3 & (x4 ? (~x6 & x7) : (x6 & ~x7));
  assign n1069 = ~n1073 & (n1071 | ~n1072) & (~n1070 | ~n1074);
  assign n1070 = x7 & ~x5 & x6;
  assign n1071 = x0 ? ~x4 : (x4 | x6);
  assign n1072 = ~x7 & x3 & x5;
  assign n1073 = ~x7 & ~x6 & ~x4 & x0 & ~x3;
  assign n1074 = x4 & ~x0 & ~x3;
  assign n1075 = n543 & ~n1076;
  assign n1076 = (~x3 | x4 | x5 | x6 | ~x7) & (x3 | ((~x6 | ~x7 | x4 | x5) & (~x4 | x6 | x7)));
  assign z024 = n1092 | ~n1096 | (x3 ? ~n1078 : ~n1086);
  assign n1078 = ~n1079 & ~n1083;
  assign n1079 = ~x1 & ((x2 & ~n1081) | (n1080 & ~n1082));
  assign n1080 = ~x2 & ~x7;
  assign n1081 = (x5 | ((x7 | (x0 ? (~x4 ^ x6) : (x4 | x6))) & (x0 | ~x4 | ~x6 | ~x7))) & (~x0 | ~x4 | ~x5 | x6 | ~x7);
  assign n1082 = (x0 | x4 | ~x5 | ~x6) & (~x0 | ~x4 | (~x5 ^ ~x6));
  assign n1083 = x1 & (x0 ? (n942 & n1084) : ~n1085);
  assign n1084 = ~x2 & ~x4;
  assign n1085 = x4 ? ((~x2 | ~x7 | (~x5 ^ ~x6)) & (x2 | x5 | ~x6 | x7)) : (x6 | ((~x5 | x7) & (x2 | x5 | ~x7)));
  assign n1086 = x2 ? n1089 : (x1 ? n1087 : n1088);
  assign n1087 = x0 ? ((~x6 | ~x7 | x4 | x5) & (x6 | x7 | ~x4 | ~x5)) : ((~x4 | x5 | ~x6 | ~x7) & (x4 | (x5 ? (~x6 ^ ~x7) : (x6 | ~x7))));
  assign n1088 = (~x4 | ((~x0 | ((x6 | x7) & (~x5 | ~x6 | ~x7))) & (x6 | ~x7 | x0 | ~x5))) & (x0 | x4 | (x5 ? (~x6 | ~x7) : (~x6 ^ x7)));
  assign n1089 = (~x6 | x7 | ~n566 | n1090) & (~x7 | n1091);
  assign n1090 = x1 ^ x5;
  assign n1091 = (x0 | ~x1 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (x1 | ((~x5 | ~x6 | x0 | x4) & (x5 | (x0 ? (~x4 ^ x6) : (x4 | x6)))));
  assign n1092 = x3 & ((n551 & ~n1094) | (n1093 & ~n1095));
  assign n1093 = x1 & ~x5;
  assign n1094 = (x0 | (x4 ? x6 : ~x2)) & (~x4 | ((x2 | x6) & (~x0 | ~x2 | ~x6)));
  assign n1095 = (x4 | x6 | ~x0 | x2) & (x0 | ~x6 | (~x2 & x4));
  assign n1096 = ~n1099 & (n1097 | n1098) & (~n653 | n1102);
  assign n1097 = x5 ^ x6;
  assign n1098 = (x0 | ~x1 | (x2 ? (x3 | x4) : (~x3 | ~x4))) & (x1 | (x0 ? (x4 | (x2 & ~x3)) : (x3 | ~x4)));
  assign n1099 = ~n1100 & (n1101 | (n902 & n626));
  assign n1100 = x4 ? (x5 | ~x6) : (~x5 | x6);
  assign n1101 = x0 & ~x3 & (~x1 ^ ~x2);
  assign n1102 = (x1 | ~x2 | x4 | x5 | ~x6) & (~x1 | ((~x4 | ~x5 | x6) & (x5 | ~x6 | x2 | x4)));
  assign z025 = ~n1114 | (x2 ? (n1110 | ~n1112) : ~n1104);
  assign n1104 = x5 ? n1107 : (x0 ? n1105 : n1106);
  assign n1105 = x1 ? ((~x3 | x4 | ~x6 | x7) & (x3 | ~x4 | x6 | ~x7)) : ((x4 | x6 | ~x7) & (~x3 | ~x4 | ~x6 | x7));
  assign n1106 = (~x4 | x6 | ((x3 | ~x7) & (x1 | (x3 & ~x7)))) & (x1 | ~x3 | x4 | ~x6 | ~x7);
  assign n1107 = (x7 | n1108) & (~n527 | ~n1109);
  assign n1108 = (x0 | ((x4 | ~x6) & (~x1 | x3 | ~x4 | x6))) & (~x4 | ~x6 | ~x0 | x1);
  assign n1109 = x7 & (x0 ? ~x4 : (x3 & x4));
  assign n1110 = ~x0 & (x1 ? (n774 & n813) : ~n1111);
  assign n1111 = (~x4 | x5 | x6 | ~x7) & (x4 | ~x6 | (x3 ? ~x5 : x7));
  assign n1112 = (n1113 | n823) & (~n661 | ~n662);
  assign n1113 = (x4 | x5 | x6 | ~x7) & (~x4 | ~x5 | ~x6 | x7);
  assign n1114 = ~n1115 & (n640 | (~n1118 & ~n1120 & n1123));
  assign n1115 = ~n1116 & ~n1117;
  assign n1116 = x5 ? (x6 | ~x7) : (~x6 | x7);
  assign n1117 = (~x1 | ((x3 | x4 | ~x0 | x2) & (x0 | ~x4))) & (x0 | ~x2 | ~x4) & (x1 | (x0 ? (x2 ? x4 : (x3 | ~x4)) : (x2 | x4)));
  assign n1118 = ~n714 & (n560 | (x2 & ~n1119));
  assign n1119 = x0 ? (x1 | x3) : (~x1 | ~x3);
  assign n1120 = n626 & (~n1122 | (n1121 & n596));
  assign n1121 = x4 & x5;
  assign n1122 = x2 ? (x4 | x5) : (~x4 | ~x5);
  assign n1123 = x0 ? (~x4 | (x1 ? (x2 | x3) : (~x2 | ~x3))) : (~x1 | x4 | (x2 & x3));
  assign z026 = n1136 | ~n1142 | (x0 ? ~n1125 : ~n1129);
  assign n1125 = ~n1126 & (~n845 | ~n979) & (n765 | n1128);
  assign n1126 = ~x1 & (x2 ? (n774 & n813) : ~n1127);
  assign n1127 = (x4 | ~x5 | x6 | ~x7) & (~x4 | x5 | (x3 ? (~x6 | ~x7) : (x6 | x7)));
  assign n1128 = (x2 | ((~x4 | x6 | x1 | ~x3) & (x4 | ~x6 | ~x1 | x3))) & (x1 | ~x2 | (x6 ? (~x3 & ~x4) : x3));
  assign n1129 = ~n1130 & ~n1132 & (x1 | x7 | n909);
  assign n1130 = ~n765 & ~n1131;
  assign n1131 = (x2 & (x1 | (~x3 & x6))) | (x3 & x4 & ~x6) | (~x2 & (~x1 | (~x4 & ~x6)));
  assign n1132 = ~n1134 & ((n804 & n684) | (n1133 & n1135));
  assign n1133 = x1 & x2;
  assign n1134 = x4 ^ x5;
  assign n1135 = ~x7 & ~x3 & x6;
  assign n1136 = ~n1008 & (n1137 | ~n1140 | (~n1138 & n1139));
  assign n1137 = ~x2 & ((~x3 & (x0 ? (~x1 ^ ~x6) : (~x1 & ~x6))) | (~x0 & ~x1 & x3 & x6));
  assign n1138 = x1 ? (~x3 | x6) : (x3 | ~x6);
  assign n1139 = ~x0 & (~x2 ^ ~x4);
  assign n1140 = (x0 | ~x1 | ~x2 | n1026) & (x2 | ~n1141 | ~x0 | x1);
  assign n1141 = x6 & x3 & ~x4;
  assign n1142 = x0 ? n1144 : (~n1149 & (n1143 | n1148));
  assign n1143 = x2 ? (x3 | ~x6) : (~x3 | x6);
  assign n1144 = x5 ? n1147 : (~n1145 | (~n1146 & ~n878));
  assign n1145 = ~x1 & ~x4;
  assign n1146 = x6 & x2 & ~x3;
  assign n1147 = (x1 | ~x2 | ~x3 | x6) & (~x1 | x2 | x3 | ~x4 | ~x6);
  assign n1148 = x1 ? (x4 | ~x5) : (~x4 | x5);
  assign n1149 = ~x6 & ((n731 & n570) | (x1 & ~n1150));
  assign n1150 = (x2 | x3 | x4 | ~x5) & (~x2 | ~x3 | ~x4 | x5);
  assign z027 = ~n1168 | n1162 | n1159 | n1152 | n1155;
  assign n1152 = ~n643 & (x0 ? ~n1153 : ~n1154);
  assign n1153 = (x2 | ((~x4 | ~x5 | x1 | ~x3) & (~x1 | (x3 ? (x4 | x5) : ~x4)))) & (x3 | x4 | x1 | ~x2);
  assign n1154 = (x3 | x4 | x1 | x2) & (~x2 | ((x1 | (x3 ? (x4 | x5) : ~x4)) & (x3 | ((~x4 | x5) & (~x1 | x4 | ~x5)))));
  assign n1155 = ~x0 & ((x4 & ~n1157) | (n1156 & ~n1158));
  assign n1156 = x2 & ~x4;
  assign n1157 = (x1 | x2 | ~x3 | ~x5 | x6) & (~x6 | ((x1 | ~x2 | ~x3 | x5) & (~x1 | x3 | (~x2 ^ ~x5))));
  assign n1158 = (x5 | x6 | ~x1 | x3) & (~x5 | ~x6 | x1 | ~x3);
  assign n1159 = ~n640 & ((n841 & ~n1161) | (~x0 & ~n1160));
  assign n1160 = (~x1 | (x2 ? (~x3 | ~x4) : x4)) & (~x3 | (x2 ? (~x4 | ~x5) : ((x4 | ~x5) & (x1 | ~x4 | x5))));
  assign n1161 = (x2 | x3 | ~x4 | ~x5) & (~x3 | (x2 ? (~x4 ^ x5) : (x4 | x5)));
  assign n1162 = ~x2 & (n1163 | (~x1 & n1166));
  assign n1163 = ~n1165 & ~x3 & ~n1164;
  assign n1164 = x1 ^ x4;
  assign n1165 = (x6 | x7 | ~x0 | x5) & (~x6 | ~x7 | x0 | ~x5);
  assign n1166 = x3 & ((n1070 & n1167) | (n525 & n658));
  assign n1167 = ~x0 & ~x4;
  assign n1168 = n1170 & (~n570 | ~n1166) & (x3 | n1169);
  assign n1169 = x0 ? ((x1 | ~x2 | ~x4 | ~x6) & (~x1 | x2 | x4 | x6)) : (x1 | (x2 ? (x4 | x6) : (~x4 | ~x6)));
  assign n1170 = (x0 | ~x1 | ~x3 | n1171) & (~x0 | x1 | n1172);
  assign n1171 = x2 ? (x4 | ~x6) : (~x4 | x6);
  assign n1172 = (x2 | x6 | (~x4 ^ x5)) & (~x2 | ~x3 | x4 | x5 | ~x6);
  assign z028 = n1180 | ~n1187 | (x1 ? ~n1174 : ~n1177);
  assign n1174 = (x2 | n1175) & (x0 | ~x2 | x3 | n1176);
  assign n1175 = (~x3 | ((x0 | ~x4 | ~x7) & (x4 | x5 | x7))) & (~x0 | x3 | x4 | x5 | ~x7) & (x0 | (x4 ? (x5 | ~x7) : x7));
  assign n1176 = x4 ? (~x5 ^ ~x7) : (~x5 | x7);
  assign n1177 = x4 ? n1178 : n1179;
  assign n1178 = (~x7 | ((~x0 | (x2 ? x3 : x5)) & (x2 | x3 | x5) & (x0 | (x2 ? (~x3 | x5) : ~x5)))) & (x0 | x7 | (x2 ? (x3 | ~x5) : (~x3 | x5)));
  assign n1179 = (~x0 | ((x2 | (~x5 ^ ~x7)) & (x7 | (x5 ? ~x2 : x3)))) & (x0 | x2 | ~x5 | x7);
  assign n1180 = ~x3 & (~n1183 | (x6 & n1181 & ~n1182));
  assign n1181 = ~x0 & ~x2;
  assign n1182 = (~x1 | ~x4 | ~x5 | x7) & (x1 | x4 | (~x5 ^ ~x7));
  assign n1183 = (n1185 | n1186) & (n524 | n1184);
  assign n1184 = (x0 | ~x1 | ~x2 | x6) & (x2 | ~x6 | ~x0 | x1);
  assign n1185 = x1 ? (x2 | ~x6) : (~x2 | x6);
  assign n1186 = (x0 | x4 | ~x5 | ~x7) & (x5 | x7 | ~x0 | ~x4);
  assign n1187 = (n671 | n1189) & (n573 | ~n1188 | n1190);
  assign n1188 = ~x1 & x3;
  assign n1189 = x0 ? ((x1 | ~x2 | ~x3 | x5) & (~x1 | x2 | x3 | ~x5)) : (~x2 | ((~x3 | (~x1 & ~x5)) & (x1 | x3 | x5)));
  assign n1190 = x2 ? (~x6 ^ ~x7) : (x6 ^ ~x7);
  assign z029 = n1193 | ~n1196 | ~n1204 | (~x0 & ~n1192);
  assign n1192 = x1 ? ((~x3 | ~x4 | x5) & (~x2 | x3 | x4 | ~x5)) : (~x4 | (~x3 ^ ~x5));
  assign n1193 = n564 & (n1195 | (~x1 & (n691 | n1194)));
  assign n1194 = x2 & (x3 ^ ~x5);
  assign n1195 = ~x5 & ~x3 & x1 & ~x2;
  assign n1196 = ~n1197 & n1201 & (~n653 | ~n681 | ~n1200);
  assign n1197 = ~n1198 & ~n1199;
  assign n1198 = x5 ^ ~x6;
  assign n1199 = (x0 | x1 | ~x3 | x4) & (~x0 | x3 | ~x4 | (x1 ^ ~x2));
  assign n1200 = ~x6 & (x1 ^ x2);
  assign n1201 = (~n559 | ~n712) & (~n543 | (~n1202 & ~n1203));
  assign n1202 = x6 & x5 & ~x3 & x4;
  assign n1203 = ~x6 & ~x5 & x3 & ~x4;
  assign n1204 = (n1205 | (~n1206 & ~n1208)) & (x2 | n1210);
  assign n1205 = x3 ^ ~x7;
  assign n1206 = ~x0 & (n1207 | (n704 & n1133));
  assign n1207 = x5 & (x1 ? (x4 & ~x6) : (~x4 & x6));
  assign n1208 = n926 & n1209;
  assign n1209 = x2 & x0 & ~x1;
  assign n1210 = (x7 | n1211 | ~x3 | x5) & (x3 | ~x7 | (x5 ? n1211 : n1212));
  assign n1211 = (~x0 | x1 | ~x4 | x6) & (x0 | ~x1 | x4 | ~x6);
  assign n1212 = (x4 | x6 | x0 | x1) & (~x0 | (x1 ? (~x4 | x6) : (x4 | ~x6)));
  assign z030 = n1227 | n1225 | n1222 | n1214 | n1217;
  assign n1214 = x6 & ((n733 & n1216) | (~n671 & ~n1215));
  assign n1215 = (~x0 | x1 | x2 | x3 | x5) & (x0 | (x1 ? (x5 | (~x2 & ~x3)) : ~x5));
  assign n1216 = ~x7 & ~x5 & ~x3 & x4;
  assign n1217 = ~x6 & ((~n1218 & ~n1219) | (~x2 & ~n1220));
  assign n1218 = x4 ^ x7;
  assign n1219 = (~x0 | ~x1 | x2 | x3 | x5) & ((~x2 & ~x3) | (x0 ? (x1 | x5) : (~x1 | ~x5)));
  assign n1220 = (~n717 | ~n699) & (x7 | ~n564 | n1221);
  assign n1221 = x1 ? (~x3 | x5) : (x3 | ~x5);
  assign n1222 = x4 & ((~n1097 & ~n1223) | (~x0 & ~n1224));
  assign n1223 = (x2 | x3 | ~x0 | x1) & (x0 | ~x1 | (~x2 & ~x3));
  assign n1224 = (~x1 | x2 | x3 | ~x5 | ~x6) & (x1 | x6 | (~x5 & (x2 | x3)));
  assign n1225 = ~n1226 & (x0 ? (x4 ? x6 : (x5 & ~x6)) : (~x5 & (x4 ^ x6)));
  assign n1226 = x1 ^ (~x2 & ~x3);
  assign n1227 = n816 & n1228;
  assign n1228 = x6 & ~x5 & ~x3 & ~x4;
  assign z031 = ~n1236 | (~x2 & (n1230 | n1233 | ~n1235));
  assign n1230 = ~x3 & (x5 ? n1231 : (n543 & ~n1232));
  assign n1231 = (x4 ^ ~x6) & (x0 ? (~x1 & x7) : (x1 & ~x7));
  assign n1232 = x4 ? (~x6 ^ ~x7) : (~x6 | x7);
  assign n1233 = n845 & n1234;
  assign n1234 = x3 & x0 & x1;
  assign n1235 = (x6 | ~x7 | x0 | ~x5) & (x1 | ((~x6 | x7 | (x0 ^ x5)) & (x0 | ~x5 | (x6 & ~x7))));
  assign n1236 = x2 ? n1237 : (n1239 & (n640 | n1238));
  assign n1237 = (x1 | ((~x0 | (x5 ? x7 : (x6 | ~x7))) & (~x5 | (~x6 ^ ~x7)) & (x0 | x5 | ~x6 | x7))) & (x0 | ((~x5 | ((x6 | ~x7) & (~x1 | ~x6 | x7))) & (~x1 | x5 | (~x6 ^ ~x7))));
  assign n1238 = (~x1 | (x0 ? (x3 | ~x5) : (~x3 | x5))) & (~x0 | x1 | (~x3 ^ ~x5));
  assign n1239 = (~x3 | (x0 ? (x1 | ~n951) : (~x1 | ~n978))) & (~x0 | ~x1 | x3 | (~n978 & ~n951));
  assign z032 = ~n1245 | (~x2 & (n1242 | (n661 & n1241)));
  assign n1241 = ~x7 & x6 & x4 & x5;
  assign n1242 = ~x4 & ((n1093 & ~n1243) | (n658 & n1244));
  assign n1243 = (x0 | x3 | ~x6 | ~x7) & (~x0 | ~x3 | (~x6 ^ x7));
  assign n1244 = ~x3 & ~x0 & ~x1;
  assign n1245 = n1247 & (~x4 | x6 | n1246 | ~n1250);
  assign n1246 = x1 ^ x7;
  assign n1247 = n1249 & (x2 | n1248);
  assign n1248 = (x6 | (~x1 ^ ~x7) | (x0 ^ ~x3)) & (~x0 | ~x6 | x7 | (x1 ^ ~x3));
  assign n1249 = (x1 | (x0 ? ((x6 | ~x7) & (~x2 | ~x6 | x7)) : (~x6 | ~x7))) & (x0 | x6 | ((~x2 | x7) & (~x1 | (~x2 & x7))));
  assign n1250 = ~x3 & ~x0 & ~x2;
  assign z033 = n1252 | n1254 | ~n1256 | (n608 & ~n1255);
  assign n1252 = ~x2 & (x0 ? n1253 : (n689 & n809));
  assign n1253 = ~x5 & ((x1 & x3 & ~x4 & ~x7) | (~x1 & ~x3 & x4 & x7));
  assign n1254 = n1044 & ((~x4 & x7 & x0 & ~x1) | (~x0 & (x1 ? (x4 ^ ~x7) : (x4 & ~x7))));
  assign n1255 = (x0 | x4 | (x1 ? (~x5 | ~x7) : (x5 | x7))) & (~x0 | x1 | ~x4 | ~x5 | x7);
  assign n1256 = (~x0 | ~x1 | x2 | x3 | x7) & ((~x2 & ~x3) | ((x1 | x7) & (x0 | ~x1 | ~x7)));
  assign z035 = ~x2 & (n1258 | ~n1259 | ~n1261);
  assign n1258 = ~x0 & ~x4 & (x1 ? (x3 & ~x5) : (~x3 & x5));
  assign n1259 = n1260 & (~n845 | ~n1244) & (~n559 | ~n661);
  assign n1260 = x0 ? (x1 | ~x3 | (x4 & x5)) : (x3 | ~x4);
  assign n1261 = (~x5 | n1205 | n1211) & (~n1167 | n1262);
  assign n1262 = (x1 | x3 | x5 | ~x6) & (~x1 | ~x3 | ~x5 | x6);
  assign z036 = ~n1267 | ~n1264 | n1266;
  assign n1264 = ~n935 & ~n1265 & (~n526 | ~n902 | n1211);
  assign n1265 = ~x0 & ((x1 & ~x2 & x3 & x4) | (~x1 & x2 & ~x3 & ~x4));
  assign n1266 = x3 & ((n696 & n746) | (n559 & n560));
  assign n1267 = ~n1270 & ~n1271 & (~n1268 | ~n1269);
  assign n1268 = ~x5 & ~x3 & x4;
  assign n1269 = x2 & ~x0 & ~x1;
  assign n1270 = ~x3 & x2 & x0 & ~x1;
  assign n1271 = ~x4 & x3 & x2 & x0 & ~x1;
  assign z037 = n1273 | n1277 | ~n1279 | (~x0 & ~n1276);
  assign n1273 = ~x1 & (x4 ? ~n1274 : (n1021 & n1250));
  assign n1274 = (~n743 | ~n943) & (x7 | n1275);
  assign n1275 = (x0 | ~x2 | ~x3 | x5 | x6) & (~x0 | x3 | ~x6 | (~x2 ^ x5));
  assign n1276 = (x1 | x2 | ~x3 | ~x4 | x5) & (~x2 | ((~x4 | ~x5 | x1 | x3) & (~x1 | x4 | (~x3 ^ ~x5))));
  assign n1277 = x3 & (x0 ? (n559 & n804) : ~n1278);
  assign n1278 = (x1 | x2 | ~x4 | ~x5 | x6) & (~x1 | ~x2 | x4 | x5 | ~x6);
  assign n1279 = ~n1280 & ~n1281 & n1286 & (n1284 | ~n1285);
  assign n1280 = ~x1 & (x0 ? (x2 & (x3 ^ ~x4)) : (x3 & ~x4));
  assign n1281 = n1283 & ((n530 & n774) | (~x3 & ~n1282));
  assign n1282 = (x6 | x7 | ~x4 | x5) & (~x6 | ~x7 | x4 | ~x5);
  assign n1283 = ~x2 & ~x0 & x1;
  assign n1284 = (x1 | ~x2 | ~x4 | x5) & (x4 | ~x5 | ~x1 | x2);
  assign n1285 = ~x6 & x0 & ~x3;
  assign n1286 = (~n1287 | ~n837) & (x0 | ~n1288);
  assign n1287 = ~x5 & ~x3 & ~x4;
  assign n1288 = x4 & x1 & x3;
  assign z038 = n1299 | ~n1304 | (x4 & (~n1290 | ~n1297));
  assign n1290 = x2 ? (~n1292 & (~n1291 | ~n1294)) : n1295;
  assign n1291 = ~x5 & ~x0 & x1;
  assign n1292 = ~x1 & ((n825 & n951) | (x0 & n1293));
  assign n1293 = x6 & (x3 ? (x5 & ~x7) : (~x5 & x7));
  assign n1294 = ~x7 & (x3 ^ x6);
  assign n1295 = (~n712 | ~n943) & (x3 | n1296);
  assign n1296 = (x0 | ~x1 | x5 | x6 | ~x7) & (~x0 | ~x5 | (x1 ? (x6 | x7) : (~x6 | ~x7)));
  assign n1297 = x3 ? n1298 : (~n904 | ~n746);
  assign n1298 = (x0 | ((~x1 | x2 | ~x5 | x6) & (x1 | ~x2 | x5 | ~x6))) & (x1 | ~x5 | ((x2 | ~x6) & (~x0 | ~x2 | x6)));
  assign n1299 = ~x4 & (n1302 | (n1300 & n1301 & n733));
  assign n1300 = x6 & x7;
  assign n1301 = x3 & x5;
  assign n1302 = ~x1 & ((n547 & n1070) | (~x7 & ~n1303));
  assign n1303 = (~x0 | ~x2 | ~x3 | x5 | x6) & (x0 | ~x5 | (x2 ? (x3 | x6) : (~x3 | ~x6)));
  assign n1304 = n1305 & ~n1309 & (~x3 | ~n804 | ~n728);
  assign n1305 = n1308 & ((x3 & (x5 | n1307)) | (~x3 & ~x5 & n1306) | (x5 & n1307));
  assign n1306 = (x1 | ~x2 | x4) & (~x0 | ~x1 | x2 | ~x4);
  assign n1307 = (~x2 | ~x4 | ~x0 | x1) & (x0 | x2 | (~x1 ^ ~x4));
  assign n1308 = (~x0 | x1 | x2 | x4 | x5) & (x0 | ~x2 | ~x5 | (~x1 ^ x4));
  assign n1309 = ~n1312 & ((n743 & n1311) | (n1310 & ~n920));
  assign n1310 = ~x0 & ~x5;
  assign n1311 = x5 & ~x3 & ~x4;
  assign n1312 = x1 ^ x6;
  assign z039 = n1319 | ~n1329 | (~x2 & (~n1314 | ~n1324));
  assign n1314 = x0 ? (x1 | n1318) : (~n1316 & (x1 | n1315));
  assign n1315 = (x3 | ~x4 | ~x5 | x6 | x7) & (~x6 | ((x3 | x4 | x5 | ~x7) & (~x3 | (x4 ? (x5 | x7) : (~x5 | ~x7)))));
  assign n1316 = n1317 & (n830 | (x4 & n962));
  assign n1317 = x1 & ~x3;
  assign n1318 = (x4 | x5 | ~x6 | x7) & (~x4 | ~x5 | ~x7 | (x3 ^ ~x6));
  assign n1319 = x2 & (~n1321 | (~x1 & ~n1320));
  assign n1320 = (x0 | x3 | x4 | ~x5 | ~x6) & (x6 | ((x0 | ~x5 | (x3 ^ ~x4)) & (~x0 | ~x3 | ~x4 | x5)));
  assign n1321 = ~n1323 & (~n626 | ~n1322) & (~n577 | ~n699);
  assign n1322 = x6 & x3 & ~x5;
  assign n1323 = (x0 ^ x1) & (x3 ? (~x5 & x6) : (x5 & ~x6));
  assign n1324 = n1326 & (x3 | n1325);
  assign n1325 = (~x4 | (x0 ? (x1 ? (~x5 | ~x6) : (x5 | x6)) : (x5 | ~x6))) & (x0 | x4 | x6 | (~x1 ^ x5));
  assign n1326 = (~n825 | ~n1328) & (n1097 | (~n712 & n1327));
  assign n1327 = x0 ? (x3 | x4) : (~x3 | ~x4);
  assign n1328 = ~x4 & ~x5 & (~x1 | ~x6);
  assign n1329 = ~n1330 & (~x2 | (~n1333 & ~n1334 & n1336));
  assign n1330 = ~n765 & ((n1331 & n837) | (n1167 & ~n1332));
  assign n1331 = ~x6 & ~x3 & x4;
  assign n1332 = (~x3 | ~x6 | ~x1 | x2) & (x3 | x6 | x1 | ~x2);
  assign n1333 = ~n1008 & ((n841 & n761) | (n566 & ~n726));
  assign n1334 = ~n1335 & ~x7 & n653;
  assign n1335 = (x5 | x6 | ~x1 | x4) & (~x5 | ~x6 | x1 | ~x4);
  assign n1336 = (n1337 | n1338) & (~n662 | ~n712);
  assign n1337 = x4 ? (x5 | ~x7) : (~x5 | x7);
  assign n1338 = (x0 | ~x1 | ~x3 | x6) & (x3 | ~x6 | ~x0 | x1);
  assign z040 = ~n1340 | n1352 | (x7 & ~n1359);
  assign n1340 = n1349 & ~n1346 & ~n1341 & ~n1343;
  assign n1341 = x0 & (x1 ? (n1044 & n548) : ~n1342);
  assign n1342 = (~x3 | ((~x6 | x7 | x2 | ~x4) & (~x2 | x4 | (~x6 ^ x7)))) & (x6 | x7 | x2 | x4);
  assign n1343 = ~x0 & ((x7 & ~n1344) | (n683 & ~n1345));
  assign n1344 = (~x2 | ((~x4 | ~x6 | ~x1 | x3) & (x1 | x6 | (~x3 ^ ~x4)))) & (~x1 | x2 | (x3 ? (x4 | ~x6) : (~x4 | x6)));
  assign n1345 = (x1 | ~x6 | (x2 ^ ~x4)) & (~x1 | ~x2 | ~x4 | x6);
  assign n1346 = ~x0 & (x4 ? ~n1348 : ~n1347);
  assign n1347 = (x6 | ((x1 | x2 | ~x3 | ~x5) & (~x1 | (x2 ? (x3 | ~x5) : x5)))) & (~x2 | ~x3 | ~x6 | (x1 & x5));
  assign n1348 = (x1 | ~x2 | x3 | x5 | x6) & (~x3 | ((x1 | x2 | ~x5 | ~x6) & (~x1 | (x2 ? (~x5 | x6) : (x5 | ~x6)))));
  assign n1349 = (n981 | n1350) & (~n564 | n1351);
  assign n1350 = (x2 | x4 | x0 | x1) & (~x0 | (x1 ? (x2 | x4) : (~x2 | ~x4)));
  assign n1351 = (~x1 | x2 | x3 | x5 | ~x6) & (x1 | (x2 ? (x3 | x6) : (~x5 | ~x6)));
  assign n1352 = ~x7 & (n1354 | n1357 | (~n1353 & ~n1356));
  assign n1353 = x4 ^ x6;
  assign n1354 = ~x2 & (x0 ? (n689 & n592) : ~n1355);
  assign n1355 = (x1 | ~x3 | ~x4 | x5 | x6) & (x3 | ((x4 | ~x5 | x6) & (x5 | ~x6 | ~x1 | ~x4)));
  assign n1356 = (~x0 | ~x1 | x2 | x3 | x5) & (x0 | ~x3 | (x1 ? (x2 | ~x5) : (~x2 | x5)));
  assign n1357 = x2 & ((~n877 & ~n1211) | (n1358 & n1244));
  assign n1358 = ~x6 & x4 & x5;
  assign n1359 = ~n1363 & (x3 | n1360) & (n714 | n1362);
  assign n1360 = (x0 | n1361) & (~n895 | (~n704 & ~n1121));
  assign n1361 = (x1 | ~x4 | ~x5 | (~x2 ^ ~x6)) & (x4 | x5 | ((~x1 | ~x2 | x6) & (x2 | ~x6)));
  assign n1362 = (x0 | ~x3 | (x1 ? (~x2 | x6) : (x2 | ~x6))) & (~x0 | x1 | ~x2 | x3 | ~x6);
  assign n1363 = n1365 & ((n1364 & n859) | (~x2 & ~n1040));
  assign n1364 = x5 & x6;
  assign n1365 = x3 & x0 & ~x1;
  assign z041 = ~n1385 | n1382 | n1375 | n1367 | n1372;
  assign n1367 = ~x0 & (n1368 | (~x5 & n1044 & ~n1371));
  assign n1368 = x3 & ((x5 & ~n1369) | (n934 & ~n1370));
  assign n1369 = (x7 | ((~x4 | ~x6 | x1 | ~x2) & (x6 | (x1 ? (x2 ^ ~x4) : (x2 | x4))))) & (x2 | ~x6 | ~x7 | (x1 ^ x4));
  assign n1370 = (x1 | ~x4 | x6 | ~x7) & (~x1 | x4 | (~x6 ^ ~x7));
  assign n1371 = (~x6 | ~x7 | ~x1 | x4) & (x1 | ~x4 | (~x6 ^ ~x7));
  assign n1372 = ~x2 & (x0 ? ~n1373 : ~n1374);
  assign n1373 = (~x3 | ((x5 | x7 | ~x1 | x4) & (~x5 | ~x7 | x1 | ~x4))) & (~x1 | x3 | (x4 ? (x5 | ~x7) : (~x5 | x7))) & (x1 | x5 | (~x4 ^ x7));
  assign n1374 = ((x3 ^ ~x7) | (x1 ? (~x4 | x5) : (~x4 ^ ~x5))) & (~x1 | x4 | ((~x5 | ~x7) & (x3 | x5 | x7)));
  assign n1375 = x2 & (n1376 | n1378 | (~x5 & ~n1377));
  assign n1376 = ~n835 & ((~x0 & x1 & ~x4 & x5) | (~x1 & (x0 ? (x4 ^ ~x5) : (x4 & ~x5))));
  assign n1377 = x0 ? (x1 | ~x4 | (~x3 ^ x7)) : ((x3 | x4 | ~x7) & (~x1 | (x3 ? (x4 | x7) : ~x7)));
  assign n1378 = n1380 & ((n1379 & n927) | (~x1 & ~n1381));
  assign n1379 = x4 & ~x7;
  assign n1380 = ~x0 & x5;
  assign n1381 = x3 ? (x4 | x7) : (~x4 | ~x7);
  assign n1382 = n841 & (x4 ? ~n1384 : (n596 & n1383));
  assign n1383 = x5 & (x6 ^ ~x7);
  assign n1384 = (~x2 | ~x3 | ~x5 | x6 | x7) & (x2 | ~x6 | (x5 ? x3 : ~x7));
  assign n1385 = ~n1388 & (n643 | (~n1386 & (n1164 | n1387)));
  assign n1386 = n1287 & n837;
  assign n1387 = (x0 | ~x2 | ~x3 | x5) & (x3 | ~x5 | ~x0 | x2);
  assign n1388 = ~n1389 & ((~x2 & x5 & x6 & ~x7) | (x2 & ~x6 & (x5 ^ ~x7)));
  assign n1389 = (~x0 | x1 | ~x3 | x4) & (x0 | x3 | (~x1 ^ ~x4));
  assign z042 = n1404 | ~n1406 | (x5 ? ~n1391 : ~n1398);
  assign n1391 = ~n1394 & (~n1392 | ~n841 | (~n1393 & ~n1397));
  assign n1392 = ~x3 & x4;
  assign n1393 = ~x7 & x2 & x6;
  assign n1394 = ~x0 & ((n558 & n1395) | (x2 & ~n1396));
  assign n1395 = x7 & ~x4 & ~x6;
  assign n1396 = (x1 | x3 | ~x4 | ~x6 | x7) & (~x7 | (x1 ? (x3 ? (x4 | x6) : (~x4 | ~x6)) : (x3 ? (~x4 | x6) : (x4 | ~x6))));
  assign n1397 = ~x2 & (x6 ^ ~x7);
  assign n1398 = x4 ? n1401 : (x1 ? n1400 : n1399);
  assign n1399 = x0 ? ((x2 | x3 | ~x6 | x7) & (x6 | ~x7 | ~x2 | ~x3)) : ((x3 | x6 | ~x7) & (x2 | ~x3 | ~x6 | x7));
  assign n1400 = (~x3 | x6 | x7 | ~x0 | x2) & (x0 | x3 | (x2 ? (x6 | x7) : (~x6 | ~x7)));
  assign n1401 = x0 ? (~n804 | ~n1403) : n1402;
  assign n1402 = (~x1 | ~x2 | x3 | x6 | ~x7) & (x1 | ((x2 | ~x3 | ~x6 | ~x7) & (~x2 | x3 | x6 | x7)));
  assign n1403 = x7 & ~x3 & x6;
  assign n1404 = x1 & (x0 ? (n704 & n1044) : ~n1405);
  assign n1405 = (x3 | x4 | ~x5 | x6) & (x5 | ((~x2 | ((~x4 | ~x6) & (~x3 | x4 | x6))) & (x2 | ~x3 | x4 | ~x6)));
  assign n1406 = ~n1407 & ~n1412 & ~n1416 & (n1097 | n1415);
  assign n1407 = ~n1408 & ((~n1410 & n1411) | (~x1 & ~n1409));
  assign n1408 = x4 ^ ~x6;
  assign n1409 = (~x0 | ~x2 | (x3 ? (~x5 | ~x7) : (x5 | x7))) & (x0 | x2 | x3 | ~x5 | x7);
  assign n1410 = x2 ? (~x3 | x7) : (x3 | ~x7);
  assign n1411 = x5 & ~x0 & x1;
  assign n1412 = ~n1100 & (n1414 | (n626 & n1413));
  assign n1413 = ~x7 & x2 & x3;
  assign n1414 = ~x2 & ((~x0 & x1 & x3 & ~x7) | (x0 & (x1 ? (~x3 & ~x7) : (x3 & x7))));
  assign n1415 = (x2 | (x1 ? (~x4 | (x0 & x3)) : (~x3 | x4))) & (x1 | ((~x2 | ~x3 | ~x4) & (~x0 | x3 | x4)));
  assign n1416 = ~x1 & (~n1418 | (n653 & n1417));
  assign n1417 = ~x5 & x6 & (x2 ^ x4);
  assign n1418 = (~x2 | ((x3 | ~x4 | ~x5 | x6) & (~x3 | x4 | x5 | ~x6))) & (x2 | ~x3 | ~x4 | ~x5 | x6);
  assign z043 = n1434 | ~n1437 | (x6 ? ~n1420 : ~n1424);
  assign n1420 = x0 ? (x1 | n1422) : (x1 ? n1423 : n1421);
  assign n1421 = (x2 | ((~x5 | ~x7 | ~x3 | ~x4) & (x5 | x7 | x3 | x4))) & (~x5 | ~x7 | x3 | x4) & (~x2 | (x3 ? (x5 | (~x4 ^ ~x7)) : (~x5 | ~x7)));
  assign n1422 = (~x2 | ~x3 | (x4 ? (x5 | x7) : (~x5 | ~x7))) & (x3 | ~x4 | ~x7 | (x2 & ~x5));
  assign n1423 = (x3 | ((x2 | (x4 ? (x5 | x7) : (~x5 | ~x7))) & (~x5 | ~x7 | ~x2 | ~x4))) & (~x2 | ~x3 | x4 | (~x5 ^ ~x7));
  assign n1424 = (x1 & n1425) | (~n1430 & ~n1432 & ~x1 & ~n1428);
  assign n1425 = (n835 | n1426) & (x0 | n1427);
  assign n1426 = (x4 | x5 | ~x0 | x2) & (~x4 | ~x5 | x0 | ~x2);
  assign n1427 = (~x3 | ((~x2 | (x4 ? (x5 | x7) : (~x5 | ~x7))) & (x5 | x7 | x2 | x4))) & (x2 | x3 | ~x4 | (~x5 ^ ~x7));
  assign n1428 = n1429 & ((x0 & ~x4 & (~x2 | ~x3)) | (x4 & (x3 ? ~x0 : ~x2)));
  assign n1429 = ~x5 & ~x7;
  assign n1430 = ~n1010 & ((n526 & n1044) | (x3 & ~n1431));
  assign n1431 = (x5 | x7) & (~x2 | ~x5 | ~x7);
  assign n1432 = ~n1433 & x7 & n691;
  assign n1433 = x0 ? (~x3 | x4) : (x3 | ~x4);
  assign n1434 = ~n1008 & ((n596 & ~n1436) | (~x2 & ~n1435));
  assign n1435 = (~x6 | (x3 ? ((x1 | ~x4) & (x0 | (x1 & ~x4))) : (x0 ? (~x1 ^ ~x4) : (~x1 | x4)))) & (x1 | ~x4 | (x0 ? (x3 | x6) : ~x3));
  assign n1436 = x0 ? (x1 | (x4 & x6)) : (x4 | x6);
  assign n1437 = ~n1441 & (x0 ? n1438 : (~n1444 & ~n1448));
  assign n1438 = (~n728 | ~n1439) & (~n934 | n1440);
  assign n1439 = x3 & ~x1 & x2;
  assign n1440 = (x1 | ~x3 | x4 | ~x6) & (~x1 | x3 | (~x4 ^ x6));
  assign n1441 = ~n643 & (x4 ? (n742 & ~n1443) : ~n1442);
  assign n1442 = (~x0 | ((x1 | ~x2 | ~x3 | x5) & (~x1 | x2 | x3 | ~x5))) & (x0 | ~x1 | x2 | ~x3 | ~x5);
  assign n1443 = (x3 | x5) & (x1 | ~x3 | ~x5);
  assign n1444 = ~x3 & ((n772 & ~n1446) | (n1445 & ~n1447));
  assign n1445 = x1 & ~x4;
  assign n1446 = x2 ? (~x5 | x6) : (x5 | ~x6);
  assign n1447 = x2 ? (~x5 | ~x6) : (x5 | x6);
  assign n1448 = ~x5 & n927 & (x2 ? (x4 & x6) : (x4 ^ x6));
  assign z044 = ~n1462 | ~n1470 | (x4 ? ~n1450 : ~n1455);
  assign n1450 = ~n1452 & (~n1300 | ~n1451 | ~n733);
  assign n1451 = ~x3 & ~x5;
  assign n1452 = ~x6 & ((n746 & n1453) | (~x1 & ~n1454));
  assign n1453 = ~x7 & ~x3 & x5;
  assign n1454 = (x0 | ~x2 | ~x3 | ~x5 | x7) & (x5 | ((x0 | ~x2 | x3 | ~x7) & (x2 | (x0 ? (~x3 ^ ~x7) : (~x3 | x7)))));
  assign n1455 = x6 ? (~n1457 & (x2 | n1456)) : n1459;
  assign n1456 = (~x0 | ((~x5 | ~x7 | x1 | x3) & (~x1 | x5 | x7))) & (x5 | x7 | ~x1 | ~x3) & (x0 | ~x5 | ((x3 | x7) & (x1 | ~x3 | ~x7)));
  assign n1457 = n742 & ((n750 & n927) | (~x1 & n1458));
  assign n1458 = ~x5 & (~x3 ^ x7);
  assign n1459 = (~n560 | ~n1460) & (~n742 | n1461);
  assign n1460 = x7 & ~x3 & ~x5;
  assign n1461 = (x5 | x7 | ~x1 | ~x3) & (x1 | ~x5 | (~x3 ^ ~x7));
  assign n1462 = (n640 | n1463) & (n1353 | (~n1464 & ~n1466));
  assign n1463 = x0 ? ((x1 | ~x2 | ~x3 | x4) & (~x1 | x2 | x3 | ~x4)) : ((x1 | ~x2 | x3 | ~x4) & (~x1 | x2 | (~x3 ^ ~x4)));
  assign n1464 = x5 & (n1414 | (x2 & n543 & n1465));
  assign n1465 = ~x3 & x7;
  assign n1466 = n1467 & (n1469 | (x0 & n1468));
  assign n1467 = ~x1 & ~x5;
  assign n1468 = x2 & (x3 ^ ~x7);
  assign n1469 = x7 & x3 & ~x0 & ~x2;
  assign n1470 = x0 ? n1473 : (x1 ? n1471 : n1472);
  assign n1471 = x2 ? ((~x4 | x6 | ~x7) & (~x6 | (x3 ? (~x4 ^ x7) : (x4 | x7)))) : ((x3 | ~x4 | ~x6 | x7) & (~x3 | x4 | x6 | ~x7));
  assign n1472 = x2 ? ((~x3 | (x4 ? (x6 | ~x7) : (~x6 | x7))) & (x6 | ~x7 | x3 | x4)) : ((x3 | ~x7 | (~x4 ^ x6)) & (x7 | ((~x4 | ~x6) & (~x3 | x4 | x6))));
  assign n1473 = x1 ? (~n1044 | ~n1395) : n1474;
  assign n1474 = x3 ? (x7 | (x2 ? (~x4 | ~x6) : (~x4 ^ x6))) : (x2 ? (x4 ? (x6 | ~x7) : ~x6) : (x4 ? ~x6 : (x6 | x7)));
  assign z045 = ~n1492 | n1490 | n1486 | n1476 | n1483;
  assign n1476 = ~x0 & (n1478 | (n1477 & ~n1482));
  assign n1477 = x4 & ~x5;
  assign n1478 = x5 & (x7 ? (n1479 & ~n1480) : ~n1481);
  assign n1479 = x4 & ~x6;
  assign n1480 = x1 ? (~x2 | x3) : (x2 | ~x3);
  assign n1481 = (~x1 | ((~x2 | ~x4 | ~x6) & (x4 | x6 | x2 | x3))) & (~x6 | ((x3 | ~x4) & (x1 | ~x2 | ~x3 | x4)));
  assign n1482 = (~x3 | ((~x1 | ~x2 | ~x6 | x7) & (x1 | x2 | x6 | ~x7))) & (x1 | ~x2 | x3 | (~x6 ^ x7));
  assign n1483 = ~n640 & ((~n1134 & ~n1484) | (x4 & ~n1485));
  assign n1484 = (x0 | ~x1 | x2 | ~x3) & (~x0 | x3 | (x1 ^ ~x2));
  assign n1485 = (~x0 | x1 | x2 | x3 | x5) & (x0 | (x1 ? (~x2 | (~x3 ^ ~x5)) : (~x3 ^ x5)));
  assign n1486 = x0 & (n1487 | (n845 & n979));
  assign n1487 = ~x1 & ((n943 & n1489) | (x3 & ~n1488));
  assign n1488 = x4 ? (~x5 | ((~x6 | x7) & (~x2 | x6 | ~x7))) : (x5 | ((x6 | ~x7) & (x2 | ~x6 | x7)));
  assign n1489 = x4 & x2 & ~x3;
  assign n1490 = ~x7 & ((n1268 & n1209) | (~x4 & ~n1491));
  assign n1491 = (x1 | ((~x5 | ((x2 | ~x3) & (~x0 | (x2 & ~x3)))) & (x3 | x5 | x0 | ~x2))) & (x0 | ~x1 | (x2 ? (~x3 ^ x5) : (x3 | x5)));
  assign n1492 = ~n1497 & (~x7 | n1493) & (~n837 | ~n1500);
  assign n1493 = n1496 & (x4 ? n1494 : (~n622 | n1495));
  assign n1494 = (~x0 | x1 | x2 | x3 | ~x5) & (x0 | ((x1 | ~x2 | ~x3 | ~x5) & (~x1 | x2 | x3 | x5)));
  assign n1495 = x1 ? (x2 | ~x5) : (~x2 ^ ~x5);
  assign n1496 = (~x0 | x1 | ~x3 | ~x4 | x5) & (x0 | x4 | (x1 ? (~x3 | ~x5) : (~x3 ^ x5)));
  assign n1497 = ~x0 & ((n1498 & n951) | (~x2 & ~n1499));
  assign n1498 = ~x3 & x1 & x2;
  assign n1499 = (~x1 | ((~x3 | x5 | ~x6 | x7) & (x3 | ~x5 | x6 | ~x7))) & (x1 | x3 | x5 | ~x6 | x7);
  assign n1500 = ~x7 & x6 & ~x3 & ~x5;
  assign z046 = n1506 | ~n1512 | ~n1521 | (x0 & ~n1502);
  assign n1502 = ~n1505 & (x1 | (x2 & n1503) | (~x2 & n1504));
  assign n1503 = (x3 | ~x5 | (x4 ? (x6 | x7) : (~x6 | ~x7))) & (x5 | ((~x4 | ~x6 | ~x7) & (x6 | x7 | ~x3 | x4)));
  assign n1504 = (~x3 | ~x4 | ~x5 | x6 | x7) & (x4 | ~x6 | ~x7 | (x3 & ~x5));
  assign n1505 = n576 & n588;
  assign n1506 = ~n643 & (~n1508 | (x3 & ~n1507));
  assign n1507 = (x0 | ~x1 | ~x2 | ~x4 | ~x5) & (x4 | ((x0 | ~x1 | x2 | x5) & (~x0 | x1 | (~x2 ^ x5))));
  assign n1508 = ~n1510 & (x4 | (~n1509 & (n605 | ~n1511)));
  assign n1509 = ~x5 & (x0 ? (x1 & ~x2) : (x1 ^ ~x2));
  assign n1510 = x5 & x4 & ~x0 & ~x1;
  assign n1511 = ~x3 & x0 & ~x1;
  assign n1512 = ~n1517 & ((x4 & (x6 | n1516)) | (n1513 & (n1516 | (~x4 & ~x6))));
  assign n1513 = (x1 | n1514) & (x0 | ~x1 | ~x6 | n1515);
  assign n1514 = (x0 | x2 | x3 | ~x5 | ~x6) & (~x0 | x5 | x6 | (x2 ^ ~x3));
  assign n1515 = x2 ? (~x3 | ~x5) : (x3 | x5);
  assign n1516 = (~x5 | (x0 ? (x1 ? (x2 | x3) : (~x2 | ~x3)) : (~x1 | (~x2 ^ x3)))) & (x0 | x1 | ~x2 | x5);
  assign n1517 = n1518 & (x0 ? (~x1 & n1520) : (x1 & n1519));
  assign n1518 = ~x2 & x4;
  assign n1519 = ~x6 & ~x3 & x5;
  assign n1520 = ~x5 & (~x3 ^ x6);
  assign n1521 = ~n1522 & (x0 | (~x2 & n1524) | (x2 & n1528));
  assign n1522 = ~n640 & ((n639 & n1269) | (~x2 & ~n1523));
  assign n1523 = (x0 | ~x1 | ~x3 | ~x4 | x5) & (x3 | ((~x0 | ~x4 | (x1 ^ ~x5)) & (x0 | ~x1 | x4 | ~x5)));
  assign n1524 = x5 ? (x1 | (~n1525 & ~n1526)) : n1527;
  assign n1525 = ~x7 & ~x6 & ~x3 & x4;
  assign n1526 = x3 & (x4 ? (~x6 & ~x7) : (x6 & x7));
  assign n1527 = x1 ? ((x3 | ~x4 | ~x6 | ~x7) & (~x3 | x4 | x6 | x7)) : (x4 ? (x6 | x7) : (~x6 | ~x7));
  assign n1528 = x5 ? n1529 : (~x1 | (~n1525 & ~n1526));
  assign n1529 = (~x1 | ~x3 | ~x4 | x6 | x7) & (x1 | ~x6 | ~x7 | (~x3 ^ ~x4));
  assign z047 = n1531 | ~n1536 | ~n1550 | (~x1 & ~n1535);
  assign n1531 = ~x0 & ((~n1532 & n1533) | (~x3 & ~n1534));
  assign n1532 = x2 ^ ~x4;
  assign n1533 = ~x7 & ~x5 & x1 & x3;
  assign n1534 = (~x4 | ((~x5 | ~x7 | ~x1 | x2) & (x1 | x7 | (~x2 ^ ~x5)))) & (~x1 | x4 | ~x5 | (~x2 ^ ~x7));
  assign n1535 = (x0 | ~x2 | x5 | ~x7) & (~x3 | ~x5 | (x0 ? (~x2 ^ ~x7) : (~x2 | x7)));
  assign n1536 = ~n1544 & n1547 & (n1198 | (~n1537 & n1540));
  assign n1537 = ~x3 & ((n841 & ~n1538) | (n543 & n1539));
  assign n1538 = x2 ? (~x4 | x7) : (x4 | ~x7);
  assign n1539 = x4 & (~x2 ^ x7);
  assign n1540 = ~n1542 & (~n841 | ~n1413) & (~n1541 | n1543);
  assign n1541 = ~x4 & x3 & ~x0 & ~x2;
  assign n1542 = ~x0 & x7 & (x1 ? (x2 & x3) : (~x2 & ~x3));
  assign n1543 = x1 ^ ~x7;
  assign n1544 = x1 & ((n743 & n1545) | (~x0 & ~n1546));
  assign n1545 = x7 & ~x3 & x5;
  assign n1546 = (x5 | x7 | ~x2 | x3) & (~x5 | ~x7 | x2 | ~x3);
  assign n1547 = (~n880 | ~n830) & (n1548 | n1543 | ~n1549);
  assign n1548 = x3 ^ ~x4;
  assign n1549 = ~x5 & x0 & ~x2;
  assign n1550 = ~n1551 & (x1 | (~n1554 & n1557));
  assign n1551 = ~n1097 & ((n841 & ~n1553) | (~x0 & ~n1552));
  assign n1552 = x1 ? ((~x2 | ~x3 | ~x4 | x7) & (x4 | ~x7 | x2 | x3)) : (x7 | (x2 ? (x3 | x4) : ~x3));
  assign n1553 = x2 ? (x3 | ~x7) : (x3 ? (~x4 | ~x7) : x7);
  assign n1554 = ~x0 & ((n942 & n1556) | (~n1555 & n859));
  assign n1555 = (x6 | x7 | x3 | x5) & (~x6 | ~x7 | ~x3 | ~x5);
  assign n1556 = ~x4 & ~x2 & ~x3;
  assign n1557 = (n1558 | n1559) & (~n594 | ~n601);
  assign n1558 = x3 ? (x5 | ~x7) : (~x5 | x7);
  assign n1559 = (x0 | x2 | ~x4 | ~x6) & (x4 | x6 | ~x0 | ~x2);
  assign z048 = ~n1565 | ~n1571 | (~n640 & ~n1561);
  assign n1561 = (x0 | ~x1 | n1564) & (x1 | (n1563 & (~x0 | ~n1562)));
  assign n1562 = x4 & ~x2 & x3;
  assign n1563 = (x0 | ~x4 | (x2 ? (~x3 | ~x5) : (x3 | x5))) & (x4 | ((x0 | x2 | x3 | ~x5) & (~x0 | (x2 ? (x3 | x5) : (~x3 | ~x5)))));
  assign n1564 = x2 ? (x3 ^ ~x4) : (x3 | x4);
  assign n1565 = n1569 & (x1 | n1567) & (n1566 | n1568);
  assign n1566 = x3 ^ ~x5;
  assign n1567 = (x0 | ~x2 | ~x3 | x4 | x6) & (~x6 | ((x0 | x2 | ~x3 | x4) & (~x0 | x3 | (~x2 ^ ~x4))));
  assign n1568 = x0 ? (x4 | (x1 ? (x2 | x6) : (~x2 | ~x6))) : (x1 | ~x4 | (~x2 ^ x6));
  assign n1569 = (~n560 | ~n1203) & (~n804 | ~n1465 | n1570);
  assign n1570 = (x0 | x4 | x5 | ~x6) & (~x0 | ~x4 | ~x5 | x6);
  assign n1571 = ~n1572 & (n643 | (~n1575 & (x2 | n1574)));
  assign n1572 = x1 & ((n743 & n1331) | (~x0 & ~n1573));
  assign n1573 = (~x2 | (x3 ? (~x4 | ~x6) : (x4 | x6))) & (x2 | ~x3 | ~x4 | x6);
  assign n1574 = (x3 | (x0 ? (x5 | (~x1 ^ x4)) : (~x1 | ~x4))) & (x0 | ~x3 | (x1 ? x4 : (~x4 | ~x5)));
  assign n1575 = n570 & (x0 ? (x3 & (x4 | x5)) : (~x3 & (~x4 | ~x5)));
  assign z049 = ~n1579 | (~x2 & (x5 ? ~n1578 : ~n1577));
  assign n1577 = (x1 | ~x4 | ((x3 | ~x7) & (x0 | ~x3 | x7))) & (x4 | ((~x1 | x3 | ~x7) & (~x0 | ~x3 | x7)));
  assign n1578 = x0 ? (x4 | (x1 ? (x3 | x7) : (~x3 | ~x7))) : (x1 | ~x4 | (~x3 ^ ~x7));
  assign n1579 = ~n1582 & ~n1583 & ~n1584 & (n1580 | n1581);
  assign n1580 = x0 ? (x1 | ~x4) : (~x1 | x4);
  assign n1581 = (~x2 | x3 | x7) & (~x3 | ~x7);
  assign n1582 = ~n1164 & ((~x0 & ~n1205) | (n743 & n683));
  assign n1583 = n570 & ~n807 & (x3 ? (x5 ^ ~x7) : (~x5 ^ ~x7));
  assign n1584 = n1586 & ((n543 & n1395) | (n841 & n1585));
  assign n1585 = ~x7 & x4 & x6;
  assign n1586 = x5 & ~x2 & ~x3;
  assign z050 = ~n1590 | (x4 & ~n1588) | (~n1226 & ~n1589);
  assign n1588 = (x1 | x2 | x3 | (~x0 ^ x5)) & (x0 | ~x1 | (~x2 & ~x3 & x5));
  assign n1589 = x0 ? (x4 ^ ~x5) : (~x4 ^ ~x5);
  assign n1590 = (~n816 | ~n1228) & (~n804 | ~n1051 | n1591);
  assign n1591 = (x0 | x4 | x5 | ~x7) & (~x0 | ~x4 | ~x5 | x7);
  assign z051 = n1593 | ~n1596 | (n1586 & (~n1594 | ~n1595));
  assign n1593 = ~x2 & ((x1 & (x0 ? (~x3 & x5) : (x3 & ~x5))) | (x0 & ~x1 & (x3 ^ ~x5)));
  assign n1594 = (x0 | ~x1 | x4 | ~x6 | x7) & (~x0 | x1 | ~x4 | x6 | ~x7);
  assign n1595 = (~x4 | ~x6 | ~x0 | x1) & (x4 | x6 | x0 | ~x1);
  assign n1596 = (x1 | ~x2 | ~x5) & (x0 | ((~x1 | x5 | (~x2 & ~n1268)) & (~x5 | (x1 & (x2 | ~n1268)))));
  assign z052 = ~x6 & (~n1599 | (n816 & n1598));
  assign n1598 = x7 & ~x5 & ~x3 & ~x4;
  assign n1599 = n1601 & (~n1084 | (~n1600 & (~n876 | ~n922)));
  assign n1600 = x5 & ~x3 & ~x0 & ~x1;
  assign n1601 = (x0 & x1 & (x2 | x3)) | (~x0 & ~x1 & ~x2 & ~x3 & ~x4);
  assign z053 = ~x7 & (n1227 | ~n1599);
  assign z054 = ~x0 & (~n1226 | ~n1604 | (~n1605 & n1606));
  assign n1604 = (~n704 | ~n558) & (~n804 | (~n1392 & ~n1311));
  assign n1605 = x1 ? (~x3 | x7) : (x3 | ~x7);
  assign n1606 = ~x6 & ~x5 & ~x2 & ~x4;
  assign z055 = ~n1611 | (~x6 & ~n1608) | (~x2 & ~n1610);
  assign n1608 = (~n689 | n1609) & (~n757 | ~n774 | ~n733);
  assign n1609 = (~x0 | x2 | ~x4 | ~x5 | x7) & (x0 | x5 | (x2 ? (~x4 | x7) : (x4 | ~x7)));
  assign n1610 = (~x0 | x1 | x3 | ~x4 | x5) & (x0 | x4 | ~x5 | (~x1 ^ ~x3));
  assign n1611 = ~n1612 & ~n1613 & (~n681 | ~n1181 | ~n1614);
  assign n1612 = ~x0 & (x2 ? (x1 | (~x3 & ~x4)) : ((x3 & x4) | (~x1 & (x3 | x4))));
  assign n1613 = ~x4 & ~x3 & ~x2 & x0 & ~x1;
  assign n1614 = x6 & (x1 ^ ~x3);
  assign z056 = n1616 | ~n1618 | n1625 | (x2 & ~n1624);
  assign n1616 = ~x3 & ((n728 & n733) | (~x1 & ~n1617));
  assign n1617 = (x0 | ~x2 | ~x4 | x5 | ~x6) & (~x0 | ~x5 | (x2 ? (x4 | x6) : (~x4 | ~x6)));
  assign n1618 = n1620 & (~n543 | (~n1619 & ~n1622 & ~n1623));
  assign n1619 = x3 & (~x2 ^ ~x4);
  assign n1620 = (x0 | ~x1 | ~x2 | x3) & (x1 | (x0 ? (x2 | (~x3 & ~n1621)) : (~x2 | ~x3)));
  assign n1621 = x7 & ~x6 & x4 & x5;
  assign n1622 = ~x2 & ~x4 & (x3 ^ ~x5);
  assign n1623 = x3 & ((x2 & x4 & x5 & ~x6) | (~x5 & x6 & ~x2 & ~x4));
  assign n1624 = (~x0 | x1 | x3 | x4 | x5) & (x0 | ~x4 | (x1 ? (~x3 | x5) : (x3 | ~x5)));
  assign n1625 = ~x0 & ((n676 & n1626) | (n1017 & ~n1627));
  assign n1626 = x7 & ~x6 & x4 & ~x5;
  assign n1627 = (x3 | ~x5 | ~x6 | x7) & (x6 | ~x7 | ~x3 | x5);
  assign z057 = n1633 | ~n1638 | (~x0 & (~n1629 | ~n1637));
  assign n1629 = (n1631 | ~n1632) & (~x2 | n1630);
  assign n1630 = (x1 | x3 | ~x4 | x5 | ~x6) & (~x5 | ((~x1 | (x3 ? (~x4 | ~x6) : (x4 | x6))) & (x1 | ~x3 | ~x4 | x6)));
  assign n1631 = x1 ? (~x3 | ~x6) : (x3 ^ ~x6);
  assign n1632 = ~x5 & ~x2 & ~x4;
  assign n1633 = ~x0 & (n1634 | (n570 & n1636));
  assign n1634 = ~x4 & ((n558 & n951) | (x1 & ~n1635));
  assign n1635 = (x2 | ~x3 | x5 | x6 | ~x7) & (~x2 | x3 | ~x5 | ~x6 | x7);
  assign n1636 = x4 & ((x3 & x5 & x6 & ~x7) | (~x6 & x7 & ~x3 & ~x5));
  assign n1637 = (x4 | ((x1 | x2 | x3 | ~x5) & (~x1 | (x2 ? (x3 | x5) : (~x3 | ~x5))))) & (x1 | ~x2 | ~x4 | (~x3 ^ x5));
  assign n1638 = ~n1639 & ~n1640 & n1642 & (~n543 | ~n1562);
  assign n1639 = ~x1 & ((x2 & x3 & ~x4) | (~x3 & ((~x2 & x4) | (x0 & (~x2 | x4)))));
  assign n1640 = n1209 & n1641;
  assign n1641 = ~x5 & x3 & x4;
  assign n1642 = (~n1209 | ~n1643) & (~n610 | ~n1644);
  assign n1643 = x6 & x5 & ~x3 & ~x4;
  assign n1644 = x3 & x2 & x0 & ~x1;
  assign z058 = ~n1650 | (~x1 & (n1646 | (n525 & ~n1649)));
  assign n1646 = ~x0 & (x4 ? ~n1648 : (n1044 & ~n1647));
  assign n1647 = x5 ? (~x6 | x7) : (x6 | ~x7);
  assign n1648 = (x2 | ~x3 | ~x5 | x6 | x7) & (~x2 | ~x7 | (x3 ? (~x5 | ~x6) : (x5 | x6)));
  assign n1649 = (~x2 | ~x3 | ~x5 | x6 | ~x7) & (x2 | x5 | x7 | (~x3 ^ ~x6));
  assign n1650 = ~n1651 & n1655 & n1656 & (x0 | n1654);
  assign n1651 = ~x1 & (x0 ? ~n1652 : ~n1653);
  assign n1652 = (~x2 | x3 | x4 | ~x5 | ~x6) & (~x3 | ((~x2 | (x4 ? (~x5 | ~x6) : (x5 | x6))) & (x5 | x6 | x2 | ~x4)));
  assign n1653 = (~x2 | x3 | ~x4 | x5 | ~x6) & (x2 | x4 | ((x5 | ~x6) & (x3 | ~x5 | x6)));
  assign n1654 = (x1 | ~x2 | (x3 ? (x4 | x5) : (~x4 | ~x5))) & (x2 | ((x4 | x5 | ~x1 | x3) & (~x3 | (~x4 ^ x5))));
  assign n1655 = (x0 | ~x1 | ~x2 | x3 | ~x4) & (~x0 | ((x2 | x3 | x4) & (x1 | (x2 ? (x3 | ~x4) : x4))));
  assign n1656 = ~n543 | (n1657 & (x4 | n1658));
  assign n1657 = (x2 | x3 | x4 | ~x5 | x6) & (~x3 | ((~x2 | (x4 ? (~x5 | ~x6) : (x5 | x6))) & (x5 | ~x6 | x2 | x4)));
  assign n1658 = (x2 | ~x3 | x5 | x6 | ~x7) & (~x6 | ((~x2 | (x3 ? (x5 | x7) : (~x5 | ~x7))) & (x2 | x3 | ~x5 | x7)));
  assign z059 = n1660 | n1663 | ~n1671 | (x0 & ~n1670);
  assign n1660 = x1 & ((n600 & n830) | (~x0 & ~n1661));
  assign n1661 = (x4 | n1662) & (x7 | n1446 | x3 | ~x4);
  assign n1662 = (x2 | x6 | (x3 ? (x5 | ~x7) : (~x5 | x7))) & (~x6 | ~x7 | ((~x2 | ~x3 | x5) & (x3 | ~x5)));
  assign n1663 = ~x1 & (n1664 | n1667);
  assign n1664 = x5 & ((~x2 & ~n1665) | (n885 & ~n1666));
  assign n1665 = (x0 | x3 | x4 | ~x6 | ~x7) & (x6 | ((x0 | ~x3 | ~x4 | ~x7) & (~x0 | x7 | (x3 ^ ~x4))));
  assign n1666 = (~x0 | (x4 ? (x6 | ~x7) : (~x6 | x7))) & (~x6 | ~x7 | x0 | ~x4);
  assign n1667 = ~x5 & ((n594 & n1668) | (~x3 & ~n1669));
  assign n1668 = x7 & x4 & x6;
  assign n1669 = (x0 | ~x2 | x4 | ~x6 | x7) & (x6 | ((x0 | ~x2 | ~x4 | ~x7) & (~x0 | (x2 ? (x4 | x7) : (~x4 | ~x7)))));
  assign n1670 = (~x4 | ((x1 | (x2 ? (x3 | x5) : (~x3 | ~x5))) & (x3 | x5 | ~x1 | x2))) & (x1 | x2 | x4 | x5);
  assign n1671 = ~n1672 & ~n1674 & ~n1677 & (x0 | n1676);
  assign n1672 = ~x2 & ((n592 & n661) | (n543 & ~n1673));
  assign n1673 = (x5 | x6 | x3 | ~x4) & (~x3 | x4 | (~x5 ^ x6));
  assign n1674 = ~n1134 & (n1675 | (~x0 & ~x1 & ~n1011));
  assign n1675 = x0 & ((~x1 & x2 & x3 & x6) | (x1 & ~x2 & ~x3 & ~x6));
  assign n1676 = (x1 | ((~x3 | x4 | ~x5) & (x2 | x3 | ~x4 | x5))) & (~x2 | ((~x3 | x4 | ~x5) & (~x1 | x3 | ~x4 | x5))) & (~x1 | x2 | (x3 ? (~x4 | ~x5) : (x4 | x5)));
  assign n1677 = x2 & ((n543 & ~n928) | (n1678 & ~n1679));
  assign n1678 = ~x1 & (~x3 ^ ~x6);
  assign n1679 = x0 ? (x4 | ~x5) : (~x4 | x5);
  assign z060 = ~n1695 | (x5 ? (n1681 | ~n1684) : ~n1689);
  assign n1681 = x7 & ((~n1171 & ~n1682) | (~x0 & ~n1683));
  assign n1682 = x0 ? (x1 | ~x3) : (~x1 | x3);
  assign n1683 = (~x1 | ~x2 | ~x3 | x4 | x6) & (x1 | (x2 ? (x3 ? (~x4 | ~x6) : (x4 | x6)) : (x3 ? (~x4 | x6) : (x4 | ~x6))));
  assign n1684 = (n1685 | n1687) & (x7 | ~n1686 | n1688);
  assign n1685 = x2 ^ x4;
  assign n1686 = ~x0 & x6;
  assign n1687 = (x0 | ~x1 | x3 | x6 | ~x7) & (~x0 | x1 | (x3 ? (x6 | ~x7) : (~x6 | x7)));
  assign n1688 = (x1 | (x2 ? (~x3 | x4) : (x3 | ~x4))) & (~x3 | ~x4 | ~x1 | x2);
  assign n1689 = x1 ? n1692 : (~n1691 & (x7 | n1690));
  assign n1690 = x0 ? (x3 | (x2 ? (~x4 ^ x6) : (x4 | x6))) : (x2 ? (x3 ? (x4 | x6) : (~x4 | ~x6)) : (x3 ? (x4 | ~x6) : (~x4 | x6)));
  assign n1691 = x7 & n1051 & (x0 ? (~x2 ^ ~x4) : (x2 ^ ~x4));
  assign n1692 = (~n1693 | ~n1395) & (x7 | n1694);
  assign n1693 = x3 & ~x0 & ~x2;
  assign n1694 = (x2 | ((~x4 | x6 | x0 | ~x3) & (~x0 | (x3 ? (x4 | x6) : (~x4 | ~x6))))) & (x0 | ~x2 | ~x6 | (~x3 ^ ~x4));
  assign n1695 = n1700 & (~n841 | n1696) & (x0 | n1697);
  assign n1696 = (~x2 | ~x3 | x4 | x5 | ~x6) & (x3 | ((~x5 | (x2 ? (~x4 ^ x6) : (x4 | x6))) & (x5 | ~x6 | x2 | ~x4)));
  assign n1697 = x2 ? (x1 | (~n1698 & ~n1202)) : n1699;
  assign n1698 = x3 & (x4 ? (~x5 & x6) : (x5 & ~x6));
  assign n1699 = x1 ? (~x3 | (x4 ? (~x5 | x6) : ~x6)) : (x3 | (x4 ? (~x5 | x6) : (x5 | ~x6)));
  assign n1700 = (n1701 | n1702) & (n1097 | n1703);
  assign n1701 = x5 ? (x6 | x7) : (~x6 | ~x7);
  assign n1702 = (x2 | (x0 ? (x1 ? (x3 | x4) : (~x3 | ~x4)) : (x1 ? (x3 | ~x4) : (~x3 | x4)))) & (x0 | ~x2 | x4 | (~x1 & x3));
  assign n1703 = (~x4 | (x0 ? (x1 ? (x2 | x3) : (~x2 | ~x3)) : (x1 ? ~x2 : (x2 | ~x3)))) & (x2 | x4 | (x0 ? (x1 | ~x3) : (~x1 | x3)));
  assign z061 = n1720 | n1718 | n1715 | n1705 | n1710;
  assign n1705 = ~x2 & (n1706 | (n569 & ~n1709));
  assign n1706 = ~x6 & (x0 ? ~n1708 : ~n1707);
  assign n1707 = x1 ? (~x5 | (x3 ? (~x4 | ~x7) : (~x4 ^ x7))) : ((x3 | ~x4 | ~x5 | ~x7) & (x4 | (x3 ? (~x5 ^ ~x7) : (x5 | ~x7))));
  assign n1708 = (~x1 | ~x3 | x4 | x5 | ~x7) & (x1 | x3 | (x4 ? ~x5 : (x5 | ~x7)));
  assign n1709 = (~x0 | x1 | ~x3 | ~x4 | ~x5) & (x5 | ((x1 | ~x3 | x4) & (x0 | (x1 ? (x3 | x4) : ~x3))));
  assign n1710 = ~n640 & (~n1712 | (~x1 & ~n1711));
  assign n1711 = (x0 | ~x4 | (x2 ? (x3 | ~x5) : (~x3 | x5))) & (x4 | ((x0 | ~x2 | x3 | x5) & (~x0 | ~x5 | (~x2 ^ ~x3))));
  assign n1712 = ~n1713 & ~n1714 & (~n1268 | ~n746);
  assign n1713 = x1 & ((~x2 & ~x3 & ~x5) | (~x0 & x3 & (x2 ^ x5)));
  assign n1714 = ~x1 & (x0 ? (x2 ? (~x3 & x5) : (x3 & ~x5)) : (x5 & (x2 ^ ~x3)));
  assign n1715 = ~n643 & ((n1716 & n1269) | (~x2 & ~n1717));
  assign n1716 = ~x5 & x3 & ~x4;
  assign n1717 = (~x5 | ((x0 | x1 | ~x3 | ~x4) & (~x0 | x4 | (x1 ^ ~x3)))) & (~x4 | x5 | ((x1 | x3) & (x0 | ~x1 | ~x3)));
  assign n1718 = ~n1647 & ~n1719;
  assign n1719 = (~x2 | ((x1 | x3 | x4) & (x0 | (x1 ? (~x3 | ~x4) : x3)))) & (~x1 | x2 | ((x3 | ~x4) & (x0 | ~x3 | x4)));
  assign n1720 = x2 & (n1722 | ~n1724 | (~n1116 & ~n1721));
  assign n1721 = (x1 | ~x3 | ~x4) & (x3 | x4 | x0 | ~x1);
  assign n1722 = ~n1543 & n1723 & n539;
  assign n1723 = ~x5 & x6;
  assign n1724 = (~n712 | ~n1725) & (n1205 | n1408 | n814);
  assign n1725 = x7 & ~x6 & ~x4 & x5;
  assign z062 = ~n1743 | (x2 ? ~n1736 : ~n1727);
  assign n1727 = x4 ? (n1733 & (x1 | n1732)) : n1728;
  assign n1728 = ~n1731 & (x5 | n1729) & (n823 | n1730);
  assign n1729 = x6 ? (x7 | (x0 ? (~x1 | ~x3) : (x1 | x3))) : (~x7 | ((x1 | x3) & (~x0 | (x1 & x3))));
  assign n1730 = (x3 | ~x5 | x6 | ~x7) & (x5 | ~x6 | x7);
  assign n1731 = ~x0 & x3 & x5 & (x6 ^ x7);
  assign n1732 = (~x0 | ((x5 | ~x6 | ~x7) & (x3 | ~x5 | x7))) & (x5 | ((x3 | ~x6 | ~x7) & (x0 | ~x3 | (~x6 ^ x7))));
  assign n1733 = (~n658 | ~n1734) & (n640 | n1735);
  assign n1734 = ~x3 & x0 & x1;
  assign n1735 = (~x1 | x3 | x5) & (~x5 | (x0 ? (x1 | ~x3) : (~x1 ^ ~x3)));
  assign n1736 = x4 ? (~n1737 & ~n1738) : (~n1739 & ~n1740);
  assign n1737 = ~n643 & (x0 ? (~x1 & (x3 ^ ~x5)) : (~x3 & (x1 | x5)));
  assign n1738 = n825 & ((~x5 & ~x6 & ~x7) | (~x1 & ((~x6 & ~x7) | (~x5 & x6 & x7))));
  assign n1739 = ~n640 & (x0 ? (~x1 & x3) : ((~x3 & ~x5) | (x1 & x3 & x5)));
  assign n1740 = ~x1 & (n1742 | (~x0 & n1741));
  assign n1741 = ~x6 & (x3 ? (~x5 & x7) : (x5 & ~x7));
  assign n1742 = ~x7 & x6 & x5 & x0 & ~x3;
  assign n1743 = n1750 & (x2 | n1745) & (n1744 | n1749);
  assign n1744 = x3 ^ x4;
  assign n1745 = x1 ? (x0 | (~n1746 & ~n1748)) : n1747;
  assign n1746 = x6 & ~x3 & x5;
  assign n1747 = (x0 | ~x3 | x4 | x5 | ~x6) & (x6 | ((x3 | ~x4 | x5) & (~x0 | ((~x4 | x5) & (~x3 | x4 | ~x5)))));
  assign n1748 = ~x6 & ~x5 & x3 & x4;
  assign n1749 = (x0 | ~x5 | (x1 ? (~x2 | ~x6) : (x2 | x6))) & (~x0 | x1 | ~x2 | x5 | ~x6);
  assign n1750 = (n1353 | n1751) & (x3 | ~n570 | n1752);
  assign n1751 = (~x0 | ~x1 | x2 | x3 | ~x5) & (x0 | ~x2 | ~x3 | (x1 ^ ~x5));
  assign n1752 = (x0 | ~x6 | (x4 ^ ~x5)) & (~x0 | ~x4 | ~x5 | x6);
  assign z063 = n1760 | ~n1765 | ~n1768 | (~x7 & ~n1754);
  assign n1754 = ~n1758 & (~x6 | (n1756 & (x1 | n1755)));
  assign n1755 = x2 ? ((x4 | x5 | x0 | x3) & (~x0 | ((x4 | ~x5) & (x3 | ~x4 | x5)))) : ((~x3 | ~x4 | x5) & (x0 | ((~x3 | x4 | ~x5) & (~x4 | x5))));
  assign n1756 = (~n1268 | ~n746) & (n1134 | n1757);
  assign n1757 = (~x2 | ~x3 | ~x0 | x1) & (x0 | (x1 ? (~x2 ^ x3) : (x2 | x3)));
  assign n1758 = n560 & n1759;
  assign n1759 = ~x6 & x5 & ~x3 & x4;
  assign n1760 = ~n640 & (n1762 | n1764 | (~x1 & ~n1761));
  assign n1761 = x3 ? ((x0 | x2 | ~x4 | x5) & (~x0 | ~x2 | x4 | ~x5)) : (x0 ? (x2 ? (~x4 | x5) : (x4 | ~x5)) : (~x5 | (~x2 ^ x4)));
  assign n1762 = ~n1134 & (n880 | (n742 & ~n1763));
  assign n1763 = x1 ^ ~x3;
  assign n1764 = n746 & n1641;
  assign n1765 = (n1014 | n1766) & (n1134 | n1767);
  assign n1766 = (x0 | x1 | ~x2 | ~x3) & (x2 | x3 | ~x0 | ~x1);
  assign n1767 = (x0 | ~x1 | ~x2 | ~x3 | ~x7) & (x1 | ((~x3 | ~x7 | x0 | x2) & (~x0 | (x2 ? (x3 | ~x7) : (~x3 | x7)))));
  assign n1768 = ~n1773 & ~n1776 & (~n1769 | n1770);
  assign n1769 = ~x6 & x7;
  assign n1770 = (x1 | n1771) & (~x1 | x2 | ~n681 | n1772);
  assign n1771 = x2 ? (~x5 | (x0 ? (x3 | x4) : (~x3 | ~x4))) : (~x4 | ((x3 | x5) & (~x0 | (x3 & x5))));
  assign n1772 = x0 & ~x3;
  assign n1773 = ~x2 & ((~x4 & ~n1774) | (n1012 & ~n1775));
  assign n1774 = (x0 | ~x1 | ~x5 | x7) & (x1 | ((~x5 | ~x7 | x0 | x3) & (~x0 | (x3 ? (~x5 | ~x7) : (x5 | x7)))));
  assign n1775 = x3 ? (x5 | ~x7) : (~x5 ^ ~x7);
  assign n1776 = x2 & (x0 ? (n1188 & n635) : ~n1777);
  assign n1777 = (x1 | x3 | ~x4 | x5 | ~x7) & (~x5 | ((x1 | x3 | ~x4 | x7) & (~x1 | x4 | (x3 ^ ~x7))));
  assign z064 = ~n1787 | ~n1798 | (~x1 & (n1779 | ~n1782));
  assign n1779 = x0 & ((n1070 & n1780) | (n1301 & ~n1781));
  assign n1780 = ~x4 & x2 & ~x3;
  assign n1781 = (x2 | ~x6 | ~x7) & (~x4 | ((~x6 | ~x7) & (~x2 | x6 | x7)));
  assign n1782 = n1785 & (~n588 | ~n1783) & (n1198 | n1784);
  assign n1783 = ~x3 & ~x0 & x2;
  assign n1784 = (x0 | ~x2 | ~x3 | ~x4 | x7) & (~x0 | x2 | x3 | x4 | ~x7);
  assign n1785 = (~n549 | ~n1786) & (~n1300 | ~n653 | n1685);
  assign n1786 = ~x7 & ~x4 & ~x6;
  assign n1787 = ~n1788 & ~n1795 & (n714 | n1791);
  assign n1788 = ~n643 & (x2 ? ~n1790 : ~n1789);
  assign n1789 = (x0 | ((~x1 | (x3 ? (x4 | ~x5) : x5)) & (x5 | ((x3 | x4) & (x1 | ~x3 | ~x4))))) & (~x4 | ~x5 | x1 | x3) & (~x0 | (x1 ? (x4 | (~x3 ^ x5)) : (~x4 | (x3 & ~x5))));
  assign n1790 = (x1 | (x3 ? (x4 | ~x5) : (~x4 | x5))) & (x0 | ~x1 | (~x4 ^ ~x5));
  assign n1791 = (~n1792 | ~n1269) & (x2 | n1793 | n1794);
  assign n1792 = x7 & x3 & x6;
  assign n1793 = x1 ? (~x6 | ~x7) : (x6 | x7);
  assign n1794 = x0 ^ ~x3;
  assign n1795 = x2 & ((~x0 & ~n1796) | (n841 & ~n1797));
  assign n1796 = x1 ? ((~x5 | ~x6 | x3 | x4) & (x5 | x6 | ~x3 | ~x4)) : (x4 | x6 | (~x3 ^ x5));
  assign n1797 = (~x3 | ~x4 | x5 | ~x6) & (x3 | ~x5 | (~x4 ^ ~x6));
  assign n1798 = ~n1799 & (~n543 | (x4 & n1802) | (~x4 & n1803));
  assign n1799 = ~x2 & ((~n1134 & ~n1800) | (~x5 & ~n1801));
  assign n1800 = (x0 | x1 | ~x3 | ~x6) & (x3 | x6 | ~x0 | ~x1);
  assign n1801 = (x0 | ~x1 | ~x3 | x4 | x6) & (x1 | ((x0 | x3 | ~x4 | x6) & (~x0 | ~x3 | (~x4 ^ x6))));
  assign n1802 = x2 ? ((x3 | x6 | x7) & (~x6 | ~x7 | ~x3 | ~x5)) : ((x3 | ~x6 | ~x7) & (x6 | x7 | ~x3 | ~x5));
  assign n1803 = (x3 | x7 | ((x5 | x6) & (x2 | ~x5 | ~x6))) & (~x2 | ~x3 | ~x6 | ~x7);
  assign z065 = ~n1816 | n1813 | n1805 | n1810;
  assign n1805 = ~x0 & (n1806 | (n570 & ~n1809));
  assign n1806 = x1 & (x3 ? ~n1808 : ~n1807);
  assign n1807 = (~x2 | ~x4 | ~x5 | x6 | ~x7) & (x4 | x7 | ((x5 | ~x6) & (x2 | ~x5 | x6)));
  assign n1808 = (~x6 | ~x7 | ~x4 | ~x5) & (~x2 | x5 | x6 | (~x4 ^ ~x7));
  assign n1809 = (x3 | x4 | x5 | ~x6 | ~x7) & (~x3 | ((~x5 | ~x6 | ~x7) & (x6 | x7 | x4 | x5)));
  assign n1810 = ~n1008 & (x2 ? ~n1812 : ~n1811);
  assign n1811 = (x6 | ((~x3 | ((x1 | ~x4) & (x0 | (x1 & ~x4)))) & (~x0 | x3 | (~x1 & x4)))) & (x0 | x3 | ~x6 | (~x1 ^ ~x4));
  assign n1812 = (x1 | ((~x0 | x4 | (~x3 ^ ~x6)) & (~x4 | x6 | x0 | ~x3))) & (x0 | ~x6 | ((x3 | ~x4) & (~x1 | ~x3 | x4)));
  assign n1813 = x2 & ((~n823 & ~n1814) | (~x1 & ~n1815));
  assign n1814 = (~x3 | ~x4 | ~x5 | x7) & (x3 | (x4 ? (x5 | x7) : (~x5 | ~x7)));
  assign n1815 = (x0 | x3 | x4 | x5 | x7) & (~x3 | ((x5 | ~x7 | ~x0 | ~x4) & (x0 | x4 | (~x5 ^ x7))));
  assign n1816 = ~n1817 & (n1014 | n1823) & (x2 | n1819);
  assign n1817 = n841 & (~n996 | (n778 & ~n1818));
  assign n1818 = x3 ? (~x5 | (~x4 ^ ~x7)) : (~x4 | x7);
  assign n1819 = x0 ? n1822 : (~n1821 & (n1008 | n1820));
  assign n1820 = x1 ? (~x3 | x4) : (x3 | ~x4);
  assign n1821 = x7 & x5 & x4 & ~x1 & x3;
  assign n1822 = x1 ? ((x3 | ~x4 | ~x5 | ~x7) & (~x3 | x4 | x5 | x7)) : (x4 | ~x7 | (~x3 ^ x5));
  assign n1823 = x0 ? ((x1 | ~x2 | ~x3 | x6) & (~x1 | x2 | x3 | ~x6)) : ((x1 | x3 | x6) & (x2 | (~x3 ^ ~x6)));
  assign z066 = ~n1844 | n1840 | ~n1833 | n1825 | n1830;
  assign n1825 = ~x3 & ((~x1 & ~n1826) | (n543 & ~n1829));
  assign n1826 = (~x4 | n1827) & (x0 | x4 | ~x5 | n1828);
  assign n1827 = (~x0 | x2 | x5 | x6 | ~x7) & (~x5 | ((x0 | ~x2 | ~x6 | x7) & (~x0 | (x2 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n1828 = x2 ? (~x6 ^ ~x7) : (~x6 | x7);
  assign n1829 = (~x7 | (x2 ? (x5 | (~x4 ^ ~x6)) : (~x5 | (~x4 ^ x6)))) & (x5 | x7 | (x2 ? (~x4 | x6) : (x4 | ~x6)));
  assign n1830 = x3 & (~n1832 | (~n1097 & ~n1831));
  assign n1831 = (~x2 | x4 | x7 | ~x0 | x1) & (x0 | ((~x1 | x2 | ~x4 | x7) & (x1 | ~x2 | x4 | ~x7)));
  assign n1832 = (~n560 | ~n817) & (x0 | n640 | n1284);
  assign n1833 = ~n1837 & (x2 | (~n1834 & ~n1836));
  assign n1834 = n1835 & (x0 ? (x1 ? (~x3 & ~x7) : (x3 & x7)) : (x1 ? (~x3 & x7) : (x3 & ~x7)));
  assign n1835 = ~x4 & ~x6;
  assign n1836 = ~x7 & n597 & ((x1 & ~x3) | (~x0 & ~x1 & x3));
  assign n1837 = ~n643 & ((n841 & ~n1839) | (~x0 & ~n1838));
  assign n1838 = (~x1 | ~x2 | ~x3 | x4 | ~x5) & (x1 | x2 | x3 | ~x4 | x5);
  assign n1839 = (x3 | x4 | ~x5) & (~x2 | ~x3 | ~x4 | x5);
  assign n1840 = ~x0 & ((n804 & ~n1841) | n1842 | n1843);
  assign n1841 = (x3 | (x4 ? (~x5 | x6) : (x5 | ~x6))) & (~x5 | ~x6 | ~x3 | x4);
  assign n1842 = ~n1353 & ((n876 & n632) | (~x1 & n1194));
  assign n1843 = n728 & n1498;
  assign n1844 = n1847 & (~n841 | n1845) & (n1040 | n1846);
  assign n1845 = (~x6 | ((x4 | x5 | ~x2 | ~x3) & (x2 | (x3 ? (~x4 | ~x5) : (x4 | x5))))) & (~x2 | ~x4 | x6 | (~x3 ^ ~x5));
  assign n1846 = x1 ? ((x0 | ~x2 | x7) & (x3 | ~x7 | ~x0 | x2)) : ((~x2 ^ x3) | (~x0 ^ x7));
  assign n1847 = (n981 | n1848) & (~n1300 | ~n1029 | ~n746);
  assign n1848 = (~x2 | ~x4 | x0 | ~x1) & (~x0 | x2 | (~x1 ^ x4));
  assign z067 = n1851 | n1859 | ~n1865 | (~n1850 & ~n1864);
  assign n1850 = x4 ? (x6 | ~x7) : (~x6 | x7);
  assign n1851 = ~x5 & (n1852 | ~n1856 | (~n682 & ~n1855));
  assign n1852 = x7 & (x6 ? ~n1853 : (n1145 & ~n1854));
  assign n1853 = x0 ? (x1 | (x2 ? (x3 | x4) : (~x3 | ~x4))) : (~x1 | ~x4 | (~x2 ^ ~x3));
  assign n1854 = x0 ? (~x2 | ~x3) : (x2 | x3);
  assign n1855 = (~x0 | x2 | x3 | ~x4 | x7) & (x0 | ((x2 | ~x3 | ~x4 | ~x7) & (~x2 | x4 | (~x3 ^ x7))));
  assign n1856 = (n1312 | n1858) & (~n1029 | ~n560 | ~n1857);
  assign n1857 = ~x6 & ~x7;
  assign n1858 = (x0 | ~x3 | (x2 ? (x4 | ~x7) : (~x4 | x7))) & (~x0 | x2 | x3 | ~x4 | ~x7);
  assign n1859 = x5 & ((~x1 & ~n1860) | (n543 & ~n1863));
  assign n1860 = x2 ? n1862 : (~n1861 & (n604 | ~n898));
  assign n1861 = x7 & x6 & ~x4 & ~x0 & ~x3;
  assign n1862 = (~x6 | ~x7 | ~x3 | x4) & (x6 | x7 | x3 | ~x4);
  assign n1863 = x2 ? ((x3 | ~x4 | ~x6 | x7) & (~x3 | x4 | x6 | ~x7)) : ((x3 | x4 | ~x6 | x7) & (~x3 | (x4 ? (~x6 | ~x7) : (x6 | x7))));
  assign n1864 = (~x0 | ((x1 | ~x2 | ~x3 | x5) & (~x1 | x2 | x3 | ~x5))) & (x1 | x2 | ((~x3 | ~x5) & (x0 | x3 | x5)));
  assign n1865 = ~n1868 & (~n841 | n1866) & (n1205 | n1867);
  assign n1866 = (x2 | ~x3 | x4 | x5 | ~x7) & (x3 | ((x2 | ~x5 | (~x4 ^ x7)) & (x5 | x7 | (~x2 & x4))));
  assign n1867 = x1 ? ((x2 | x4 | x5) & (x0 | ~x4 | (~x2 ^ x5))) : (~x2 | ~x5);
  assign n1868 = ~x0 & ((~n1090 & ~n1869) | (n683 & ~n1870));
  assign n1869 = (x2 | ~x3 | x4 | ~x7) & (~x2 | (x3 ? (~x4 | ~x7) : (x4 | x7)));
  assign n1870 = (~x1 | x2 | ~x4 | x5) & (x1 | (x2 ? (~x4 | x5) : ~x5));
  assign z068 = n1877 | n1880 | ~n1883 | (~x2 & ~n1872);
  assign n1872 = ~n1876 & (x3 | (~n1874 & (~x1 | n1873)));
  assign n1873 = (~x4 | ((~x6 | ~x7 | ~x0 | ~x5) & (x0 | x5 | (~x6 ^ ~x7)))) & (~x0 | x4 | ~x5 | (~x6 ^ x7));
  assign n1874 = n772 & ((n1769 & n1875) | (~x0 & n659));
  assign n1875 = x0 & x5;
  assign n1876 = n852 & ((x4 & x5 & x7) | (~x1 & ~x4 & ~x7));
  assign n1877 = ~n823 & (x5 ? ~n1878 : ~n1879);
  assign n1878 = (~x2 | x3 | ~x4 | (~x6 ^ x7)) & (x4 | ((~x2 | ~x3 | ~x6 | ~x7) & (x2 | ((x6 | ~x7) & (~x3 | ~x6 | x7)))));
  assign n1879 = (x2 | x3 | x4 | ~x6 | x7) & (~x2 | ((~x6 | ~x7 | ~x3 | ~x4) & (x3 | x4 | (~x6 ^ ~x7))));
  assign n1880 = x5 & ((~n1744 & ~n1881) | (~x0 & ~n1882));
  assign n1881 = (x0 | ~x1 | ~x2 | x6) & (~x0 | x1 | (~x2 ^ x6));
  assign n1882 = (x1 | ~x2 | ~x3 | ~x4 | x6) & (x2 | x3 | ((~x4 | x6) & (~x1 | x4 | ~x6)));
  assign n1883 = ~n1884 & ~n1886 & ~n1889 & (n1353 | n1888);
  assign n1884 = n1885 & ((n828 & n813) | (x7 & ~n1841));
  assign n1885 = x2 & ~x0 & ~x1;
  assign n1886 = ~n627 & ((n816 & n867) | (n1429 & ~n1887));
  assign n1887 = (x2 | x4 | ~x0 | ~x1) & (~x2 | ~x4 | (x0 & x1));
  assign n1888 = (x0 | ((x2 | ~x3 | x5) & (x1 | ~x2 | x3 | ~x5))) & (x2 | x5 | (x3 ? x1 : ~x0));
  assign n1889 = ~x5 & ((~n615 & n1890) | (~n682 & n1891));
  assign n1890 = x2 & (~x0 | ~x1);
  assign n1891 = ~x4 & ~x3 & ~x0 & ~x2;
  assign z069 = n1896 | ~n1904 | (x2 ? ~n1900 : ~n1893);
  assign n1893 = n1895 & (x3 | n1894);
  assign n1894 = (x1 | ~x4 | x7 | (~x0 & ~x5)) & (x0 | ~x7 | ((~x4 | x5) & (~x1 | x4 | ~x5)));
  assign n1895 = (x0 & x3 & (x1 | ~n867)) | (~n670 & ~n867) | (~x3 & (~x0 | ~x1));
  assign n1896 = ~x2 & (x0 ? ~n1897 : ~n1899);
  assign n1897 = x1 ? (~n774 | ~n951) : (n1898 & (~n774 | ~n942));
  assign n1898 = (x3 | x4 | x6 | ~x7) & (~x3 | ~x4 | ~x6 | x7);
  assign n1899 = (x1 | x3 | x4 | ~n942) & (~x1 | (x3 ? (x4 | ~n942) : n1113));
  assign n1900 = ~n1902 & (x0 ? (~n1188 | ~n635) : n1901);
  assign n1901 = (~x1 | ~x3 | ~x4 | x5 | ~x7) & (x3 | x4 | ((~x5 | x7) & (x1 | x5 | ~x7)));
  assign n1902 = ~n1134 & ((~n1205 & ~n823) | (n626 & n1903));
  assign n1903 = x3 & ~x7;
  assign n1904 = (n640 | (~n1905 & ~n1906)) & (~n570 | n1907);
  assign n1905 = ~n710 & (x2 ? ~n856 : (x3 & ~n1134));
  assign n1906 = n1044 & ((x0 & ((~x4 & ~x5) | (x1 & x4 & x5))) | (~x4 & ((x1 & ~x5) | (~x0 & ~x1 & x5))));
  assign n1907 = (~n978 | ~n1908) & (~n1910 | (~n959 & ~n1909));
  assign n1908 = ~x4 & x0 & ~x3;
  assign n1909 = x3 & (~x4 ^ ~x5);
  assign n1910 = x7 & ~x0 & ~x6;
  assign z070 = n1912 | ~n1919 | ~n1927 | (~n643 & ~n1914);
  assign n1912 = n689 & (x0 ? (n859 & n951) : ~n1913);
  assign n1913 = (x2 | ~x4 | ~x5 | ~x6 | ~x7) & (~x2 | ((x4 | ~x6 | ~x7) & (x6 | x7 | ~x4 | ~x5)));
  assign n1914 = ~n1915 & (~n731 | ~n560) & (n1566 | n1918);
  assign n1915 = ~x0 & (n1917 | (~x4 & ~n1916));
  assign n1916 = x2 ? (x3 | x5) : (~x3 | ~x5);
  assign n1917 = ~x5 & x4 & ~x3 & ~x1 & ~x2;
  assign n1918 = x4 ? (~x2 | (x0 & x1)) : (x2 | (~x0 & ~x1));
  assign n1919 = ~n1921 & n1924 & (n1926 | (n1920 & n1566));
  assign n1920 = x3 ? (~x4 | ~x5) : (x4 | x5);
  assign n1921 = ~n1134 & (n1923 | (~n784 & n1922));
  assign n1922 = x3 & ~x0 & ~x1;
  assign n1923 = ~x6 & ~x3 & ~x2 & x0 & x1;
  assign n1924 = (~n588 | ~n733) & (~n1209 | (~n662 & ~n1925));
  assign n1925 = x7 & x6 & x3 & ~x5;
  assign n1926 = (~x0 | x1 | x2 | x6 | x7) & (x0 | ~x1 | ~x2 | ~x6 | ~x7);
  assign n1927 = ~n1928 & ~n1930 & n1933 & (n856 | n1184);
  assign n1928 = ~n714 & ((~n1794 & ~n1929) | (n1792 & n816));
  assign n1929 = (~x6 | ~x7 | ~x1 | x2) & (x6 | x7 | x1 | ~x2);
  assign n1930 = ~n1932 & (n1931 | (n543 & n1518));
  assign n1931 = ~x4 & x2 & x0 & ~x1;
  assign n1932 = x3 ? (~x5 | x6) : (x5 | ~x6);
  assign n1933 = (n1934 | ~n626 | ~n1051) & (~n1250 | n1935);
  assign n1934 = x2 ? (~x4 | x5) : (x4 | ~x5);
  assign n1935 = (x1 | x5 | ~x6 | ~x7) & (x6 | x7 | ~x1 | ~x5);
  assign z071 = x3 ? (~n1945 | ~n1956) : (~n1937 | ~n1959);
  assign n1937 = (x2 | n1942) & (~x2 | n1938) & (n1218 | n1941);
  assign n1938 = (n640 | n1939) & (x1 | n1940);
  assign n1939 = (~x4 | ~x5 | ~x0 | x1) & (x4 | x5 | x0 | ~x1);
  assign n1940 = (~x0 | x4 | ~x5 | ~x6 | ~x7) & (x0 | ((x4 | ~x7 | (~x5 ^ x6)) & (x7 | ((~x5 | ~x6) & (~x4 | x5 | x6)))));
  assign n1941 = (~x6 | ((x2 | ~x5 | ~x0 | x1) & (x0 | (x1 ? ~x5 : (x2 | x5))))) & (~x0 | x5 | x6 | (x1 & x2));
  assign n1942 = x0 ? n1943 : (x6 ? n1944 : n1014);
  assign n1943 = (x6 | x7 | ~x4 | ~x5) & (~x6 | ((x1 | x4 | x5 | ~x7) & (~x1 | (x4 ? (x5 | x7) : (~x5 | ~x7)))));
  assign n1944 = (x1 | ~x4 | ~x5 | x7) & (x5 | ~x7 | ~x1 | x4);
  assign n1945 = n1955 & ~n1953 & ~n1951 & ~n1946 & ~n1949;
  assign n1946 = ~x1 & ((n951 & n1948) | (x2 & ~n1947));
  assign n1947 = (x0 | x4 | ~x5 | x6 | x7) & (~x0 | ~x4 | x5 | (~x6 ^ ~x7));
  assign n1948 = x4 & ~x0 & ~x2;
  assign n1949 = ~x1 & ((n525 & n978) | (~x0 & n1950));
  assign n1950 = ~x4 & x7 & (x5 ^ ~x6);
  assign n1951 = ~n1198 & ~n1952;
  assign n1952 = (x1 | x2 | (x0 ? (~x4 ^ ~x7) : (~x4 | x7))) & (x0 | ~x1 | ((x4 | x7) & (~x2 | ~x4 | ~x7)));
  assign n1953 = ~n1116 & (n1931 | (~x0 & x4 & ~n1954));
  assign n1954 = x1 ^ ~x2;
  assign n1955 = (~n529 | ~n951) & (~n1364 | ~n543 | n1538);
  assign n1956 = (n1014 | n1957) & (x2 | n1958);
  assign n1957 = x0 ? (x1 | x2) : (~x1 | ~x2);
  assign n1958 = (x0 | x1 | ~x5 | (~x4 ^ ~x7)) & (~x0 | ~x1 | x4 | x5 | x7);
  assign n1959 = ~n1960 & ~n1962 & (x5 | n1218 | ~n1885);
  assign n1960 = ~n1008 & ~n1961;
  assign n1961 = x0 ? (x4 | (x1 ^ ~x2)) : (~x1 | ~x4);
  assign n1962 = n632 & ((n525 & n526) | (n1429 & n1167));
  assign z072 = n1984 | n1981 | ~n1975 | n1964 | ~n1970;
  assign n1964 = ~x1 & (n1965 | n1968 | n1969);
  assign n1965 = ~x0 & ((n934 & ~n1898) | (n1966 & ~n1967));
  assign n1966 = x2 & x5;
  assign n1967 = (x6 | x7 | x3 | x4) & (~x6 | ~x7 | ~x3 | ~x4);
  assign n1968 = ~n1040 & ((~x3 & ~x7 & x0 & ~x2) | (~x0 & x7 & (~x2 ^ ~x3)));
  assign n1969 = n526 & n564 & (x2 ? (x3 & x6) : ~x6);
  assign n1970 = ~n1971 & (n981 | n1974);
  assign n1971 = ~x5 & (x2 ? ~n1973 : ~n1972);
  assign n1972 = (x0 | ~x1 | ~x3 | x4 | ~x6) & ((~x0 ^ ~x1) | (x3 ? (x4 | x6) : (~x4 | ~x6)));
  assign n1973 = (~x0 | x1 | ~x3 | ~x4 | ~x6) & (x0 | ((x4 | x6 | x1 | x3) & (~x1 | ((~x4 | x6) & (x3 | x4 | ~x6)))));
  assign n1974 = x0 ? (x1 | ~x2 | (~x4 ^ x7)) : (~x1 | x2 | (~x4 ^ ~x7));
  assign n1975 = ~n1976 & (n643 | (~x1 & n1979) | (x1 & n1980));
  assign n1976 = x5 & (x0 ? (~x1 & ~n1977) : ~n1978);
  assign n1977 = x2 ? (x4 | x6) : (~x4 | ~x6);
  assign n1978 = (x1 | ~x2 | x4 | ~x6) & (~x4 | ((~x1 | (x2 ? (~x3 | ~x6) : (x3 | x6))) & (x1 | ~x2 | ~x3 | x6)));
  assign n1979 = (~x0 | x4 | x5 | (x2 ^ ~x3)) & (~x4 | ((x0 | (x2 ? x5 : (x3 | ~x5))) & (~x0 | ~x2 | ~x3 | ~x5)));
  assign n1980 = (x0 | ((x2 | x3 | ~x4 | x5) & (~x2 | x4 | ~x5))) & (~x0 | x2 | x3 | ~x4 | ~x5);
  assign n1981 = ~n640 & (x0 ? ~n1983 : ~n1982);
  assign n1982 = (~x1 | ~x4 | ~x5 | (x2 ^ ~x3)) & (x4 | ((x3 | x5 | ~x1 | x2) & (x1 | (x2 ? (~x3 | x5) : ~x5))));
  assign n1983 = (~x1 | x2 | x3 | x4 | ~x5) & (x1 | ~x4 | x5 | (x2 & x3));
  assign n1984 = x1 & (x4 ? (~n1701 & n1988) : ~n1985);
  assign n1985 = (~n600 | ~n951) & (~n1986 | n1987);
  assign n1986 = ~x0 & ~x7;
  assign n1987 = (~x5 | ~x6 | x2 | ~x3) & (~x2 | x5 | (~x3 ^ ~x6));
  assign n1988 = x3 & ~x0 & x2;
  assign z073 = ~n2005 | ~n1999 | n1990 | n1996;
  assign n1990 = ~x0 & (n1991 | n1993 | n1995);
  assign n1991 = x5 & (x4 ? ~n1992 : (n1300 & n979));
  assign n1992 = (x1 | x2 | ~x3 | ~x6 | x7) & ((x2 ? (~x3 | ~x6) : (x3 | x6)) | (~x1 ^ x7));
  assign n1993 = ~n1994 & (n1203 | (~x3 & ~n1097));
  assign n1994 = x1 ? (x2 | ~x7) : (~x2 | x7);
  assign n1995 = n558 & n830;
  assign n1996 = ~n1198 & (n1997 | (n828 & ~n1543 & ~n1998));
  assign n1997 = x3 & ((x0 & ~x1 & x2 & ~x7) | (~x0 & (x1 ? (x2 ^ ~x7) : (~x2 & x7))));
  assign n1998 = x0 ^ ~x2;
  assign n1999 = (~n841 | n2002) & (~x1 | n2000) & (x1 | n2001);
  assign n2000 = (x0 | ~x2 | (x3 ? (x5 | x7) : (~x5 | ~x7))) & (~x0 | x2 | x3 | ~x5 | ~x7);
  assign n2001 = x0 ? ((~x2 | x3 | ~x5 | x7) & (x2 | ~x3 | x5 | ~x7)) : (~x3 | (x2 ? (~x5 ^ x7) : (x5 | x7)));
  assign n2002 = (~n2003 | ~n951) & (~n2004 | (x3 & x4));
  assign n2003 = x4 & x2 & x3;
  assign n2004 = (x5 ^ ~x6) & (~x2 ^ x7);
  assign n2005 = x3 ? n2007 : (~n2006 & (~n670 | ~n816));
  assign n2006 = ~n1543 & ((n1477 & n743) | (~x0 & ~n1934));
  assign n2007 = (~n1209 | ~n717) & (x2 | n2008);
  assign n2008 = (x0 | ~x1 | ~x4 | ~x5 | ~x7) & (~x0 | x7 | (x1 ? (x4 | x5) : (~x4 | ~x5)));
  assign z074 = n2028 | n2025 | n2010 | ~n2014;
  assign n2010 = ~n643 & (n2012 | ~n2013 | (~x1 & ~n2011));
  assign n2011 = (x0 | x4 | x5 | (~x2 ^ ~x3)) & (~x0 | ~x2 | ~x3 | ~x4 | ~x5);
  assign n2012 = x4 & ((~x2 & ~x3 & x0 & ~x1) | (~x0 & (x1 ? (~x2 & x3) : (x2 & ~x3))));
  assign n2013 = (~n1287 | ~n746) & (x4 | ~n743 | n1763);
  assign n2014 = ~n2016 & n2020 & (x0 ? n2015 : n2019);
  assign n2015 = (~x1 | x2 | x3 | ~x4 | x6) & (x1 | ((x4 | ~x6 | ~x2 | ~x3) & (x2 | (x3 ? (~x4 | x6) : (x4 | ~x6)))));
  assign n2016 = x2 & ((~n2017 & ~n2018) | (n626 & n946));
  assign n2017 = x3 ? (~x4 | x7) : (x4 | ~x7);
  assign n2018 = (x0 | ~x1 | ~x5 | x6) & (x5 | ~x6 | ~x0 | x1);
  assign n2019 = x1 ? ((~x2 | x3 | ~x4 | x6) & (x2 | ~x3 | x4 | ~x6)) : (~x4 | x6 | (~x2 ^ ~x3));
  assign n2020 = (~x5 | ~n2021 | n2022) & (n2023 | ~n2024);
  assign n2021 = x4 & ~x3 & ~x0 & ~x2;
  assign n2022 = x1 ? (x6 | x7) : (~x6 | ~x7);
  assign n2023 = x1 ? (~x2 ^ ~x3) : (x2 | ~x3);
  assign n2024 = x6 & x5 & ~x0 & x4;
  assign n2025 = ~x4 & ((n1269 & n2026) | (~x6 & ~n2027));
  assign n2026 = x6 & ~x3 & ~x5;
  assign n2027 = x0 ? (x5 | (x1 ? (x2 | ~x3) : (~x2 | x3))) : (x1 | ~x5 | (~x2 ^ ~x3));
  assign n2028 = ~n640 & (~n2029 | (~x5 & n566 & ~n2023));
  assign n2029 = ~n2030 & (~n1209 | ~n1311) & (~n1167 | n2023);
  assign n2030 = x4 & ~x3 & x2 & x0 & ~x1;
  assign z075 = ~n2041 | n2039 | n2032 | n2036;
  assign n2032 = ~x1 & (n2033 | (n1300 & ~n2035));
  assign n2033 = ~x6 & ((n600 & n670) | (x7 & ~n2034));
  assign n2034 = x0 ? (~x5 | (x2 ? (x3 | ~x4) : (~x3 | x4))) : (x5 | (x2 ? (~x3 | x4) : (~x3 ^ ~x4)));
  assign n2035 = (x0 | x2 | x3 | ~x4 | ~x5) & (~x2 | (~x3 ^ ~x4) | (~x0 ^ x5));
  assign n2036 = ~x5 & (x2 ? ~n2037 : ~n2038);
  assign n2037 = (~x0 | x1 | x3 | ~x4 | ~x7) & ((~x3 ^ ~x4) | (x0 ? (x1 | x7) : (~x1 | ~x7)));
  assign n2038 = (x0 | ~x1 | x3 | ~x4 | ~x7) & (~x0 | x4 | (x1 ? (~x3 ^ x7) : (~x3 | ~x7)));
  assign n2039 = x1 & ((n600 & n1725) | (n1986 & ~n2040));
  assign n2040 = (~x2 | ~x3 | ~x4 | ~x5 | ~x6) & ((x2 ^ ~x4) | (x3 ? (x5 | x6) : (~x5 | ~x6)));
  assign n2041 = ~n2042 & ~n2044 & ~n2046 & (x2 | n2045);
  assign n2042 = ~n1532 & ((n841 & n1903) | (~x0 & ~n2043));
  assign n2043 = x1 ? (~x3 | ~x7) : (x3 | x7);
  assign n2044 = x4 & n742 & (x1 ? (~x3 & ~x7) : (x3 ^ x7));
  assign n2045 = ((x1 ^ ~x7) | (x0 ? (x3 | ~x4) : (~x3 | x4))) & (x3 | x4 | (x0 ? (x1 | x7) : (~x1 | ~x7)));
  assign n2046 = n551 & ((~n1744 & ~n2048) | (n742 & n2047));
  assign n2047 = ~x7 & x3 & ~x4;
  assign n2048 = x0 ? (~x2 | ~x7) : (x2 | x7);
  assign z076 = n2062 | ~n2065 | (x1 ? ~n2050 : ~n2053);
  assign n2050 = ~n609 & (x0 | (~x2 & n2052) | (x2 & n2051));
  assign n2051 = x3 ? ((x6 | ~x7 | ~x4 | ~x5) & (x4 | (x5 ? (~x6 | x7) : (x6 | ~x7)))) : ((~x4 | x5 | ~x6 | x7) & (x4 | ~x5 | x6 | ~x7));
  assign n2052 = (~x5 | ((~x3 | ~x4 | ~x6 | x7) & (x3 | x6 | (~x4 ^ ~x7)))) & (~x3 | x5 | (x4 ? (x6 | ~x7) : (~x6 | x7)));
  assign n2053 = x3 ? (~n2054 & n2056) : (~n2059 & ~n2060);
  assign n2054 = ~n882 & ~n2055;
  assign n2055 = (~x6 | ~x7 | ~x4 | x5) & (x6 | x7 | x4 | ~x5);
  assign n2056 = (~n658 | ~n2057) & (~n1070 | ~n2058);
  assign n2057 = x4 & x0 & ~x2;
  assign n2058 = ~x4 & ~x0 & x2;
  assign n2059 = ~x0 & ((n658 & n859) | (n1070 & n1084));
  assign n2060 = n2061 & ((n1300 & n1156) | (~x2 & ~n1850));
  assign n2061 = x0 & ~x5;
  assign n2062 = ~n2063 & ~n2064;
  assign n2063 = x5 ? (~x6 | ~x7) : (x6 | x7);
  assign n2064 = (~x0 | ~x1 | x2 | x3 | x4) & (x1 | (x0 ? (x2 ? (x3 | ~x4) : (~x3 | x4)) : (x2 ? (~x3 ^ ~x4) : (x3 | ~x4))));
  assign n2065 = n2068 & (~n543 | n2066) & (x1 | n2067);
  assign n2066 = (~x2 | x4 | ~x6 | (~x3 ^ x5)) & (~x4 | ((x5 | x6 | ~x2 | x3) & (x2 | ~x5 | (x3 ^ ~x6))));
  assign n2067 = (x0 | x2 | ~x3 | ~x4 | ~x5) & (~x2 | ((x0 | x3 | ~x4 | x5) & (~x0 | x4 | (~x3 ^ x5))));
  assign n2068 = (n1010 | n2069) & (n1353 | n2070);
  assign n2069 = (x3 | x5 | ~x1 | x2) & (x1 | (x2 ? (~x3 | ~x5) : (~x3 ^ x5)));
  assign n2070 = (~x0 | x1 | x2 | x3 | x5) & (x0 | ~x1 | ~x3 | (~x2 ^ ~x5));
  assign z077 = ~n2080 | (x7 & (n2072 | n2078));
  assign n2072 = ~x0 & (n2073 | ~n2076 | (~n1480 & ~n1100));
  assign n2073 = ~n2075 & ~x6 & n2074;
  assign n2074 = x1 & x5;
  assign n2075 = x2 ? (~x3 | ~x4) : (x3 | x4);
  assign n2076 = (n1954 | n2077) & (~n704 | ~n558);
  assign n2077 = (x3 | ~x4 | ~x5 | x6) & (x5 | ~x6 | ~x3 | x4);
  assign n2078 = x0 & ((n576 & n1358) | (~x1 & ~n2079));
  assign n2079 = (~x2 | ~x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (x5 | ~x6 | x3 | x4) & (x2 | ~x4 | x6 | (x3 & ~x5));
  assign n2080 = ~n2081 & (x0 ? n2088 : n2084);
  assign n2081 = ~n1097 & (~n2083 | (x7 & ~n2082));
  assign n2082 = x1 ? ((x3 | x4 | ~x0 | x2) & (x0 | ~x3 | (~x2 ^ x4))) : (x0 ? (x2 ? (x3 | ~x4) : (~x3 | x4)) : (x2 ? (~x3 ^ ~x4) : (x3 | ~x4)));
  assign n2083 = x1 ? ((x2 | x3 | ~x4) & (x0 | ((x3 | x4) & (~x2 | ~x3 | ~x4)))) : ((~x3 | (x0 ? (~x2 ^ x4) : (x2 | x4))) & (x3 | ~x4 | x0 | ~x2));
  assign n2084 = x2 ? n2086 : (~n2087 & (n1100 | n2085));
  assign n2085 = x1 ^ x3;
  assign n2086 = x1 ? ((x3 | ~x4 | ~x5 | x6) & (~x3 | x4 | x5 | ~x6)) : ((~x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (x5 | ~x6 | x3 | x4));
  assign n2087 = ~x6 & x5 & x4 & ~x1 & x3;
  assign n2088 = x1 ? (~n704 | ~n1044) : (~n1623 & ~n2089);
  assign n2089 = ~x3 & (x4 ? (~x5 & x6) : (x5 & ~x6));
  assign z078 = ~n2096 | n2105 | ~n2107 | (~x1 & ~n2091);
  assign n2091 = x2 ? (x0 ? n740 : n2092) : n2093;
  assign n2092 = x3 ? ((x4 | ~x5 | ~x6 | x7) & (~x4 | x5 | x6 | ~x7) & ((~x6 ^ ~x7) | (~x4 ^ ~x5))) : (x4 ? (x5 ? (x6 | ~x7) : (~x6 | x7)) : (x5 ? (~x6 ^ ~x7) : (x6 | ~x7)));
  assign n2093 = (~n658 | ~n2094) & (x0 | n2095);
  assign n2094 = x4 & x0 & ~x3;
  assign n2095 = x3 ? (x4 ? (x5 ? (~x6 | x7) : (~x6 ^ ~x7)) : (x5 ? (x6 | ~x7) : (~x6 | x7))) : ((~x6 | ~x7 | ~x4 | ~x5) & ((~x4 ^ x6) | (~x5 ^ x7)));
  assign n2096 = ~n2098 & ~n2100 & n2102 & (n1532 | n2097);
  assign n2097 = (x0 | ~x1 | ~x3 | ~x5 | x6) & (~x6 | ((x3 | x5 | x0 | ~x1) & (~x0 | x1 | (~x3 ^ x5))));
  assign n2098 = ~n1097 & (x0 ? (~x1 & ~n2075) : (x1 & ~n2099));
  assign n2099 = x2 ? (x3 | ~x4) : (~x3 | x4);
  assign n2100 = ~n2101 & ~x6 & n841;
  assign n2101 = (x2 | ~x3 | x4 | ~x5) & (~x2 | x3 | (~x4 ^ ~x5));
  assign n2102 = (n1282 | n2103) & (n1701 | n2104);
  assign n2103 = (x2 | ~x3 | ~x0 | x1) & (~x1 | ((x2 | x3) & (x0 | ~x2 | ~x3)));
  assign n2104 = x0 ? (x1 | ((x3 | x4) & (~x2 | ~x3 | ~x4))) : (~x1 | (x2 ? (x3 | ~x4) : (~x3 | x4)));
  assign n2105 = n543 & (x2 ? (n828 & n813) : ~n2106);
  assign n2106 = (~x3 | ~x4 | ~x5 | ~x6 | ~x7) & (x3 | x4 | (x5 ? (x6 | ~x7) : (~x6 | x7)));
  assign n2107 = ~n2108 & (n643 | (n2111 & (~x4 | n2110)));
  assign n2108 = x1 & ((n600 & n728) | (~x5 & ~n2109));
  assign n2109 = (x0 | ~x2 | ~x3 | ~x4 | ~x6) & (~x0 | x2 | (x3 ? (x4 | x6) : (~x4 | ~x6)));
  assign n2110 = (x0 | ~x1 | ~x2 | ~x3 | ~x5) & (~x0 | x3 | (x1 ? (x2 | ~x5) : x5));
  assign n2111 = x2 ? (x4 | n2113) : ((~x4 | n2113) & (~x0 | x4 | ~n2112));
  assign n2112 = ~x5 & (x1 ^ x3);
  assign n2113 = (x0 | ~x1 | (~x3 ^ x5)) & (~x3 | ~x5 | ~x0 | x1);
  assign z079 = n2115 | n2119 | ~n2123 | (~n1116 & ~n2122);
  assign n2115 = ~x1 & (x2 ? ~n2116 : ~n2117);
  assign n2116 = (x0 | x3 | x4 | ~n951) & (~x4 | ~n978 | ~x0 | ~x3);
  assign n2117 = (x3 | n2118) & (~x4 | ~n978 | x0 | ~x3);
  assign n2118 = (x0 | x4 | x5 | ~x7) & (~x0 | ~x4 | ~x5 | x6);
  assign n2119 = ~n640 & (n1905 | n2121 | (~x3 & ~n2120));
  assign n2120 = x1 ? (x2 | (x5 ? ~x0 : x4)) : (x0 ? ((x4 | x5) & (~x2 | ~x4 | ~x5)) : (~x5 | (x2 & x4)));
  assign n2121 = n1188 & (x0 ? (x2 ? (x4 & ~x5) : (~x4 & x5)) : (x2 ? (x4 ^ ~x5) : (x4 & ~x5)));
  assign n2122 = (x1 | ((~x0 | (x4 ? ~x3 : ~x2)) & (~x2 | x3 | x4) & (x0 | ((x3 | ~x4) & (x2 | ~x3 | x4))))) & (~x1 | x2 | x3 | ~x4) & (x0 | ((~x2 | ~x3 | ~x4) & (~x1 | x3 | x4)));
  assign n2123 = ~n2125 & ~n2127 & (~n1017 | n2124);
  assign n2124 = (x0 | x3 | ~x5 | ~x6) & (~x0 | x5 | (x3 ? x7 : (x6 | ~x7)));
  assign n2125 = ~n2126 & (x0 ? ~x1 : x2);
  assign n2126 = (x3 | ~x4 | ~x5 | ~x6 | x7) & (~x3 | x4 | x5 | x6 | ~x7);
  assign n2127 = ~n2128 & ((~x1 & (~n1794 | (~x2 & ~n2129))) | (~x2 & ~n1794));
  assign n2128 = (x4 | ~x5 | ~x6 | x7) & (x6 | ~x7 | ~x4 | x5);
  assign n2129 = x0 ^ x3;
  assign z080 = n2131 | ~n2140 | ~n2146 | (~n1701 & ~n2139);
  assign n2131 = ~x0 & (n2136 | (x7 & (n2132 | ~n2134)));
  assign n2132 = ~x1 & (x2 ? ~n2133 : ~n928);
  assign n2133 = (x5 | x6 | ~x3 | x4) & (x3 | (x4 ? (x5 | ~x6) : (~x5 | x6)));
  assign n2134 = (~n559 | ~n2135) & (n1408 | n2069);
  assign n2135 = x3 & x1 & x2;
  assign n2136 = ~x7 & ((~n1097 & ~n2137) | (~x1 & ~n2138));
  assign n2137 = (x3 | x4 | ~x1 | x2) & (x1 | (x2 ? (x3 | ~x4) : (~x3 | x4)));
  assign n2138 = (x2 | ~x3 | ~x4 | ~x5 | x6) & (~x2 | x3 | x4 | x5 | ~x6) & ((~x2 ^ ~x3) | (x4 ? (x5 | ~x6) : (~x5 | x6)));
  assign n2139 = (~x0 | x1 | ~x2 | ~x3 | ~x4) & ((x0 ? (x1 | x3) : (~x1 | ~x3)) | (~x2 ^ x4));
  assign n2140 = ~n2141 & ~n2142 & n2143 & (n1036 | n2077);
  assign n2141 = ~n1097 & ~n2139;
  assign n2142 = ~n1138 & n681 & n743;
  assign n2143 = (~n588 | ~n2144) & (~n746 | ~n2145);
  assign n2144 = ~x3 & ~x2 & x0 & ~x1;
  assign n2145 = ~x6 & x5 & x3 & x4;
  assign n2146 = n2149 & (n643 | (n2148 & (n1134 | n2147)));
  assign n2147 = (x0 | ~x1 | ~x2 | x3) & (~x0 | x2 | (~x1 ^ x3));
  assign n2148 = (~n639 | ~n1209) & (n1934 | n1119);
  assign n2149 = (n740 | n1036) & (n2147 | (n1100 & n1282));
  assign z081 = n2151 | n2158 | ~n2163 | (~n1116 & ~n2162);
  assign n2151 = ~x2 & (n2156 | (x0 & (n2152 | n2154)));
  assign n2152 = ~x1 & ((n1392 & n2153) | (n774 & n951));
  assign n2153 = x5 & (~x6 ^ ~x7);
  assign n2154 = ~x5 & n1445 & (n2155 | n1903);
  assign n2155 = x7 & ~x3 & ~x6;
  assign n2156 = ~x0 & (x1 ? ~n2157 : ~n2126);
  assign n2157 = (~x3 | ~x4 | ~x5 | ~x6 | x7) & (x3 | x5 | (x4 ? (~x6 | x7) : (x6 | ~x7)));
  assign n2158 = ~n640 & ((~x1 & ~n2159) | ~n2161 | (x1 & ~n2160));
  assign n2159 = x4 ? (x2 ? (~x3 | x5) : ((x3 | x5) & (~x0 | ~x3 | ~x5))) : ((x0 | ~x3 | ~x5) & (~x2 | (~x3 ^ ~x5)));
  assign n2160 = (~x4 | ((x2 | x3 | ~x5) & (x0 | ~x3 | (~x2 ^ ~x5)))) & (x0 | ~x2 | x4 | (~x3 ^ x5));
  assign n2161 = (~x1 | x2 | x3 | x4) & (x1 | ((~x2 | x3 | ~x4) & (~x0 | x2 | ~x3 | x4)));
  assign n2162 = x3 ? ((~x2 & ~x4) ? (x0 | ~x1) : x1) : ((~x0 | (x1 ? (x2 | ~x4) : x4)) & (x1 | x2 | x4) & (x0 | ~x1 | ~x2 | ~x4));
  assign n2163 = ~n2164 & (~x2 | (~n2165 & (~n699 | ~n845)));
  assign n2164 = ~n2128 & (x3 ? ~n1957 : ~n1954);
  assign n2165 = ~x1 & ((n1392 & n978) | (x3 & ~n1113));
  assign z082 = ~n2173 | n2179 | (x3 ? ~n2182 : ~n2167);
  assign n2167 = x2 ? n2170 : (~n2168 & n2169);
  assign n2168 = n750 & (x0 ? (~x1 & n597) : (x1 & ~n1353));
  assign n2169 = n1282 & (~n529 | ~n951);
  assign n2170 = (x1 | n2172) & (x0 | ~x1 | n2171);
  assign n2171 = (x4 | ~x5 | ~x6 | x7) & (x6 | ~x7 | ~x4 | x5) & ((~x6 ^ ~x7) | (~x4 ^ ~x5));
  assign n2172 = x4 ? ((~x5 | ~x6 | ~x7) & (x0 | x6 | (~x5 ^ x7))) : ((x5 | x6 | x7) & (~x0 | ((x6 | x7) & (x5 | ~x6 | ~x7))));
  assign n2173 = x6 ? (~n2175 & (~x4 | n2174)) : n2178;
  assign n2174 = x2 ? (~x3 | ~x5 | (~x0 ^ x1)) : (x3 | x5);
  assign n2175 = n1145 & (n2177 | (x2 & ~n2176));
  assign n2176 = x0 ? (x3 ^ ~x5) : (x3 | x5);
  assign n2177 = x5 & x3 & ~x0 & ~x2;
  assign n2178 = (~x3 | x5 | n1350) & (~x5 | ((~n804 | n1327) & (x3 | n1350)));
  assign n2179 = ~n643 & ((~x3 & ~n2181) | (~x1 & n2180));
  assign n2180 = x3 & ((~x0 & ~x2 & x4 & ~x5) | (x0 & x2 & ~x4 & x5));
  assign n2181 = (x1 | ((x5 | ((x2 | x4) & (~x0 | ~x2 | ~x4))) & (x0 | ~x5 | (~x2 ^ x4)))) & (~x0 | x2 | ((x4 | x5) & (~x1 | ~x4 | ~x5)));
  assign n2182 = x1 ? (x0 | n2189) : (n2183 & n2186);
  assign n2183 = (n1701 | n2184) & (n1116 | n2185);
  assign n2184 = x0 ? (~x2 | ~x4) : (x2 | x4);
  assign n2185 = x0 ? (x2 | ~x4) : (~x2 | x4);
  assign n2186 = (n640 | n2187) & (n697 | n2188);
  assign n2187 = (x0 | ~x2 | ~x4 | x5) & (x4 | ~x5 | ~x0 | x2);
  assign n2188 = (x5 | x6 | ~x0 | x4) & (~x5 | ~x6 | x0 | ~x4);
  assign n2189 = ((x2 ? (~x4 | x5) : (x4 | ~x5)) | (~x6 ^ ~x7)) & (x2 | x4 | x5 | x6 | ~x7) & ((~x2 ^ x4) | (x5 ? (x6 | ~x7) : (~x6 | x7)));
  assign z083 = ~n2206 | (x2 ? (~n2197 | ~n2199) : ~n2191);
  assign n2191 = x0 ? n2194 : (x3 ? n2192 : n2193);
  assign n2192 = x6 ? (((~x1 ^ ~x4) | (~x5 ^ x7)) & (x1 | ~x4 | ~x5 | ~x7) & (x5 | x7 | ~x1 | x4)) : (x4 ? (x5 | x7) : (~x5 | ~x7));
  assign n2193 = (~x1 & (x4 ^ (x6 & ~x7))) | (x5 & (x6 ^ x7)) | (~x5 & (x6 ^ ~x7)) | (x6 & x7 & x1 & ~x4);
  assign n2194 = (x3 | n2195) & (x1 | ~x3 | n2196);
  assign n2195 = x6 ? ((x4 | ~x5 | ~x7) & (~x4 | x5 | x7) & (x1 | (x7 ? ~x5 : ~x4))) : ((x5 | x7 | ~x1 | x4) & ((~x1 ^ ~x4) | (~x5 ^ x7)));
  assign n2196 = (~x6 | ~x7 | ~x4 | x5) & (x6 | x7 | x4 | ~x5) & ((~x4 ^ ~x5) | (~x6 ^ x7));
  assign n2197 = (~n699 | ~n845) & (n643 | n2198);
  assign n2198 = (~x0 | x1 | ~x3 | ~x4 | ~x5) & (x0 | ((x4 | x5 | x1 | x3) & (~x1 | (x3 ? (x4 | ~x5) : (~x4 | x5)))));
  assign n2199 = (n1566 | n2200) & (x1 | (~n2201 & n2203));
  assign n2200 = x0 ? (x1 | (x4 ? (~x6 ^ ~x7) : (~x6 | x7))) : (x1 ? (x4 ? (x6 | x7) : (~x6 | ~x7)) : (x6 | (~x4 ^ ~x7)));
  assign n2201 = ~x0 & (n2202 | (n1392 & n942));
  assign n2202 = x3 & ((x6 & x7 & ~x4 & ~x5) | (~x6 & ~x7 & x4 & x5));
  assign n2203 = (~n943 | ~n2204) & (n1218 | n2205);
  assign n2204 = ~x4 & x0 & x3;
  assign n2205 = (x5 | x6 | ~x0 | x3) & (~x5 | ~x6 | x0 | ~x3);
  assign n2206 = x2 ? n2214 : (n2207 & n2211);
  assign n2207 = (~n727 | ~n2209) & (n2208 | n2210);
  assign n2208 = x1 ^ ~x4;
  assign n2209 = ~x7 & ~x4 & ~x5;
  assign n2210 = (x0 | x3 | ~x5 | ~x7) & (x5 | x7 | ~x0 | ~x3);
  assign n2211 = x5 ? ((x7 | n2213) & (~x0 | ~x7 | n2212)) : (~x7 | n2213);
  assign n2212 = x1 ? (x3 | ~x4) : (~x3 | x4);
  assign n2213 = (x0 | x1 | ~x3 | ~x4) & (x3 | x4 | ~x0 | ~x1);
  assign n2214 = x3 ? (~n543 | n2216) : n2215;
  assign n2215 = (~x0 | x1 | x4 | x5 | ~x7) & (x0 | ~x5 | (x1 ? (~x4 ^ ~x7) : (x4 | ~x7)));
  assign n2216 = x4 ? (x5 ^ ~x7) : (x5 | x7);
  assign z084 = n2235 | n2232 | ~n2225 | n2218 | n2221;
  assign n2218 = ~x5 & (x1 ? ~n2219 : ~n2220);
  assign n2219 = (x0 | (x2 ? (x4 | x6) : (~x4 | ~x6))) & (x2 | ((x3 | ~x4 | ~x6) & (x4 | x6 | ~x0 | ~x3)));
  assign n2220 = (x0 | ~x2 | x4 | ~x6) & (~x3 | ~x4 | (x0 ? (~x2 ^ ~x6) : (~x2 | x6)));
  assign n2221 = ~x3 & (x5 ? ~n2222 : (n1181 & ~n2224));
  assign n2222 = (~x2 | ~x6 | n2223) & (x6 | ((~n1145 | n2048) & (x2 | n2223)));
  assign n2223 = (~x0 | x1 | ~x4 | x7) & (x0 | ~x1 | x4 | ~x7);
  assign n2224 = (x1 | ~x4 | x6 | ~x7) & (~x1 | x7 | (x4 ^ ~x6));
  assign n2225 = ~n2226 & (~x3 | n2230);
  assign n2226 = ~n1218 & ((n793 & ~n2228) | (~n2227 & ~n2229));
  assign n2227 = x2 ^ ~x3;
  assign n2228 = x1 ? (~x5 | x6) : (~x5 ^ ~x6);
  assign n2229 = (x5 | ~x6 | ~x0 | x1) & (x0 | (x1 ? (~x5 | x6) : (~x5 ^ ~x6)));
  assign n2230 = (~n1209 | ~n830) & (x0 | n682 | n2231);
  assign n2231 = (~x2 | (x4 ? (x5 | ~x7) : (~x5 | x7))) & (x2 | x4 | x5 | ~x7);
  assign n2232 = x5 & ((n543 & n2234) | (~x1 & ~n2233));
  assign n2233 = (~x3 | ((x0 | ~x2 | ~x4 | ~x6) & (~x0 | (x2 ? (x4 | x6) : (~x4 | ~x6))))) & (x0 | x2 | ((~x4 | x6) & (x3 | x4 | ~x6)));
  assign n2234 = x2 & x3 & (x4 ^ x6);
  assign n2235 = ~n671 & (x0 ? ~n2236 : ~n2237);
  assign n2236 = (x1 | ~x2 | ((x5 | x6) & (~x3 | ~x5 | ~x6))) & (x2 | ((~x5 | x6 | x1 | ~x3) & (x3 | (x1 ? (~x5 ^ ~x6) : (x5 | ~x6)))));
  assign n2237 = (x1 | ~x2 | ~x5 | x6) & (~x6 | ((x3 | x5 | x1 | x2) & (~x1 | (~x2 ^ x5))));
  assign z085 = ~n2245 | n2255 | (x3 ? ~n2257 : ~n2239);
  assign n2239 = x7 ? (~n2244 & (x2 | n2243)) : n2240;
  assign n2240 = x2 ? n2241 : n2242;
  assign n2241 = (x0 | x1 | ~x4 | x5 | ~x6) & ((x0 ? (x1 | x4) : (~x1 | ~x4)) | (~x5 ^ ~x6));
  assign n2242 = (~x0 | ~x1 | ~x4 | x5 | ~x6) & (x0 | x4 | (x1 ? (x5 | x6) : (~x5 | ~x6)));
  assign n2243 = (x0 | ~x1 | ~x4 | x5 | x6) & (~x5 | ((x0 | ~x1 | ~x4 | ~x6) & (~x0 | x1 | (~x4 ^ x6))));
  assign n2244 = n570 & ((n525 & n1364) | (n904 & n1167));
  assign n2245 = n2253 & ~n2251 & ~n2246 & ~n2249;
  assign n2246 = ~n1198 & (x1 ? ~n2248 : ~n2247);
  assign n2247 = (x0 | ~x2 | x3 | x4 | x7) & (~x3 | (x0 ? (x2 ? (~x4 | x7) : (x4 | ~x7)) : (~x4 | (~x2 ^ ~x7))));
  assign n2248 = (x0 | ~x2 | x3 | ~x7) & (x2 | x7 | (x0 ? (x3 | x4) : (~x3 ^ x4)));
  assign n2249 = ~x0 & ((n918 & ~n1150) | (~x7 & ~n2250));
  assign n2250 = (~x1 | ~x2 | (x3 ? (~x4 | ~x5) : (x4 | x5))) & (x2 | ((~x1 | ~x3 | ~x4 | x5) & (x1 | ~x5 | (~x3 ^ x4))));
  assign n2251 = ~n1008 & ((n1141 & n746) | (~x2 & ~n2252));
  assign n2252 = (x0 | ~x1 | x3 | x4 | ~x6) & (~x0 | x1 | ~x4 | (~x3 ^ ~x6));
  assign n2253 = (~x7 | n2254) & (x7 | ~n1269 | ~x3 | x5);
  assign n2254 = (x0 | ~x1 | x2 | ~x3 | ~x5) & (x3 | (x0 ? (x1 ? (x2 | ~x5) : (~x2 | x5)) : (x1 | (~x2 ^ ~x5))));
  assign n2255 = x0 & ((n979 & n2209) | (~x1 & ~n2256));
  assign n2256 = (x2 | x3 | x4 | x5 | ~x7) & (x7 | ((x4 | x5 | x2 | ~x3) & (~x5 | (x2 ? (x3 ^ ~x4) : (x3 | x4)))));
  assign n2257 = n2261 & (x1 | (~n2258 & ~n2260));
  assign n2258 = ~x7 & (x0 ? (~x2 & ~n2259) : (x2 & n559));
  assign n2259 = x4 ? (x5 | x6) : (~x5 | ~x6);
  assign n2260 = n943 & n2058;
  assign n2261 = (~n813 | ~n746) & (~n619 | n1097 | n882);
  assign z086 = ~n2279 | (x3 ? ~n2263 : (n2271 | ~n2274));
  assign n2263 = n2269 & (x1 | (~n2265 & (~n2264 | ~n2268)));
  assign n2264 = ~x7 & (x2 ^ ~x5);
  assign n2265 = ~n640 & (n2266 | (~x4 & (~n882 | ~n2267)));
  assign n2266 = ~x5 & x4 & ~x0 & x2;
  assign n2267 = x0 ? (x2 | x5) : (~x2 | ~x5);
  assign n2268 = ~x6 & ~x0 & x4;
  assign n2269 = (~n746 | ~n830) & (n643 | n2270);
  assign n2270 = (x2 | ((x0 | ~x1 | x4) & (~x4 | ~x5 | ~x0 | x1))) & (x0 | ~x1 | ((x4 | ~x5) & (~x2 | ~x4 | x5)));
  assign n2271 = x0 & ((~x6 & ~n2272) | (~x1 & n2273));
  assign n2272 = (~x1 | x2 | ~x4 | x5 | ~x7) & (x1 | x4 | ~x5 | (~x2 ^ ~x7));
  assign n2273 = x2 & x6 & (x4 ? (x5 & x7) : (~x5 & ~x7));
  assign n2274 = n2277 & (x6 ? (x7 ? n2276 : n2275) : (x7 ? n2275 : n2276));
  assign n2275 = (x0 | x1 | ~x2 | ~x4 | x5) & (x4 | (x0 ? (~x1 | x2) : (x1 | (x2 & ~x5))));
  assign n2276 = (x0 | ~x1 | ~x2 | x4) & (x2 | ~x4 | ~x0 | x1);
  assign n2277 = (~n830 | ~n1269) & (n538 | n2278);
  assign n2278 = (x0 | ~x1 | ~x4 | x7) & (x4 | ~x7 | ~x0 | x1);
  assign n2279 = x6 ? (~n2280 & n2281) : (~n2284 & n2285);
  assign n2280 = n1188 & (x0 ? (~x2 & ~n714) : (x2 & n1121));
  assign n2281 = ~n2282 & ~n2283 & (~n1268 | ~n733);
  assign n2282 = x4 & x3 & x2 & x0 & ~x1;
  assign n2283 = ~x0 & ((x3 & x4 & ~x1 & ~x2) | (x1 & ~x3 & (x2 ^ ~x4)));
  assign n2284 = ~n2085 & ((~x4 & ~x5 & x0 & ~x2) | (~x0 & x4 & (~x2 | x5)));
  assign n2285 = (~n1716 | ~n1269) & (~x4 | ~n622 | n2286);
  assign n2286 = x1 ? (x2 | ~x5) : ~x2;
  assign z087 = ~n2293 | ~n2304 | (x4 ? ~n2299 : ~n2288);
  assign n2288 = (x0 | n2289) & (~n1857 | ~n1451 | ~x0 | ~n632);
  assign n2289 = x7 ? (n2085 | n2291) : (n2290 | ~n2292);
  assign n2290 = x1 ^ ~x5;
  assign n2291 = x2 ? (x5 | ~x6) : (~x5 | x6);
  assign n2292 = ~x6 & x2 & x3;
  assign n2293 = ~n2295 & (n643 | (~n2294 & (~n622 | n2298)));
  assign n2294 = n731 & n1269;
  assign n2295 = x2 & ((n2296 & n699) | (~x1 & ~n2297));
  assign n2296 = x7 & ~x4 & ~x5;
  assign n2297 = (~x4 | ((~x0 | x3 | ~x5 | x7) & (x0 | x5 | ~x7))) & (x0 | x4 | ((x5 | x7) & (~x3 | ~x5 | ~x7)));
  assign n2298 = (~x1 | x2 | ~x4 | x5) & (x1 | ~x2 | x4 | ~x5);
  assign n2299 = ~n2300 & (~n1310 | n2303);
  assign n2300 = x5 & ((n1283 & n2302) | (n841 & ~n2301));
  assign n2301 = (~x6 | ~x7 | ~x2 | x3) & (x6 | x7 | x2 | ~x3);
  assign n2302 = ~x3 & (x6 ^ ~x7);
  assign n2303 = (x1 | x2 | ~x3 | ~x6 | x7) & (~x1 | ~x2 | (x3 ? (x6 | ~x7) : (~x6 | x7)));
  assign n2304 = ~n2306 & (n671 | n2305);
  assign n2305 = x0 ? ((~x1 | x2 | x3 | ~x5) & (x1 | ((~x3 | x5) & (~x2 | (~x3 & x5))))) : ((~x1 | (x2 ? ~x5 : (~x3 | x5))) & (~x2 | x3 | ~x5) & (x1 | x2 | (~x3 ^ ~x5)));
  assign n2306 = ~x2 & (x0 ? ~n2308 : ~n2307);
  assign n2307 = x1 ? (x7 | (x3 ^ (x4 & x5))) : ((x3 | ~x4 | ~x5 | x7) & (~x3 | x4 | x5 | ~x7));
  assign n2308 = (x4 | ((x1 | ~x3 | ~x5 | x7) & (x5 | (x1 ? (x3 ^ ~x7) : (x3 | x7))))) & (x1 | ~x7 | ((x3 | (~x4 & ~x5)) & (~x4 | ~x5)));
  assign z088 = n2310 | n2319 | ~n2324 | (~x0 & ~n2323);
  assign n2310 = ~x3 & (n2311 | (x2 & (n2314 | n2318)));
  assign n2311 = ~x2 & (x0 ? ~n2312 : ~n2313);
  assign n2312 = (~x1 | x4 | x5 | x6 | ~x7) & (~x4 | ((~x5 | ~x6 | x7) & (x1 | x6 | (~x5 ^ ~x7))));
  assign n2313 = (~x1 | ~x4 | x5 | x6 | x7) & (x4 | ((~x5 | ~x6 | ~x7) & (x1 | x5 | (~x6 ^ x7))));
  assign n2314 = n2315 & (x0 ? n2316 : n2317);
  assign n2315 = ~x1 & x6;
  assign n2316 = x4 & (x5 ^ ~x7);
  assign n2317 = ~x4 & (~x5 ^ ~x7);
  assign n2318 = n962 & x4 & n543;
  assign n2319 = x3 & ((n527 & ~n2321) | (n2320 & ~n2322));
  assign n2320 = x6 & ~x0 & x1;
  assign n2321 = (x0 | x4 | ~x5 | (~x2 ^ ~x7)) & (~x4 | (x2 ^ ~x7) | (x0 ^ x5));
  assign n2322 = (~x2 | ~x4 | x5 | ~x7) & (x2 | (x4 ? (x5 | x7) : (~x5 | ~x7)));
  assign n2323 = (~x2 | ((~x4 | ~x5 | x1 | x3) & (~x1 | (x3 ? (~x4 | ~x5) : (x4 | x5))))) & (x1 | x2 | x5 | (~x3 ^ x4));
  assign n2324 = ~n2326 & ~n2328 & ~n2331 & (~n543 | n2325);
  assign n2325 = (x3 | ~x4 | ~x6 | (x2 ^ ~x5)) & (x2 | x5 | x6 | (~x3 & x4));
  assign n2326 = ~x1 & ((n559 & n594) | (x2 & ~n2327));
  assign n2327 = (x0 | ~x3 | ~x5 | ~x6) & (x3 | ((x0 | x4 | ~x5 | x6) & (~x0 | ((x5 | x6) & (x4 | ~x5 | ~x6)))));
  assign n2328 = ~n1198 & (n2330 | (x1 & (n600 | n2329)));
  assign n2329 = ~x4 & x3 & ~x0 & x2;
  assign n2330 = x4 & x3 & ~x2 & ~x0 & ~x1;
  assign n2331 = n841 & (x2 ? (x3 & ~x5) : n2332);
  assign n2332 = ~x4 & x5;
  assign z089 = ~n2348 | n2346 | n2344 | n2334 | n2340;
  assign n2334 = x4 & (n2338 | (~x1 & (n2335 | n2336)));
  assign n2335 = ~x0 & ((n596 & n813) | (x3 & ~n1647));
  assign n2336 = n2337 & ((n757 & n1044) | (x2 & ~n1558));
  assign n2337 = x0 & ~x6;
  assign n2338 = x1 & ((n530 & n600) | (n1310 & ~n2339));
  assign n2339 = x3 ? (~x6 | ~x7) : (x2 ? (~x6 | x7) : (x6 | ~x7));
  assign n2340 = ~n2341 & ((~n1176 & n2343) | (~x2 & ~n2342));
  assign n2341 = x0 ^ ~x6;
  assign n2342 = (~x4 | ((x1 | ~x3 | ~x7) & (~x1 | x3 | ~x5 | x7))) & (x1 | ~x3 | x5 | x7) & (x4 | (x1 & x5) | (x3 ^ ~x7));
  assign n2343 = x3 & ~x1 & x2;
  assign n2344 = n1167 & (x5 ? ~n2345 : (n569 & n576));
  assign n2345 = (~x1 | ~x2 | x3 | ~x6 | x7) & (x6 | ((x2 | x3 | x7) & (x1 | (~x3 ^ ~x7))));
  assign n2346 = ~x4 & ((n1792 & n733) | (~x1 & ~n2347));
  assign n2347 = (x0 | ~x2 | x3 | ~x6 | ~x7) & (~x0 | x2 | x6 | (~x3 ^ ~x7));
  assign n2348 = n2358 & ~n2356 & ~n2354 & ~n2349 & ~n2351;
  assign n2349 = ~x3 & ~n2350;
  assign n2350 = (x0 | x1 | x2 | ~x4 | x6) & (x4 | ((x0 | ~x1 | ~x2 | x6) & (~x0 | ~x6 | (x1 ^ ~x2))));
  assign n2351 = ~n765 & ((n733 & n2352) | (n841 & ~n2353));
  assign n2352 = x6 & ~x3 & x4;
  assign n2353 = (x2 | x3 | ~x4 | ~x6) & (x4 | x6 | ~x2 | ~x3);
  assign n2354 = n1392 & ~n2355;
  assign n2355 = (~x0 | ~x1 | x2 | x5 | ~x6) & (x0 | ~x2 | ~x5 | (~x1 ^ ~x6));
  assign n2356 = x4 & ~n2357 & ((x3 & ~x7) | (x2 & ~x3 & x7));
  assign n2357 = x0 ? (x1 | ~x6) : (~x1 | x6);
  assign n2358 = ~x3 | ((~n626 | ~n696) & (~n2359 | ~n746));
  assign n2359 = ~x4 & x6;
  assign z090 = n2361 | ~n2366 | ~n2375 | (n619 & ~n2365);
  assign n2361 = ~x5 & (n2362 | (n689 & ~n2364));
  assign n2362 = x3 & ((n837 & n1395) | (~x1 & ~n2363));
  assign n2363 = x0 ? (x7 | ((~x4 | x6) & (~x2 | x4 | ~x6))) : (~x7 | ((x4 | ~x6) & (x2 | ~x4 | x6)));
  assign n2364 = (x0 | x2 | ~x4 | ~x6 | x7) & (~x2 | ((x6 | x7 | x0 | x4) & ((~x4 ^ x6) | (~x0 ^ x7))));
  assign n2365 = (x0 | ~x2 | x3 | x4 | ~x5) & (x5 | ((x3 | x4 | x0 | x2) & (~x0 | ~x4 | (x2 ^ ~x3))));
  assign n2366 = ~n2368 & ~n2370 & n2372 & (x1 | n2367);
  assign n2367 = (~x0 | x2 | x4 | x5 | x7) & (x0 | ~x5 | ((~x4 | x7) & (x2 | x4 | ~x7)));
  assign n2368 = ~n765 & (n2369 | (n1167 & (n632 | n1439)));
  assign n2369 = x4 & ~x3 & ~x2 & x0 & x1;
  assign n2370 = ~n1218 & ((x0 & n551) | (n543 & n2371));
  assign n2371 = x2 & ~x5;
  assign n2372 = (n2373 | n2374) & (~n635 | ~n733);
  assign n2373 = x0 ? (x2 | x3) : (~x2 | ~x3);
  assign n2374 = (~x1 | x4 | ~x5 | x7) & (x1 | ~x4 | x5 | ~x7);
  assign n2375 = (n1353 | n2376) & (~n1411 | n2378);
  assign n2376 = (~x5 | x7 | ~n543 | n2227) & (x5 | n2377);
  assign n2377 = (~x0 | ~x7 | (x1 ? (x2 | x3) : (~x2 | ~x3))) & (x0 | x1 | x2 | ~x3 | x7);
  assign n2378 = (x2 | x3 | ~x4 | ~x6 | x7) & (~x7 | ((~x3 | ~x4 | x6) & (~x2 | (~x4 ^ x6))));
  assign z091 = n2380 | n2394 | (x2 ? ~n2390 : ~n2386);
  assign n2380 = ~x1 & (n2381 | (~x0 & (n2383 | n2384)));
  assign n2381 = x0 & (x2 ? (n828 & n943) : ~n2382);
  assign n2382 = (x3 | x4 | x5 | ~x6 | ~x7) & (~x3 | x6 | x7 | (x4 ^ ~x5));
  assign n2383 = n865 & (n1216 | (x3 & n886));
  assign n2384 = n813 & n2385;
  assign n2385 = x4 & ~x2 & ~x3;
  assign n2386 = n2389 & (x6 | n2387) & (~n922 | ~n2388);
  assign n2387 = (~x0 | x1 | ~x3 | ~x5 | ~x7) & (x0 | ((~x5 | ~x7 | x1 | x3) & (~x1 | ((x5 | ~x7) & (~x3 | ~x5 | x7)))));
  assign n2388 = ~x3 & x6 & (x5 ^ ~x7);
  assign n2389 = (~x0 | x3 | (x1 ? (x5 | x6) : ~x5)) & (x1 | ~x5 | ~x6) & (x0 | x5 | (x1 ? ~x6 : (~x3 | x6)));
  assign n2390 = ~n2391 & ~n2392 & ~n2393 & (~n813 | ~n661);
  assign n2391 = n1686 & ((~x1 & ~x3 & x5 & x7) | (x3 & (x1 ? (x5 ^ x7) : (~x5 & ~x7))));
  assign n2392 = ~x0 & x1 & ((x5 & ~x6) | (~x3 & ~x5 & x6));
  assign n2393 = ~x1 & ((x0 & x5 & x6) | (~x5 & ~x6 & (~x0 | x3)));
  assign n2394 = n632 & ((n942 & n2204) | (~x6 & ~n2395));
  assign n2395 = (~x3 | ((~x5 | ~x7 | x0 | ~x4) & (~x0 | x4 | x5))) & (x0 | x3 | x7 | (~x4 ^ ~x5));
  assign z092 = ~n2410 | ~n2404 | n2397 | ~n2401;
  assign n2397 = ~n640 & (n2398 | n2399 | (n1181 & ~n2400));
  assign n2398 = ~x1 & ((~x3 & x4 & ~x0 & ~x2) | (x0 & (x2 ? (~x3 & ~x4) : (x3 & x4))));
  assign n2399 = ~x0 & x1 & ~x2 & (x3 ^ x4);
  assign n2400 = (x1 | x3 | x4 | ~x5) & (~x1 | ~x3 | ~x4 | x5);
  assign n2401 = ~n2403 & (~n1270 | ~n2402) & (~n733 | ~n2145);
  assign n2402 = ~x7 & ~x6 & x4 & ~x5;
  assign n2403 = ~x6 & ((~x0 & (x1 ? (x2 & ~x3) : (~x2 & x3))) | (x2 & x3 & x0 & ~x1));
  assign n2404 = ~n2405 & (x4 | (~n2407 & (~n746 | ~n2409)));
  assign n2405 = x6 & ~n2406;
  assign n2406 = (~x0 | x1 | x2 | x3 | ~x4) & (x0 | ((x1 | ~x2 | ~x3 | ~x4) & (~x1 | x2 | x3 | x4)));
  assign n2407 = n1300 & n804 & (n1875 | n2408);
  assign n2408 = ~x5 & ~x0 & ~x3;
  assign n2409 = ~x7 & ~x6 & x3 & ~x5;
  assign n2410 = ~n2413 & (n643 | (n2412 & (x4 | n2411)));
  assign n2411 = (x0 | x1 | ~x2 | x3 | ~x5) & (~x0 | ~x1 | x2 | ~x3 | x5);
  assign n2412 = (x0 | x1 | ~x2 | x3 | ~x4) & ((~x1 & x4) | (x0 ? (x2 | x3) : (~x2 | ~x3)));
  assign n2413 = ~x1 & (x0 ? ~n2414 : (n596 & n696));
  assign n2414 = (x2 | ~x3 | x4 | x5 | ~x6) & (~x2 | x3 | ~x4 | ~x5 | x6);
  assign z093 = n2416 | ~n2418 | (x2 ? ~n2426 : ~n2429);
  assign n2416 = x0 & ((n979 & n2209) | (~x1 & ~n2417));
  assign n2417 = (x2 | x3 | x4 | x5 | x7) & (~x7 | ((~x2 | ~x4 | (~x3 ^ x5)) & (x4 | x5 | x2 | ~x3)));
  assign n2418 = n2423 & (x1 | n2419) & (x0 | n2420);
  assign n2419 = x0 ? (x2 ? (x4 | (~x3 ^ ~x7)) : (~x4 | (~x3 ^ x7))) : ((x3 | ~x4 | x7) & (~x2 | ~x3 | (~x4 ^ ~x7)));
  assign n2420 = (~x1 | ~x3 | n2421) & (x1 | x3 | x4 | n2422);
  assign n2421 = (~x2 | x4 | ~x5 | x7) & (x2 | ~x4 | (~x5 ^ ~x7));
  assign n2422 = (~x5 | x7) & (~x2 | x5 | ~x7);
  assign n2423 = n2425 & (~n543 | n2424);
  assign n2424 = (x2 | x3 | x4 | ~x7) & (x7 | (x2 ? (~x3 | ~x4) : (x3 ^ ~x4)));
  assign n2425 = (~x0 | ~x1 | x2 | x3 | x7) & (x0 | ~x7 | (x1 ? (~x2 | x3) : (x2 | ~x3)));
  assign n2426 = (~n712 | ~n1621) & (x5 | (~n2427 & ~n2428));
  assign n2427 = n772 & ((n825 & n1857) | (x0 & n2302));
  assign n2428 = ~n643 & n543 & x3 & ~x4;
  assign n2429 = ~n2432 & (x7 | (~n2430 & (~n1358 | ~n866)));
  assign n2430 = n1145 & ((n1723 & n653) | (x0 & n2431));
  assign n2431 = x5 & (~x3 ^ x6);
  assign n2432 = n601 & n661;
  assign z094 = ~n2442 | (x1 ? ~n2439 : (n2434 | n2437));
  assign n2434 = ~x6 & ((n635 & n2435) | (~x2 & ~n2436));
  assign n2435 = x3 & ~x0 & x2;
  assign n2436 = (x0 | x3 | x4 | x5 | ~x7) & (~x5 | ((~x0 | (x3 ? (x4 | ~x7) : (~x4 | x7))) & (x0 | x3 | x4 | x7)));
  assign n2437 = n1364 & n859 & (x0 ? n2438 : n683);
  assign n2438 = x3 & x7;
  assign n2439 = ~n2440 & (~n600 | ~n2402);
  assign n2440 = ~x0 & (x2 ? (n828 & n978) : ~n2441);
  assign n2441 = (x4 | x5 | ~x6 | x7) & (~x3 | ~x4 | ~x5 | x6 | ~x7);
  assign n2442 = ~n2444 & (x2 ? (n2443 & n2448) : n2447);
  assign n2443 = (x0 | ~x1 | (x3 ? (~x4 ^ x5) : (x4 | x5))) & (x1 | (x0 ? (x3 ? (x4 | x5) : (~x4 | ~x5)) : (x3 ? (~x4 | ~x5) : (~x4 ^ x5))));
  assign n2444 = ~x2 & ((~x4 & ~n2445) | (~n623 & n2446));
  assign n2445 = (~x5 | ~x6 | ~x0 | x1) & (x0 | x5 | (x1 ? x6 : (x3 | ~x6)));
  assign n2446 = x4 & ~x0 & x3;
  assign n2447 = x0 ? (x1 ? (x3 | x4) : (~x4 | (~x3 & x5))) : (x1 ? (x3 | ~x4) : (~x3 | x4));
  assign n2448 = (~n592 | ~n661) & (n975 | ~n2449);
  assign n2449 = ~x0 & (~x1 ^ ~x4);
  assign z095 = n2451 | ~n2456 | ~n2461 | (~x2 & ~n2455);
  assign n2451 = ~x5 & (n2452 | (n1029 & n1769 & n1269));
  assign n2452 = ~x2 & ((x6 & ~n2453) | (n1285 & ~n2454));
  assign n2453 = (x0 | ~x1 | x4 | ~x7) & (x1 | ~x4 | x7 | (~x0 & x3));
  assign n2454 = x1 ? (~x4 | ~x7) : (x4 | x7);
  assign n2455 = (~x0 | ~x1 | x3 | x4 | x5) & (x0 | ((~x1 | (x3 ? (x4 | ~x5) : (~x4 | x5))) & (x1 | ~x3 | x4 | x5)));
  assign n2456 = n2458 & (n1198 | (~n932 & (~x4 | n2457)));
  assign n2457 = x0 ? (x3 | (x1 ^ ~x2)) : (x1 | ~x3);
  assign n2458 = ~x2 | (n2459 & (x5 | x6 | n2460));
  assign n2459 = (x0 | x1 | x4 | (~x3 ^ x5)) & ((~x3 ^ ~x5) | (x0 ? (x1 | x4) : (~x1 | ~x4)));
  assign n2460 = (x0 | x3 | (~x1 ^ x4)) & (~x3 | ~x4 | ~x0 | x1);
  assign n2461 = ~n2462 & (~x5 | (~n2465 & (~n543 | n2469)));
  assign n2462 = ~x2 & (x5 ? ~n2464 : (n772 & n2463));
  assign n2463 = ~x6 & (x0 | ~x3);
  assign n2464 = (x0 | ~x1 | x3 | x4 | x6) & (~x6 | ((~x3 | ~x4 | x0 | ~x1) & (x1 | ((x3 | x4) & (~x0 | (x3 & x4))))));
  assign n2465 = ~x1 & ((~n2466 & n2467) | (x7 & ~n2468));
  assign n2466 = x0 ? (~x2 | x3) : (x2 | ~x3);
  assign n2467 = ~x7 & (x4 ^ ~x6);
  assign n2468 = (~x0 | x2 | x3 | ~x4 | x6) & ((x2 ? (~x4 | ~x6) : (x4 | x6)) | (x0 ^ x3));
  assign n2469 = (x4 | ~x6 | (x2 ? (x3 ^ ~x7) : (x3 | x7))) & (x2 | ~x4 | x6 | (~x3 ^ ~x7));
  assign z096 = n2471 | n2478 | ~n2487 | (~n1408 & ~n2482);
  assign n2471 = ~n1353 & (n2473 | ~n2474 | (~x0 & ~n2472));
  assign n2472 = (x1 | x2 | ~x3 | x5 | x7) & (~x5 | ((x1 | x2 | ~x3 | ~x7) & (x7 | (x1 ? (x2 ^ ~x3) : (~x2 | ~x3)))));
  assign n2473 = ~x3 & (x1 ? (~x2 & (x5 | ~x7)) : ((~x5 & x7) | (x2 & (~x5 | x7))));
  assign n2474 = (~n1209 | ~n2476) & (~n1188 | (~n2475 & ~n2477));
  assign n2475 = x2 & (x5 ^ ~x7);
  assign n2476 = x7 & x3 & ~x5;
  assign n2477 = x7 & ~x2 & ~x5;
  assign n2478 = ~x3 & (n2480 | (~n605 & ~n2479));
  assign n2479 = (x0 | ~x1 | ~x4 | x6 | x7) & (~x0 | x1 | x4 | ~x6 | ~x7);
  assign n2480 = ~x2 & (x0 ? (n1445 & n978) : ~n2481);
  assign n2481 = (~x1 | ~x4 | ~x5 | x6 | ~x7) & (x1 | x4 | x5 | ~x6 | x7);
  assign n2482 = ~n2486 & (n2484 | n2485) & (n605 | n2483);
  assign n2483 = (x3 | x7 | ~x0 | x1) & (x0 | ~x1 | ~x7);
  assign n2484 = x3 & x7;
  assign n2485 = (x0 | ~x1 | ~x2 | x5) & (x2 | ~x5 | ~x0 | x1);
  assign n2486 = ~x7 & x5 & ~x2 & ~x0 & ~x1;
  assign n2487 = ~n2488 & ~n2491 & (~x5 | n697 | n2490);
  assign n2488 = ~n2489 & ~x5 & n927;
  assign n2489 = (~x0 | x2 | x4 | x6 | x7) & (x0 | ((~x2 | x4 | ~x6 | ~x7) & (x2 | ~x4 | x6 | x7)));
  assign n2490 = (~x0 | x1 | ~x3 | x4) & (x0 | (x1 ? (~x3 | ~x4) : (x3 | x4)));
  assign n2491 = ~x5 & ((n2492 & n1269) | (n743 & ~n2493));
  assign n2492 = x7 & x3 & x4;
  assign n2493 = (~x4 | ~x7 | ~x1 | x3) & (x4 | x7 | x1 | ~x3);
  assign z097 = n2495 | n2503 | ~n2506 | (~n1008 & ~n2498);
  assign n2495 = ~n765 & (x2 ? ~n2497 : ~n2496);
  assign n2496 = (x0 | ((~x3 | x6) & (x1 | ~x4 | (~x3 & x6)))) & (x1 | ~x3 | ~x4 | x6) & (~x0 | ~x1 | x3 | x4 | ~x6);
  assign n2497 = (x0 & (x1 | (~x3 & ~x4 & x6))) | (~x0 & ~x1 & (x3 | ~x6)) | (~x6 & (x3 | (x1 & x4)));
  assign n2498 = ~n2501 & ~n2502 & (x0 | (n2499 & n2500));
  assign n2499 = (x1 | ~x2 | ~x3 | x6) & (x3 | ~x6 | ~x1 | x2);
  assign n2500 = (~x1 | x6 | (x2 ? (~x3 | ~x4) : (x3 | x4))) & (x1 | x2 | x3 | x4 | ~x6);
  assign n2501 = x0 & ~x2 & ((~x3 & ~x6) | (~x1 & x3 & x6));
  assign n2502 = n560 & n2352;
  assign n2503 = ~n2504 & ~n2505;
  assign n2504 = x2 ? (x5 | x7) : (~x5 | ~x7);
  assign n2505 = (x0 | ~x1 | x3 | ~x4 | x6) & (x1 | x4 | (x0 ? (~x3 | x6) : (~x3 ^ ~x6)));
  assign n2506 = ~n2514 & ~n2512 & ~n2510 & ~n2507 & ~n2508;
  assign n2507 = n845 & n902 & n922;
  assign n2508 = ~x6 & ((n1268 & n733) | (n1365 & ~n2509));
  assign n2509 = x2 ? ~x5 : (x4 | x5);
  assign n2510 = ~n1164 & ((n1746 & n743) | (~x0 & ~n2511));
  assign n2511 = (~x2 | x3 | ~x5 | x6) & (x2 | ~x3 | x5 | ~x6);
  assign n2512 = ~n1820 & n2513;
  assign n2513 = ~x0 & ((x6 & x7 & ~x2 & ~x5) | (~x6 & ~x7 & x2 & x5));
  assign n2514 = x6 & n570 & (n2515 | (n681 & n622));
  assign n2515 = x5 & ~x0 & x3;
  assign z098 = n2517 | ~n2524 | ~n2532 | (~n643 & ~n2521);
  assign n2517 = ~x3 & (n2518 | (n560 & n662));
  assign n2518 = ~x5 & ((n742 & n2519) | (~x2 & ~n2520));
  assign n2519 = x6 & x7 & (x1 ^ ~x4);
  assign n2520 = (x0 | x1 | x4 | x6 | ~x7) & (~x0 | ~x4 | (x1 ? (x6 | x7) : (~x6 | ~x7)));
  assign n2521 = n2522 & ~n2523 & (x2 | n791 | n1820);
  assign n2522 = x0 ? (x3 | (x1 ? (x2 | ~x4) : x4)) : (~x3 | (x1 ? (x2 | ~x4) : (~x2 ^ ~x4)));
  assign n2523 = n570 & ((n2332 & n825) | (n1477 & n622));
  assign n2524 = n2526 & n2529 & (~x5 | ~n1188 | n2525);
  assign n2525 = (x0 | x2 | x4 | ~x6 | ~x7) & (~x0 | ~x2 | x6 | x7);
  assign n2526 = x2 ? (~n543 | n2527) : (n2341 | n2528);
  assign n2527 = x3 ? (~x4 | x6) : (x4 | ~x6);
  assign n2528 = x1 ? (x3 | x4) : (~x3 | ~x4);
  assign n2529 = (n647 | n2530) & (n856 | n2531);
  assign n2530 = (~x2 | ~x6 | ~x0 | x1) & (x0 | x6 | (x1 ^ ~x2));
  assign n2531 = (~x0 | x1 | ~x2 | ~x6 | ~x7) & (x0 | x6 | x7 | (x1 ^ ~x2));
  assign n2532 = ~n2536 & (x6 | n2533);
  assign n2533 = (~n1268 | ~n816) & (~n2332 | (~n2534 & ~n2535));
  assign n2534 = x3 & ~x2 & x0 & ~x1;
  assign n2535 = ~x0 & (x1 ? (x2 & x3) : (~x2 & ~x3));
  assign n2536 = ~n640 & ((n543 & n2537) | (~x1 & ~n2538));
  assign n2537 = x2 & (x3 ? (~x4 & ~x5) : (x4 & x5));
  assign n2538 = (x0 | ~x2 | x3 | x4 | ~x5) & (~x0 | ~x3 | x5 | (~x2 ^ ~x4));
  assign z099 = ~n2545 | (x1 ? ~n2540 : ~n2555);
  assign n2540 = ~n2544 & (x0 | (n2542 & (~n706 | n2541)));
  assign n2541 = (x2 | x3 | x4 | ~x7) & (~x2 | ~x3 | (~x4 ^ ~x7));
  assign n2542 = (~n1070 | ~n2385) & (n643 | n2543);
  assign n2543 = (~x2 | x3 | ~x4 | x5) & (x2 | ~x3 | x4 | ~x5);
  assign n2544 = n600 & n931;
  assign n2545 = ~n2546 & ~n2548 & ~n2550 & (x1 | n2552);
  assign n2546 = ~n1205 & ~n2547;
  assign n2547 = x1 ? ((x4 | x5 | ~x0 | x2) & (x0 | (x2 ? (x4 | x5) : (~x4 | ~x5)))) : ((~x2 | ~x4 | ~x5) & (x4 | x5 | x0 | x2));
  assign n2548 = ~n671 & ~n2549;
  assign n2549 = x1 ? ((x3 | ~x5 | ~x0 | x2) & (x0 | (x2 ? (x3 | ~x5) : x5))) : ((~x2 | ~x3 | x5) & (x3 | ~x5 | x0 | x2));
  assign n2550 = ~n714 & ((n841 & n2551) | (n742 & ~n2043));
  assign n2551 = x7 & ~x2 & x3;
  assign n2552 = n2554 & (~n2264 | ~n2553) & (~n547 | ~n635);
  assign n2553 = ~x4 & x0 & x3;
  assign n2554 = (x4 | x7 | ~x0 | x3) & (x0 | x2 | ~x3 | ~x4 | ~x7);
  assign n2555 = ~n2557 & (n1218 | n2558) & (~n1364 | n2556);
  assign n2556 = (x0 | ~x2 | ~x3 | x4 | x7) & (~x0 | ~x4 | (x2 ? (~x3 | ~x7) : (x3 | x7)));
  assign n2557 = ~n640 & ((n1181 & n639) | (x0 & n1268));
  assign n2558 = (x0 | ~x2 | x3 | x5 | ~x6) & (~x0 | x2 | ~x3 | ~x5 | x6);
  assign z100 = ~n2567 | n2574 | (x1 ? ~n2560 : ~n2564);
  assign n2560 = ~n2563 & (x0 | (~n2561 & (~n658 | ~n1780)));
  assign n2561 = ~x2 & (n2562 | (~x3 & ~n2055));
  assign n2562 = ~x7 & x6 & ~x5 & x3 & x4;
  assign n2563 = n600 & n1626;
  assign n2564 = (~x2 | ~x3 | n2566) & (x0 | x2 | x3 | ~n2565);
  assign n2565 = ~x4 & (x5 ? (x6 & ~x7) : (~x6 & x7));
  assign n2566 = (x0 | x4 | ~x5 | x6 | ~x7) & (~x4 | ((~x0 | (x5 ? (~x6 | ~x7) : (x6 | x7))) & (x0 | x5 | ~x6 | x7)));
  assign n2567 = ~n2568 & ~n2572 & ~n2573 & (x1 | n2571);
  assign n2568 = ~x3 & ((~n1198 & ~n2569) | (~n1957 & n2570));
  assign n2569 = x0 ? (~x4 | (x1 ^ ~x2)) : (x1 | x4);
  assign n2570 = x6 & x4 & ~x5;
  assign n2571 = (~x0 | x4 | ((x3 | x5) & (~x2 | ~x3 | ~x5))) & (x3 | ~x4 | ~x5 | (x0 & x2));
  assign n2572 = n1317 & ((n681 & n743) | (~x0 & ~n1134));
  assign n2573 = x3 & ~n2259 & (~x0 | n804);
  assign n2574 = ~n1353 & ((n746 & n2575) | (~x1 & ~n2576));
  assign n2575 = x7 & x3 & x5;
  assign n2576 = x0 ? (~x5 | (x2 ? (x3 | x7) : (~x3 | ~x7))) : (x5 | (x2 ? (x3 | ~x7) : (~x3 | x7)));
  assign z101 = n2588 | ~n2590 | (x1 ? ~n2578 : ~n2582);
  assign n2578 = ~n2581 & (x0 | (~n2580 & (x3 | n2579)));
  assign n2579 = x7 ? ((x2 | ~x4 | x5 | ~x6) & (x4 | ~x5 | x6)) : ((x5 | x6 | x2 | ~x4) & (~x2 | (x4 ? (~x5 | x6) : (x5 | ~x6))));
  assign n2580 = ~x6 & n1301 & ((x4 & ~x7) | (x2 & ~x4 & x7));
  assign n2581 = n588 & n594;
  assign n2582 = x2 ? (x6 | n2587) : n2583;
  assign n2583 = x3 ? (n2585 | (~n1395 & ~n2584)) : n2586;
  assign n2584 = x4 & (x6 ^ ~x7);
  assign n2585 = x0 ^ x5;
  assign n2586 = (x0 | ~x4 | x5 | x6 | x7) & (x4 | ((~x0 | ~x5 | ~x6 | x7) & (x0 | ~x7 | (~x5 ^ ~x6))));
  assign n2587 = (x0 | ~x3 | ~x4 | ~x5 | x7) & (~x7 | (x0 ? (x3 ? (~x4 | x5) : (x4 | ~x5)) : (x4 | (~x3 ^ ~x5))));
  assign n2588 = x0 & ((n592 & n576) | (x5 & ~n2589));
  assign n2589 = (~x1 | x2 | x3 | ~x4 | ~x6) & (x4 | ((x2 | x3 | x6) & (x1 | ~x3 | (x2 ^ ~x6))));
  assign n2590 = ~n2591 & ~n2597 & ~n2598 & (n1218 | n2594);
  assign n2591 = ~x0 & (x1 ? ~n2593 : ~n2592);
  assign n2592 = (x2 | ~x3 | ~x4 | ~x5 | x6) & (x4 | (x2 ? (x3 ? (x5 | x6) : (~x5 | ~x6)) : (x5 | ~x6)));
  assign n2593 = (x5 | ~x6 | ~x2 | ~x4) & (x2 | ~x5 | (x3 ? (x4 | ~x6) : (~x4 | x6)));
  assign n2594 = (x5 | n2595) & (~x2 | ~x5 | ~x6 | n2596);
  assign n2595 = (~x0 | ~x1 | x2 | x3 | x6) & (x0 | ~x6 | (x1 ? (x2 | ~x3) : ~x2));
  assign n2596 = x0 ? x1 : (~x1 | ~x3);
  assign n2597 = ~x4 & ((n904 & ~n823) | (n1380 & n1006));
  assign n2598 = n772 & ((n653 & n706) | (x0 & n1723));
  assign z102 = n2609 | ~n2613 | (x4 ? ~n2605 : ~n2600);
  assign n2600 = x0 ? (~n2602 & (x5 | n2601)) : n2603;
  assign n2601 = (~x1 | x2 | ~x3 | x6 | ~x7) & (x7 | ((x2 | (x6 ? x3 : x1)) & (x1 | (x3 & (~x2 | ~x6)))));
  assign n2602 = x7 & n551 & ((x2 & (~x3 | x6)) | (~x3 & x6) | (~x2 & x3 & ~x6));
  assign n2603 = x5 ? (~x7 | (n2604 & (~n885 | n1312))) : (x7 | n2604);
  assign n2604 = (~x1 | x6 | (~x2 & x3)) & (x1 | x2 | x3 | ~x6);
  assign n2605 = x0 ? (x1 | n2608) : (~n2606 & ~n2607);
  assign n2606 = ~x2 & ((n943 & n927) | (n689 & n942));
  assign n2607 = n2475 & ((x3 & ~x6) | (x1 & (x3 | ~x6)));
  assign n2608 = (x2 | ~x3 | (x5 ? ~x7 : (x6 | x7))) & (~x6 | ~x7 | ~x2 | ~x5) & (x5 | x7 | ((x3 | ~x6) & (~x2 | (x3 & ~x6))));
  assign n2609 = ~n1008 & (n2611 | ~n2612 | (x4 & ~n2610));
  assign n2610 = (~x0 | x1 | ~x2 | ~x3 | x6) & (x0 | x2 | (x1 ? x3 : (~x3 | ~x6)));
  assign n2611 = ~x2 & ((x0 & x1 & ~x3 & ~x6) | (~x0 & (x1 ? (x3 & x6) : ~x6)));
  assign n2612 = x0 | ~x2 | ((~x6 | ~n828) & (x1 | (~x6 & ~n828)));
  assign n2613 = ~n2615 & (n1548 | n2614);
  assign n2614 = (x0 | ~x1 | ~x2 | x5 | ~x6) & (x1 | ((~x0 | ~x2 | ~x5 | x6) & (x0 | (x2 ? (x5 | x6) : (~x5 | ~x6)))));
  assign n2615 = ~x2 & (n2616 | n2617 | (n704 & n699));
  assign n2616 = x0 & ~x1 & (x3 ? (~x5 & x6) : (x5 & ~x6));
  assign n2617 = x1 & ((x5 & x6 & x0 & ~x3) | (~x5 & ~x6 & ~x0 & x3));
  assign z103 = ~n2629 | n2626 | n2619 | n2624;
  assign n2619 = ~x2 & (~n2622 | (~x3 & ~n2620));
  assign n2620 = (~x5 | n2621) & (x5 | x6 | ~n1167 | n1543);
  assign n2621 = (x0 | ~x1 | ~x6 | ~x7) & (~x0 | x6 | x7 | (x1 ^ ~x4));
  assign n2622 = (~n866 | ~n2402) & (n640 | n2623);
  assign n2623 = (x0 | ~x1 | ~x3 | x4) & (~x0 | x1 | x3 | (~x4 ^ x5));
  assign n2624 = x1 & (x0 ? (n1044 & n696) : ~n2625);
  assign n2625 = x2 ? (x3 ? (~x4 | ~x6) : (x4 | x6)) : (~x4 | (x3 ? (~x5 | x6) : (x5 | ~x6)));
  assign n2626 = x2 & ((n601 & n866) | (~x1 & ~n2627));
  assign n2627 = (~n1070 | ~n2094) & (n640 | (n1433 & n2628));
  assign n2628 = (~x4 | ~x5 | ~x0 | x3) & (x4 | x5 | x0 | ~x3);
  assign n2629 = ~n2632 & (n643 | (n2631 & (x2 | n2630)));
  assign n2630 = (~x4 | ~x5 | x1 | x3) & (~x0 | ((x1 | ~x3 | ~x4 | x5) & (~x1 | x4 | (~x3 ^ x5))));
  assign n2631 = (x1 | x2 | ~x3 | x4) & (~x1 | ((x3 | ~x4 | ~x0 | x2) & (x0 | (x2 ? (~x3 ^ x4) : (x3 | x4)))));
  assign n2632 = ~x1 & (x6 ? ~n2633 : ~n2634);
  assign n2633 = (x2 | ~x3 | ~x4 | (x0 & ~x5)) & (x3 | x4 | (~x2 & (~x0 | x5)));
  assign n2634 = (x0 | x2 | x3 | (~x4 ^ x5)) & (~x2 | ~x3 | (~x4 & (x0 | ~x5)));
  assign z104 = n2641 | n2643 | ~n2645 | (~x3 & ~n2636);
  assign n2636 = ~n2637 & (~n560 | ~n1621) & (n643 | n2640);
  assign n2637 = ~x0 & ((n943 & n2638) | (~x2 & ~n2639));
  assign n2638 = ~x4 & ~x1 & x2;
  assign n2639 = (x1 | ~x4 | x5 | x6 | ~x7) & (~x1 | ~x5 | ~x6 | (x4 ^ ~x7));
  assign n2640 = (~x0 | ((x1 | ~x2 | ~x4 | x5) & (~x1 | x2 | x4 | ~x5))) & (x0 | ~x1 | x2 | x4 | x5);
  assign n2641 = x1 & ((n2435 & n2209) | (~x2 & ~n2642));
  assign n2642 = (x4 | ((~x0 | x5 | (x3 ^ ~x7)) & (x0 | x3 | ~x5 | x7))) & (x0 | ~x4 | ~x7 | (~x3 ^ ~x5));
  assign n2643 = ~x1 & (x3 ? (~n765 & ~n2185) : ~n2644);
  assign n2644 = x0 ? ((~x2 | ~x4 | ~x5 | x7) & (x2 | x4 | (~x5 ^ x7))) : ((x2 | ~x4 | ~x5 | x7) & (~x2 | x4 | x5 | ~x7));
  assign n2645 = n2646 & (~n825 | n2651) & (x1 | n2650);
  assign n2646 = ~n2649 & (~n746 | ~n2647) & (~n743 | ~n2648);
  assign n2647 = x7 & ~x3 & ~x4;
  assign n2648 = ~x7 & ~x3 & x4;
  assign n2649 = ~x0 & ((~x2 & x3 & ~x4 & ~x7) | (x2 & x4 & (x3 ^ ~x7)));
  assign n2650 = (x4 | x7 | ~x0 | ~x3) & (~x7 | (~x3 ^ ~x4) | (~x0 ^ ~x2));
  assign n2651 = x1 ? (n640 | n2652) : (~n1518 | ~n813);
  assign n2652 = x2 ? (x4 | ~x5) : (~x4 | x5);
  assign z105 = n2654 | n2656 | ~n2664 | (~x0 & ~n2659);
  assign n2654 = n898 & ((n576 & n1358) | (~x1 & ~n2655));
  assign n2655 = x2 ? ((x5 | ~x6 | x3 | x4) & (~x3 | (x4 ? (~x5 | ~x6) : (x5 | x6)))) : ((~x3 | x4 | ~x5 | x6) & (x3 | ~x4 | x5 | ~x6));
  assign n2656 = ~x1 & ((x5 & ~n2657) | (n2061 & ~n2658));
  assign n2657 = (x6 | (x0 ? (~x3 | ~x4) : (x2 ? (~x3 | x4) : (x3 | ~x4)))) & (~x0 | ~x4 | ~x6 | (x2 & x3));
  assign n2658 = (~x4 | ~x6 | ~x2 | x3) & (x6 | (x2 ? (~x3 ^ ~x4) : (~x3 | x4)));
  assign n2659 = ~n2663 & (~x4 | (n2661 & (~n570 | ~n2660)));
  assign n2660 = ~x7 & (x3 ? (~x5 & x6) : (x5 & ~x6));
  assign n2661 = (~n576 | ~n943) & (n627 | n2662);
  assign n2662 = (x1 | x2 | x5 | ~x7) & (~x1 | ~x2 | ~x5 | x7);
  assign n2663 = n828 & (x1 ? (~x7 & ~n538) : (x7 & ~n1447));
  assign n2664 = ~n2665 & n2667 & (n975 | n823 | n1685);
  assign n2665 = ~x0 & ~n2666;
  assign n2666 = (x5 | (x2 ? (x3 | ~x4) : (x4 | (x3 ^ ~x6)))) & (x2 | ~x4 | ((~x5 | ~x6) & (~x3 | (~x5 & ~x6))));
  assign n2667 = (n2259 | n2373) & (~n837 | ~n960);
  assign z106 = n2675 | ~n2677 | (~x0 & ~n2669);
  assign n2669 = x5 ? (~n2671 & (~x2 | n2670)) : n2672;
  assign n2670 = (~x1 | x3 | x4 | x6 | x7) & (~x4 | ((x1 | ~x3 | ~x6 | x7) & (~x7 | (x1 ? (~x3 ^ x6) : (x3 | x6)))));
  assign n2671 = n1084 & ((~x6 & ~x7 & ~x1 & x3) | (x6 & (x1 ? (x3 ^ x7) : (~x3 & ~x7))));
  assign n2672 = (~x2 | n2673) & (x1 | x2 | ~x4 | ~n2674);
  assign n2673 = (x1 | ~x3 | ~x4 | ~x6 | ~x7) & (x4 | ((x1 | ~x3 | x6 | x7) & (~x1 | (x3 ? (~x6 | x7) : (x6 | ~x7)))));
  assign n2674 = x7 & (x3 ^ x6);
  assign n2675 = x1 & (x0 ? (n1044 & n559) : ~n2676);
  assign n2676 = (x2 | ((~x5 | ((x4 | x6) & (x3 | ~x4 | ~x6))) & (~x3 | ((~x4 | x5 | ~x6) & (~x5 | x6))))) & (x3 | x5 | (x4 ? ~x2 : ~x6));
  assign n2677 = ~n2678 & ~n2681 & ~n2685 & (n1097 | n2684);
  assign n2678 = ~x1 & (x0 ? ~n2680 : ~n2679);
  assign n2679 = x2 ? ((x5 | x6 | x3 | x4) & (~x3 | ~x5 | (x4 & x6))) : (x3 ? (x5 | ~x6) : (~x5 | x6));
  assign n2680 = x4 ? (x2 ? (x5 | (x3 ^ ~x6)) : (~x5 | (~x3 & ~x6))) : ((x3 | ~x5 | x6) & (~x2 | ~x3 | x5 | ~x6));
  assign n2681 = n841 & (x2 ? ~n2683 : ~n2682);
  assign n2682 = (x3 | ~x6 | (x4 ? (x5 | ~x7) : (~x5 | x7))) & (x6 | ((x3 | ~x4 | ~x5 | x7) & (~x3 | (x4 ? (x5 | x7) : (~x5 | ~x7)))));
  assign n2683 = (~x3 | x4 | x5 | x6 | ~x7) & (x3 | ((x6 | x7 | ~x4 | ~x5) & (x4 | ~x6 | (~x5 ^ x7))));
  assign n2684 = x0 ? (x2 | x4 | (~x1 ^ x3)) : (~x2 | (x1 ? ~x3 : (x3 | ~x4)));
  assign n2685 = ~n765 & ((n744 & n1269) | (x4 & ~n2686));
  assign n2686 = (~x1 | x2 | x3 | x6) & (~x0 | x1 | ~x2 | ~x3 | ~x6);
  assign z107 = n2688 | ~n2691 | n2697 | (n1188 & ~n2700);
  assign n2688 = ~x0 & (n952 | (x1 & (n2689 | ~n2690)));
  assign n2689 = x2 & (n2562 | (~n643 & (n828 | n731)));
  assign n2690 = (~n1562 | ~n813) & (n640 | (~n545 & ~n2537));
  assign n2691 = ~n2694 & (x2 ? n2692 : (~n2695 & n2696));
  assign n2692 = (x1 | ~x3 | ~n728) & (x0 | ~x1 | n2693);
  assign n2693 = (~x5 | ~x6 | ~x3 | x4) & (x5 | x6 | x3 | ~x4);
  assign n2694 = ~n627 & ((~x4 & ~x5 & x1 & ~x2) | (~x1 & x4 & (x2 ^ x5)));
  assign n2695 = n1145 & ((n1723 & n536) | (~x0 & ~n975));
  assign n2696 = (~x0 | x1 | x3 | x4 | x6) & (x0 | ~x1 | ~x3 | ~x4 | ~x6);
  assign n2697 = ~x3 & ((~x2 & ~n2698) | (n570 & ~n2699));
  assign n2698 = (~x6 | (x4 ^ ~x5) | (~x1 ^ x7)) & (~x4 | x6 | (~x1 ^ ~x7));
  assign n2699 = x4 ? (~x5 | (~x6 ^ x7)) : (~x6 ^ ~x7);
  assign n2700 = x4 ? ((x6 | ~x7 | x2 | x5) & (~x2 | ((~x6 | ~x7) & (~x5 | x6 | x7)))) : ((~x6 ^ x7) | (x2 ^ ~x5));
  assign z108 = n2706 | ~n2710 | (~x2 & ~n2702);
  assign n2702 = ~n2704 & (x0 ? n2703 : (~n1317 | ~n2209));
  assign n2703 = (x5 | x7 | x3 | x4) & (~x1 | ((x4 | x5 | x7) & (x3 | (x4 ? (x5 | ~x7) : x7))));
  assign n2704 = ~n710 & (x3 ? (n674 | n2705) : ~n1337);
  assign n2705 = ~x4 & (x5 ^ ~x7);
  assign n2706 = ~x3 & (n2708 | (~n815 & ~n2707));
  assign n2707 = (x0 | x1 | x4 | x5 | x7) & (~x5 | (x0 & x1) | (~x4 ^ x7));
  assign n2708 = x1 & ((n813 & n2058) | (n743 & n2709));
  assign n2709 = x5 & x6 & (~x4 ^ ~x7);
  assign n2710 = ~n2711 & (n710 | n1190 | x5 | ~n1029);
  assign n2711 = n1890 & (n2712 | (~x7 & ~n856));
  assign n2712 = x7 & (x4 ^ ~x5);
  assign z109 = ~n2719 | n2714 | (~x6 & n681 & ~n2718);
  assign n2714 = ~x2 & (n2715 | (n588 & n712));
  assign n2715 = x1 & (x5 ? (n622 & ~n2717) : ~n2716);
  assign n2716 = (x6 | x7 | x0 | x4) & (~x0 | x3 | (x4 & x6));
  assign n2717 = (~x6 & ~x7) | (~x4 & (~x6 | ~x7));
  assign n2718 = x0 ? (x1 | x3) : ((x3 | ~x7) & (x1 | ~x3 | x7));
  assign n2719 = n710 | (n2721 & (n1205 | ~n2720));
  assign n2720 = x5 & (~x4 ^ ~x6);
  assign n2721 = x3 ? (x4 ? (x5 | ~x6) : (~x5 | x6)) : (x4 ? (~x5 ^ ~x6) : (x5 | ~x6));
  assign z110 = x5 ? (~n2732 & (n2723 | n2724)) : ~n2725;
  assign n2723 = ~x4 & (x6 ^ ~x7);
  assign n2724 = x4 & (~x6 ^ ~x7);
  assign n2725 = ~n2727 & (n2726 | n2730) & (~n596 | n2731);
  assign n2726 = x2 ^ x3;
  assign n2727 = ~x2 & (~n2729 | (x0 & ~n2728));
  assign n2728 = (~x4 | (x1 ? (x3 | ~x6) : (~x3 | (~x6 & x7)))) & (~x1 | x4 | x6 | (x3 & x7));
  assign n2729 = (~x3 | x4 | x6 | ~x7) & (x0 | ~x4 | (x6 ? ~x3 : x7));
  assign n2730 = (~x6 & (x4 | (~x0 & ~x1 & ~x7))) | (x0 & x1) | (~x4 & x6);
  assign n2731 = (x0 & (x1 | (x4 & ~x6))) | (x4 & ~x6 & x7) | (~x4 & (x6 | (~x0 & ~x7)));
  assign n2732 = x0 & x1 & (x2 | x3);
  assign z111 = n2734 | ~n2739 | (~x4 & ~n2736);
  assign n2734 = ~x7 & ((n746 & n960) | (~n1198 & ~n2735));
  assign n2735 = (x2 | ((x1 | ~x3) & (x0 | (~x3 & ~x4)))) & (x0 | ((~x2 | x3 | x4) & (x1 | (x3 & x4))));
  assign n2736 = (x5 | x7 | n2738) & (~x5 | ~x7 | ~n841 | n2737);
  assign n2737 = ~x2 & ~x3;
  assign n2738 = x0 ? (x1 ? (x2 | ~x3) : ~x2) : (~x1 | (~x2 ^ ~x3));
  assign n2739 = ~n2740 & ~n2741 & n2743 & (~n670 | ~n2435);
  assign n2740 = ~x2 & ((~x0 & x5 & x7) | (~x3 & ((x5 & x7) | (x0 & ~x5 & ~x7))));
  assign n2741 = n2742 & (n2475 | (n526 & n902));
  assign n2742 = x4 & x0 & ~x1;
  assign n2743 = (~n845 | ~n829) & (x0 | ~x2 | ~n526);
  assign z112 = ~n2746 | n2751 | n2754 | (~x6 & ~n2745);
  assign n2745 = x0 ? ((x1 | ~x2 | ~x3 | x7) & (~x1 | x2 | x3)) : (~x2 | (x1 ? (~x3 | x7) : (x3 | ~x7)));
  assign n2746 = ~n2747 & ~n2749 & ~n2750 & (~n626 | ~n1135);
  assign n2747 = ~n2748 & ~x7 & n742;
  assign n2748 = (x1 | ~x3 | x4 | x5 | ~x6) & (~x1 | x3 | ~x4 | (~x5 ^ x6));
  assign n2749 = ~x6 & ((~x0 & x1 & x7) | (~x1 & (x3 ? x7 : x0)));
  assign n2750 = ~n710 & n902 & x6 & ~x7;
  assign n2751 = ~x0 & (x4 ? ~n2752 : (n1317 & n2753));
  assign n2752 = (~x1 | x2 | x3 | ~x6 | x7) & (x1 | x6 | (x2 ? (~x3 | x7) : (x3 | ~x7)));
  assign n2753 = ~x7 & (x2 ^ ~x6);
  assign n2754 = ~x2 & ((n1244 & n1725) | (x0 & ~n2755));
  assign n2755 = (~x1 | ~x3 | x4 | ~n904) & (x1 | x3 | ~x4 | ~n978);
  assign z113 = ~n2762 | (~x0 & (~n2757 | ~n2761));
  assign n2757 = (~n2758 | ~n1439) & (~x7 | (~n2759 & (~n728 | ~n1439)));
  assign n2758 = ~x7 & x6 & ~x4 & x5;
  assign n2759 = ~x3 & ((n704 & n804) | (x1 & ~n2760));
  assign n2760 = (x2 | x4 | ~x5 | ~x6) & (x5 | x6 | ~x2 | ~x4);
  assign n2761 = (x1 | ~x2 | ~x3 | ~x4 | x7) & (x3 | ((x2 | ~x4 | ~x7) & (~x1 | x4 | (~x2 ^ ~x7))));
  assign n2762 = ~n2763 & n2764 & ~n2767 & (~n619 | n2768);
  assign n2763 = ~x3 & ((x0 & ~x7 & (~x1 ^ ~x2)) | (~x0 & ~x1 & x2 & x7));
  assign n2764 = ~n2766 & (~n560 | ~n2765) & (~n610 | ~n2144);
  assign n2765 = ~x7 & ~x3 & ~x4;
  assign n2766 = x3 & ((~x0 & ((~x2 & x7) | (x1 & x2 & ~x7))) | (~x1 & ((~x2 & x7) | (x0 & x2 & ~x7))));
  assign n2767 = ~x7 & ((n959 & n746) | (n1549 & ~n1820));
  assign n2768 = (~x0 | x2 | x3 | ~x4 | ~x5) & (x0 | x4 | (x2 ? (~x3 | x5) : (x3 | ~x5)));
  assign z114 = ~n2771 | n2774 | (~x1 & (~n2770 | ~n2776));
  assign n2770 = (x0 | x2 | x3 | ~x4) & (~x3 | (x0 ? (~x2 | x4) : (~x2 ^ ~x4)));
  assign n2771 = ~n2772 & n2773 & (x0 | ~x1 | n2726);
  assign n2772 = n1291 & ((n902 & n1786) | (n596 & n1668));
  assign n2773 = ~n1270 & (~n993 | ~n2144) & (~n1287 | ~n560);
  assign n2774 = ~x0 & ((n1133 & n959) | (~x1 & n2775));
  assign n2775 = ~x2 & (x3 ? (x4 & ~x5) : (~x4 & x5));
  assign n2776 = (~n549 | ~n926) & (~x6 | ~n1167 | n1515);
  assign z115 = n2778 | ~n2783 | (~x3 & ~n2782);
  assign n2778 = ~x2 & (n2779 | (n1241 & n1244));
  assign n2779 = ~x4 & ((n841 & ~n2780) | (x1 & ~n2781));
  assign n2780 = (~x3 | x5 | ~x6 | x7) & (x3 | ~x5 | x6 | ~x7);
  assign n2781 = (x0 | x5 | (x3 ? (x6 | ~x7) : (~x6 | x7))) & (~x0 | x3 | ~x5 | ~x6 | x7);
  assign n2782 = (x0 | ~x5 | (x1 ? (~x2 | ~x4) : x4)) & (x1 | ~x4 | ((x2 | x5) & (~x0 | (x2 & x5)))) & (x4 | ((x1 | ~x2) & (~x0 | ~x1 | x2 | x5)));
  assign n2783 = ~n2785 & n2788 & (~n632 | n2784);
  assign n2784 = (~x0 | x3 | x4 | ~x5 | x6) & (x0 | ((x5 | x6 | x3 | x4) & (~x3 | (x4 ? (~x5 | x6) : (x5 | ~x6)))));
  assign n2785 = ~x1 & ((n878 & ~n2786) | (x6 & ~n2787));
  assign n2786 = (x0 | x3 | ~x4 | ~x5) & (x4 | x5 | ~x0 | ~x3);
  assign n2787 = x0 ? ((~x2 | ~x3 | ~x4 | x5) & (x4 | ~x5 | x2 | x3)) : (x4 | (x2 ? (~x3 | ~x5) : (x3 | x5)));
  assign n2788 = (~x3 | n2789) & (~x2 | x3 | ~x4 | n2790);
  assign n2789 = (x1 | ~x2 | ~x4 | ~x5) & (x0 | ((~x1 | x2 | ~x4 | x5) & ((~x2 & ~x5) | (~x1 ^ x4))));
  assign n2790 = (~x5 | x6 | x7 | ~x0 | x1) & (x0 | x5 | (x1 ? (~x6 | ~x7) : (x6 | x7)));
  assign z116 = n2806 | (~x2 & (~n2792 | n2799 | ~n2802));
  assign n2792 = n2796 & ~n2793 & ~n2795;
  assign n2793 = ~x1 & ((n825 & n728) | (x0 & n2794));
  assign n2794 = ~x3 & (x4 ? (~x5 & ~x6) : (x5 & x6));
  assign n2795 = ~x0 & ((~x4 & x5 & (x1 | ~x3)) | (~x1 & x3 & (x4 ^ ~x5)));
  assign n2796 = (~x6 | n1134 | ~n2797) & (~x0 | n2798);
  assign n2797 = x3 & ~x0 & x1;
  assign n2798 = (~x1 | x3 | ~x4 | x5) & (x1 | ~x3 | x4 | ~x5);
  assign n2799 = ~x5 & ((x4 & ~n2800) | (n1167 & ~n2801));
  assign n2800 = x0 ? (x1 | (x3 ? (x6 | ~x7) : (~x6 | x7))) : (~x1 | x3 | (~x6 ^ x7));
  assign n2801 = (x1 | x3 | ~x6 | x7) & (~x1 | ~x3 | x6 | ~x7);
  assign n2802 = (n2803 | n2804) & (~n526 | ~n689 | n2805);
  assign n2803 = x4 ? (x6 | x7) : (~x6 | ~x7);
  assign n2804 = x0 ? (x1 ? (x3 | ~x5) : (~x3 | x5)) : (x3 | x5);
  assign n2805 = x0 ? (x4 | x6) : (~x4 | ~x6);
  assign n2806 = x2 & (n2810 | ~n2812 | n2807 | n2809);
  assign n2807 = ~x7 & ((n559 & n1244) | (~x4 & ~n2808));
  assign n2808 = (x0 | x1 | x3 | x5 | ~x6) & ((~x3 ^ x5) | (x0 ? (x1 | ~x6) : (~x1 | x6)));
  assign n2809 = ~x1 & ((~n615 & n1380) | (~n1353 & ~n2176));
  assign n2810 = ~n2811 & x7 & n1392;
  assign n2811 = (~x0 | x1 | ~x5 | x6) & (x0 | x5 | (~x1 ^ ~x6));
  assign n2812 = ~n2813 & ~n2814 & (~n1358 | ~n866);
  assign n2813 = ~x1 & ((x4 & ~x5 & ~x0 & x3) | (x0 & (x3 ? (x4 & x5) : (~x4 & ~x5))));
  assign n2814 = ~x0 & x1 & (x3 ? (x4 & ~x5) : (x4 ^ ~x5));
  assign z117 = ~n2821 | ~n2828 | (~x3 & ~n2816);
  assign n2816 = ~n2818 & (~n704 | ~n816) & (~x5 | n2817);
  assign n2817 = (x1 | x2 | (x0 ^ (x4 | x6))) & (x0 | ~x1 | ((~x2 | x4 | ~x6) & (~x4 | x6)));
  assign n2818 = ~n1954 & (n2820 | (x0 & ~n2819));
  assign n2819 = x4 ? (~x5 | ~x6) : (x5 | x6);
  assign n2820 = ~x6 & x5 & ~x0 & ~x4;
  assign n2821 = (~x3 | n2825) & (n765 | (n2823 & (x3 | n2822)));
  assign n2822 = (~x0 | x1 | x2 | x4 | x6) & (x0 | ((x1 | ~x4 | ~x6) & (x4 | x6 | ~x1 | ~x2)));
  assign n2823 = (~n2446 | n2824) & (n1408 | (~n587 & ~n1101));
  assign n2824 = x1 ? ~x6 : (x2 | x6);
  assign n2825 = ~n2827 & (~n577 | ~n816) & (~n543 | ~n2826);
  assign n2826 = ~x5 & (~x4 ^ ~x6);
  assign n2827 = ~x1 & ((~x5 & ~x6 & ~x0 & ~x4) | (x0 & (x4 ? (~x5 & x6) : (x5 & ~x6))));
  assign n2828 = x1 ? (~n2563 & ~n2833) : (~n2829 & ~n2831);
  assign n2829 = ~n2830 & ((x2 & x4 & ~x6) | (~x0 & (x4 | (x2 & x6))));
  assign n2830 = x3 ? (~x5 | x7) : (x5 | ~x7);
  assign n2831 = x0 & ((n1070 & n2385) | (x3 & ~n2832));
  assign n2832 = (x2 | ~x4 | ~x5 | x6 | x7) & (x4 | ~x6 | (~x5 ^ x7));
  assign n2833 = ~x0 & (n2835 | n2836 | (n1044 & n2834));
  assign n2834 = x7 & ~x4 & x6;
  assign n2835 = x3 & ~x4 & ~x6 & (x5 ^ x7);
  assign n2836 = x4 & x6 & (x3 ? (x5 & ~x7) : (~x5 & x7));
  assign z118 = ~n2850 | n2848 | n2845 | n2838 | n2842;
  assign n2838 = ~x2 & (n2839 | (n727 & n931));
  assign n2839 = ~x3 & ((x5 & ~n2840) | (n1310 & ~n2841));
  assign n2840 = x0 ? (x1 | (x4 ? (~x6 | x7) : (x6 | ~x7))) : (~x1 | x7 | (~x4 ^ x6));
  assign n2841 = (x1 | ~x4 | x6 | ~x7) & (~x1 | (~x6 ^ ~x7));
  assign n2842 = ~n1218 & (~n2844 | (~x2 & ~n2843));
  assign n2843 = (~x3 | ((x0 | x5 | (~x1 ^ ~x6)) & (~x0 | x1 | ~x5 | x6))) & (~x0 | x3 | (x1 ? (~x5 | x6) : (x5 | ~x6)));
  assign n2844 = (x0 | ~x1 | ~x2 | x5 | ~x6) & (x1 | ((~x0 | ~x2 | ~x5 | x6) & (x0 | ((~x5 | ~x6) & (~x2 | x5 | x6)))));
  assign n2845 = ~n671 & (~n2847 | (n1467 & ~n2846));
  assign n2846 = (x3 | x6 | ~x0 | x2) & (x0 | ~x2 | ~x6);
  assign n2847 = (~x0 | ~x1 | x2 | x3 | ~x6) & ((~x2 & ~x3) | (x0 ? (x1 | ~x6) : (~x1 | x6)));
  assign n2848 = ~x6 & (n1510 | (x0 & ~x4 & n2849));
  assign n2849 = ~x5 & (x1 ^ x2);
  assign n2850 = (~n2851 | ~n895) & (~n1686 | n2852);
  assign n2851 = ~x6 & (x3 ? (~x4 & ~x5) : (x4 & x5));
  assign n2852 = (~x1 | ~x4 | ~x5) & (x4 | x5 | x1 | x2);
  assign z119 = ~n2859 | n2865 | n2866 | (~x1 & ~n2854);
  assign n2854 = x2 ? (x0 | ~n992) : (~n2855 & n2856);
  assign n2855 = ~n1097 & ((~x4 & ~x7 & x0 & ~x3) | (~x0 & x7 & (~x3 | x4)));
  assign n2856 = (~n2857 | ~n951) & (n765 | n2858);
  assign n2857 = ~x4 & ~x0 & x3;
  assign n2858 = (~x0 | x3 | ~x4 | x6) & (x0 | ~x3 | x4 | ~x6);
  assign n2859 = ~n2860 & ~n2863 & (x5 | ~n793 | n1543);
  assign n2860 = n543 & ((~n2861 & n2862) | (n1556 & n951));
  assign n2861 = ~x4 & ~x2 & ~x3;
  assign n2862 = ~x7 & (x5 ^ ~x6);
  assign n2863 = ~n2737 & ((n841 & n1429) | (~x0 & ~n2864));
  assign n2864 = x1 ? (x5 | ~x7) : (~x5 | x7);
  assign n2865 = n632 & (x0 ? (x3 & n2209) : (~x3 & ~n1337));
  assign n2866 = ~n1198 & ~n2867;
  assign n2867 = (x2 | x3 | (x0 ? (~x1 | ~x7) : (x1 | x7))) & (~x0 | x1 | ~x7 | (~x2 & ~x3));
  assign z120 = n2873 | n2876 | (~x2 & (n2869 | n2870));
  assign n2869 = x0 & ((n813 & n945) | (n530 & n944));
  assign n2870 = ~x0 & ((n658 & n2871) | (n2315 & ~n2872));
  assign n2871 = ~x4 & x1 & ~x3;
  assign n2872 = x3 & (x4 | (x5 & ~x7));
  assign n2873 = ~n640 & (n2874 | n2875 | n880 | n2330);
  assign n2874 = ~x1 & (x2 | (x0 & x3));
  assign n2875 = n1287 & n733;
  assign n2876 = ~n643 & (~n2877 | (n560 & n1268));
  assign n2877 = (~x0 | x1 | x2 | x3 | x4) & (x0 | ~x1 | (~x2 & ~x3 & ~x4));
  assign z121 = n2879 | ~n2882 | (x7 & (n2330 | ~n2881));
  assign n2879 = n1084 & (n2880 | (n951 & n1234));
  assign n2880 = n626 & (n1500 | (x3 & n1383));
  assign n2881 = x0 ? (x1 & (x2 | x3)) : (~x1 & ~x2);
  assign n2882 = ~n2883 & (~n816 | ~n2648);
  assign n2883 = n1084 & ~n1566 & ~x7 & n626;
  assign z122 = ~n2891 | n2890 | n2885 | n2887;
  assign n2885 = ~x4 & (x3 ? ~n2886 : (n1723 & n816));
  assign n2886 = (~x0 | ~x1 | x2 | x5 | x6) & (x0 | ~x5 | (x1 ? (~x2 | ~x6) : (x2 | x6)));
  assign n2887 = ~x4 & ((n837 & n2888) | (n1910 & ~n2889));
  assign n2888 = ~x7 & x6 & x3 & ~x5;
  assign n2889 = (x3 | x5 | x1 | x2) & (~x3 | ~x5 | ~x1 | ~x2);
  assign n2890 = x4 & ((x0 & (~x1 | (~x2 & ~x3))) | (~x1 & ~x2 & ~x3) | (x2 & x3 & ~x0 & x1));
  assign n2891 = x0 ? (x4 | (x1 & ~n576)) : (x1 | ~n2892);
  assign n2892 = ~x2 & ~x4 & (x3 ^ x5);
  assign z123 = ~n2896 | (~x0 & ~n2894) | (n1084 & ~n2895);
  assign n2894 = (x2 | x3 | x4 | (~x1 ^ x5)) & (~x3 | ((x1 | ~x2 | ~x4 | ~x5) & (x4 | (x1 ? (x2 ^ ~x5) : (x2 | x5)))));
  assign n2895 = (~x0 | ~x1 | ~x3 | x5 | x6) & (x0 | (x1 ? (x3 ? (x5 | ~x6) : (~x5 | x6)) : (x3 ? (~x5 | x6) : (x5 | ~x6))));
  assign n2896 = ~n2897 & n2901 & (~x6 | (~n2899 & ~n2900));
  assign n2897 = ~n2898 & ~x6 & n1167;
  assign n2898 = (x1 | x2 | x3 | x5 | ~x7) & (~x1 | ~x3 | (x2 ? (~x5 | x7) : (x5 | ~x7)));
  assign n2899 = x0 & ((n979 & n2209) | (n717 & n676));
  assign n2900 = ~x0 & ((n635 & n1439) | (n576 & n809));
  assign n2901 = x0 ? (x1 ? (x2 | x3) : (~x2 | ~x3)) : ((x3 | ~x4 | x1 | x2) & (~x1 | (x2 ? x3 : (~x3 | ~x4))));
  assign z124 = n2903 | ~n2911 | (n772 & ~n2908);
  assign n2903 = ~x4 & (n2905 | (n560 & n2904));
  assign n2904 = x7 & x6 & ~x3 & x5;
  assign n2905 = x1 & ((~x2 & ~n2906) | (~x0 & n2907));
  assign n2906 = (x0 | x3 | ~x5 | ~x6 | ~x7) & (x5 | ((x0 | ~x3 | x6 | x7) & (~x0 | (x3 ? (~x6 | x7) : (x6 | ~x7)))));
  assign n2907 = x2 & ((x6 & x7 & ~x3 & ~x5) | (~x6 & ~x7 & x3 & x5));
  assign n2908 = (~x2 | n2910) & (~x5 | ~n2909 | ~x0 | x2);
  assign n2909 = ~x6 & (~x3 ^ x7);
  assign n2910 = (~x0 | x3 | ~x5 | ~x6 | x7) & (x0 | x5 | (x3 ? (~x6 | x7) : (x6 | ~x7)));
  assign n2911 = x2 ? n2914 : (x0 ? n2912 : n2913);
  assign n2912 = x3 ? ((x5 | x6 | ~x1 | x4) & (~x5 | ~x6 | x1 | ~x4)) : ((~x4 | x5) & (~x1 | (~x5 & ~x6)));
  assign n2913 = (x3 & (x4 | (x5 & x6))) | (~x4 & (x1 | (~x3 & ~x5)));
  assign n2914 = n2916 & (~n772 | n2915);
  assign n2915 = (~x0 | x3 | ~x5 | x6) & (x0 | x5 | (~x3 ^ x6));
  assign n2916 = (x3 | (x0 ? (x1 | (x4 & x5)) : ((~x4 | ~x5) & (~x1 | (~x4 & ~x5))))) & (x0 | ~x3 | x4 | (x1 & x5));
  assign z125 = n2918 | ~n2920 | n2926 | (~x0 & ~n2930);
  assign n2918 = n898 & ((n559 & n676) | (~x2 & ~n2919));
  assign n2919 = (x1 | ~x3 | ~x4 | ~x5 | x6) & (x4 | ((x1 | x3 | ~x5 | ~x6) & (~x1 | x5 | (~x3 ^ ~x6))));
  assign n2920 = ~n2923 & (x0 ? n2921 : n2922);
  assign n2921 = (~x1 | x2 | x3 | ~x4 | ~x5) & (x1 | ((x2 | x4 | (~x3 ^ ~x5)) & (~x4 | ((~x3 | x5) & (~x2 | (~x3 & x5))))));
  assign n2922 = (x4 | ((~x3 | x5 | (~x1 ^ ~x2)) & (x1 | ~x2 | (x3 & ~x5)))) & (~x1 | ~x4 | ((x3 | ~x5) & (x2 | (x3 & ~x5))));
  assign n2923 = x2 & ((n543 & ~n928) | (~n2924 & n2925));
  assign n2924 = x0 ? (x3 | ~x5) : (~x3 | x5);
  assign n2925 = ~x1 & (~x4 ^ ~x6);
  assign n2926 = ~x2 & (~n2928 | (~x0 & ~n2927));
  assign n2927 = (x1 | x3 | x4 | x5 | ~x6) & (~x1 | ((x3 | x4 | ~x5 | x6) & (x5 | ~x6 | ~x3 | ~x4)));
  assign n2928 = (n752 | n2929) & (~n661 | ~n728);
  assign n2929 = x0 ? (~x1 | x5) : (x1 | ~x5);
  assign n2930 = ~n2931 & ((~x2 & n981) | ~n2933 | (x2 & n1932));
  assign n2931 = ~x1 & ((n1556 & n951) | (n2932 & ~n2504));
  assign n2932 = x4 & (~x3 ^ x6);
  assign n2933 = ~x7 & x1 & ~x4;
  assign z126 = n2945 | ~n2948 | (x4 ? ~n2941 : ~n2935);
  assign n2935 = ~n2938 & (x2 | (~n2937 & (x3 | n2936)));
  assign n2936 = (~x0 | x7 | (x1 ? (x5 | x6) : (~x5 | ~x6))) & (~x7 | ((x5 | ~x6 | ~x0 | x1) & (x0 | (x1 ? (~x5 | ~x6) : (x5 | x6)))));
  assign n2937 = n927 & ((x0 & ~x5 & x6 & ~x7) | (~x0 & ~x6 & (x5 ^ ~x7)));
  assign n2938 = n2940 & (n2388 | n2939);
  assign n2939 = ~x7 & ~x6 & x3 & x5;
  assign n2940 = x2 & ~x0 & x1;
  assign n2941 = x1 ? (~x7 | n2942) : (x7 ? n2943 : n2944);
  assign n2942 = (x0 | ~x2 | ~x3 | x5 | x6) & (~x0 | x2 | x3 | ~x5 | ~x6);
  assign n2943 = x2 ? (x0 ? (x3 ? (~x5 | x6) : (x5 | ~x6)) : (~x5 | (~x3 ^ ~x6))) : ((~x5 | ~x6 | ~x0 | x3) & (x0 | x5 | (~x3 ^ ~x6)));
  assign n2944 = (~x5 | ((~x0 | (x2 ? (x3 | ~x6) : x6)) & (x2 | ((x3 | x6) & (x0 | ~x3 | ~x6))))) & (x0 | ~x2 | x5 | (~x3 ^ ~x6));
  assign n2945 = ~x2 & ((x3 & ~n2946) | (n653 & ~n2947));
  assign n2946 = x0 ? (x5 | (x1 & (x4 | x6))) : (~x4 | ~x5 | (~x1 ^ ~x6));
  assign n2947 = x1 ? (~x4 | ~x5) : (x5 | ~x6);
  assign n2948 = ~n2949 & ~n2952 & ~n2954 & (n1198 | n2951);
  assign n2949 = x2 & ((n696 & n699) | (~x1 & ~n2950));
  assign n2950 = (~x3 | ((~x0 | ~x5 | ~x6) & (x5 | x6 | x0 | x4))) & (x0 | x3 | ~x5 | (x4 & ~x6));
  assign n2951 = (~x2 | x3 | x4 | ~x0 | x1) & (x0 | ~x3 | (x1 ? (~x2 | ~x4) : (x2 | x4)));
  assign n2952 = ~n2259 & ~n2953;
  assign n2953 = (x2 | x3 | ~x0 | ~x1) & (x0 | ~x3 | (x1 ^ ~x2));
  assign n2954 = ~n1564 & (n2955 | (~x0 & n1093));
  assign n2955 = ~x6 & x5 & x0 & ~x1;
  assign z127 = ~n2963 | n2969 | (x5 ? ~n2972 : ~n2957);
  assign n2957 = x3 ? n2960 : (~n2958 & (x1 | n2959));
  assign n2958 = ~n1998 & ((n1445 & n1857) | (n1300 & n772));
  assign n2959 = (~x0 | x2 | x4 | x6 | x7) & (~x4 | ((~x2 | x6 | x7) & (x0 | ((x6 | x7) & (x2 | ~x6 | ~x7)))));
  assign n2960 = x2 ? n2961 : n2962;
  assign n2961 = (~x6 | ~x7 | ~x0 | x1) & (x0 | ((~x4 | x6 | x7) & (~x1 | x4 | ~x6 | ~x7)));
  assign n2962 = (~x0 | x1 | ~x4 | ~x6 | ~x7) & (x0 | ~x1 | x4 | (~x6 ^ ~x7));
  assign n2963 = ~n2966 & (n643 | (x0 & n2964) | (~x0 & n2965));
  assign n2964 = x3 ? (x4 | x5 | (~x1 ^ x2)) : ((x2 | ~x4 | ~x5) & (x1 | (x2 & ~x4)));
  assign n2965 = (x1 | ~x3 | ~x4) & (x3 | x4 | ~x1 | ~x2);
  assign n2966 = x3 & (~n2968 | (n1966 & ~n2967));
  assign n2967 = (x0 | ~x1 | ~x4 | x6) & (x4 | ~x6 | ~x0 | x1);
  assign n2968 = (~x0 | x1 | x2 | x4 | ~x6) & (x0 | x6 | (x1 ? (x2 | ~x4) : x4));
  assign n2969 = ~x3 & ((~n2341 & ~n2970) | (n1686 & ~n2971));
  assign n2970 = x1 ? (x2 | (~x4 ^ x5)) : (~x2 | x4);
  assign n2971 = x4 ? (~x1 | (~x2 & ~x5)) : (x2 | (x1 & x5));
  assign n2972 = (~n816 | ~n1525) & (n640 | n2973);
  assign n2973 = (~x3 | ~x4 | ~x0 | x1) & (x0 | ((~x1 | ~x3 | x4) & (x1 | ~x2 | x3 | ~x4)));
  assign z128 = n2975 | n2978 | ~n2986 | (~x0 & ~n2985);
  assign n2975 = ~x4 & ((~x5 & ~n2976) | (n691 & ~n2977));
  assign n2976 = (x0 | ~x1 | x2 | ~x3 | x7) & (~x7 | ((x2 | x3 | x0 | ~x1) & (x1 | (x0 ? (~x2 ^ x3) : (~x2 | ~x3)))));
  assign n2977 = (x3 | x7 | ~x0 | x1) & (x0 | ~x1 | (~x3 ^ x7));
  assign n2978 = ~x1 & (n2983 | (~x2 & (n2979 | ~n2981)));
  assign n2979 = ~n1353 & ((n526 & n653) | (x0 & n2980));
  assign n2980 = ~x5 & (~x3 ^ ~x7);
  assign n2981 = (~n2857 | ~n943) & (x7 | ~n622 | n2982);
  assign n2982 = x4 ? (~x5 ^ ~x6) : (x5 | ~x6);
  assign n2983 = n2371 & ~n2984;
  assign n2984 = (~x3 | x7 | (~x4 ^ ~x6)) & (~x0 | (x4 ? (~x6 ^ x7) : ((x6 | x7) & (~x3 | ~x6 | ~x7))));
  assign n2985 = (~x1 | ~x2 | x4 | ~x5 | x7) & (~x4 | ((x1 | x2 | ~x5 | x7) & (~x1 | ~x7 | (x2 & ~x5))));
  assign n2986 = ~n2988 & n2991 & (n671 | n2987);
  assign n2987 = (~x5 | ((x1 | ~x2) & (~x0 | (x1 ? (x2 | x3) : ~x3)))) & (x0 | x1 | x5 | (x2 & x3));
  assign n2988 = n1093 & ((~n1408 & ~n2989) | (~x0 & ~n2990));
  assign n2989 = (x0 | ~x2 | x7) & (x3 | ~x7 | ~x0 | x2);
  assign n2990 = (x2 | x3 | x4 | x6 | x7) & (~x2 | ~x3 | ~x4 | ~x6 | ~x7);
  assign n2991 = (~n837 | ~n2209) & (~n746 | ~n2992);
  assign n2992 = x7 & ~x5 & ~x3 & x4;
  assign z129 = x1 ? ~n3002 : (x3 ? ~n2994 : ~n2997);
  assign n2994 = x6 ? n2995 : (n2996 & (n1008 | n1998));
  assign n2995 = (~x0 | (x5 & (~x2 | ~x4 | x7))) & (x0 | x2 | x4 | ~x5 | ~x7) & (x5 | (~x2 & ~x4 & x7));
  assign n2996 = x0 ? (~x2 | ~x5) : (x2 | x5);
  assign n2997 = ~n2998 & ~n3000 & n3001 & (~n995 | ~n2999);
  assign n2998 = ~x0 & ((~x2 & x5 & x6 & x7) | (x2 & ~x5 & (x6 | ~x7)));
  assign n2999 = ~x6 & x7 & (x4 ^ ~x5);
  assign n3000 = ~x2 & ((n564 & n943) | (~x0 & n670));
  assign n3001 = (x0 | x5 | x6 | ~x7) & (~x0 | (x5 ? (x6 | x7) : ~x6));
  assign n3002 = ~n3003 & (~n825 | n3006) & (x3 | n3005);
  assign n3003 = ~x0 & ((n530 & n1556) | (~x6 & ~n3004));
  assign n3004 = x2 ? (~x3 | ~x7 | (~x4 ^ ~x5)) : (x3 | x7 | (~x4 ^ x5));
  assign n3005 = (x2 | ((x5 | ~x6 | ~x7) & (~x0 | ~x5 | (x6 & x7)))) & (x0 | ((~x6 & ~x7) ? (~x2 | ~x5) : x5));
  assign n3006 = (x5 | (x2 & ~x6)) & (x6 | x7 | ~x2 | ~x5);
  assign z130 = x2 ? ~n3019 : (n3008 | ~n3011);
  assign n3008 = ~x6 & ((~x5 & ~n3009) | (n526 & ~n3010));
  assign n3009 = (x0 | ~x1 | x3 | (~x4 ^ x7)) & (~x3 | ((x0 | x1 | ~x4 | x7) & (~x0 | (x1 ? (x4 | x7) : ~x7))));
  assign n3010 = (x3 | x4 | x0 | ~x1) & (~x0 | x1 | (~x3 & ~x4));
  assign n3011 = ~n3012 & ~n3015 & n3017 & (n640 | n3014);
  assign n3012 = ~x0 & ~n3013;
  assign n3013 = (x1 | ~x3 | ~x4 | ~x5 | x6) & (x3 | ((x5 | ~x6 | x1 | x4) & (~x1 | ~x5 | (~x4 ^ x6))));
  assign n3014 = (x3 | (x0 ? ~x1 : (x1 | ~x4))) & (x0 | x1 | x4 | (~x3 & ~x5));
  assign n3015 = n569 & (n712 | n3016);
  assign n3016 = ~x5 & ~x4 & ~x3 & ~x0 & x1;
  assign n3017 = ~n3018 & (~n841 | ~n744) & (~n592 | ~n661);
  assign n3018 = ~x6 & x3 & ~x0 & x1;
  assign n3019 = ~n3024 & n3020 & ~n3023;
  assign n3020 = ~n3022 & (~n712 | ~n1668) & (~n543 | ~n3021);
  assign n3021 = x6 & x3 & x4;
  assign n3022 = ~x1 & (x0 ? (x6 & (x3 ^ x4)) : (~x3 & ~x6));
  assign n3023 = ~n643 & ((~x0 & (x3 ? ~x4 : x1)) | (~x1 & (x0 ? (~x3 & ~x4) : x3)));
  assign n3024 = x6 & ((n866 & n867) | (n841 & ~n3025));
  assign n3025 = (x3 | x4 | ~x5 | ~x7) & (x5 | x7 | ~x3 | ~x4);
  assign z131 = ~n3035 | n3033 | n3027 | n3030;
  assign n3027 = ~x6 & (n3028 | (n1209 & n923));
  assign n3028 = x7 & (x4 ? (n1181 & n2112) : ~n3029);
  assign n3029 = (x0 | ~x1 | ~x2 | ~x3 | ~x5) & (~x0 | ((~x1 | x2 | ~x3 | x5) & (x1 | ~x2 | x3 | ~x5)));
  assign n3030 = ~x0 & (n3031 | (x5 & n804 & ~n2017));
  assign n3031 = x1 & (n3032 | (n674 & n1044));
  assign n3032 = x7 & ~x5 & ~x4 & x2 & x3;
  assign n3033 = n3034 & (n1598 | (x3 & n2316));
  assign n3034 = x2 & x0 & ~x1;
  assign n3035 = n3037 & ~n3041 & (x0 | ~x1 | n3036);
  assign n3036 = (x2 | x3 | x4 | ~x7) & (~x2 | ~x3 | ~x4 | x7);
  assign n3037 = ~n3039 & ~n3040 & (x1 | n1548 | n3038);
  assign n3038 = x0 ? (~x2 | x7) : (x2 | ~x7);
  assign n3039 = ~x7 & x3 & ~x2 & ~x0 & x1;
  assign n3040 = (~x0 ^ ~x2) & (x1 ? (~x3 & x7) : (x3 ^ ~x7));
  assign n3041 = ~n3042 & n1181 & ~x7 & n1723;
  assign n3042 = x1 ? (x3 | ~x4) : (~x3 ^ ~x4);
  assign z132 = n3044 | n3048 | ~n3053 | (n564 & ~n3052);
  assign n3044 = x5 & (n3045 | (~n790 & n3047));
  assign n3045 = ~x1 & ((n547 & n1668) | (x2 & ~n3046));
  assign n3046 = (x0 | x3 | x4 | x6 | ~x7) & (~x0 | x7 | (x3 ? (~x4 | x6) : (x4 | ~x6)));
  assign n3047 = ~x4 & x3 & ~x0 & x1;
  assign n3048 = ~x0 & ((n3050 & n3051) | (~x4 & ~n3049));
  assign n3049 = (x1 | x2 | x3 | x5 | ~x6) & (~x5 | ((x1 | ~x2 | x3 | ~x6) & (~x1 | ~x3 | (x2 ^ ~x6))));
  assign n3050 = ~x6 & (x1 ^ x3);
  assign n3051 = ~x5 & ~x2 & x4;
  assign n3052 = (~x3 | x5 | x6 | ~x1 | x2) & (x1 | ((~x2 | (x3 ? (x5 | ~x6) : (~x5 | x6))) & (x5 | ~x6 | x2 | x3)));
  assign n3053 = ~n3056 & n3058 & (x2 ? n3054 : n3055);
  assign n3054 = x0 ? (x1 | (x3 ? (~x4 ^ x5) : (x4 | x5))) : ((x1 | ~x3 | ~x4 | ~x5) & (~x1 | (x3 ? (x4 | x5) : (~x4 | ~x5))));
  assign n3055 = x0 ? (x3 | ~x4) : (x1 ? (~x3 ^ ~x4) : (~x3 | x4));
  assign n3056 = n1632 & ((n2155 & n626) | (n3057 & n922));
  assign n3057 = ~x7 & x3 & x6;
  assign n3058 = (~n626 | ~n1489) & (~x5 | n1744 | ~n895);
  assign z133 = ~n3071 | n3068 | n3060 | n3065;
  assign n3060 = ~x4 & (x1 ? ~n3061 : ~n3063);
  assign n3061 = (x2 | n3062) & (x0 | ~x2 | ~x3 | n1647);
  assign n3062 = (x0 | ~x3 | ~x5 | x6 | x7) & (x5 | ((x0 | x3 | x6 | ~x7) & (~x0 | ~x6 | (x3 ^ ~x7))));
  assign n3063 = (~n1693 | ~n943) & (x3 | n3064);
  assign n3064 = (x0 | x2 | x5 | x6 | ~x7) & (~x2 | ((~x0 | (x5 ? (~x6 | x7) : (x6 | ~x7))) & (x6 | x7 | x0 | ~x5)));
  assign n3065 = x6 & ((~x1 & ~n3066) | (n543 & ~n3067));
  assign n3066 = (x2 | ((~x3 | x4 | ~x5) & (~x0 | x3 | ~x4 | x5))) & (x4 | ((x0 | ~x3 | ~x5) & (~x2 | x3 | x5)));
  assign n3067 = x3 ? (~x4 | ~x5) : (x5 | (x2 ^ x4));
  assign n3068 = x4 & ((n733 & n1925) | (~x1 & ~n3069));
  assign n3069 = (~x2 | n3070) & (x3 | n1647 | x0 | x2);
  assign n3070 = (~x0 | ~x3 | ~x5 | x6 | x7) & (x0 | x3 | x5 | ~x6 | ~x7);
  assign n3071 = n3073 & (n1566 | n3072);
  assign n3072 = (x0 & (x6 ? ~x4 : x2)) | (x4 & (x1 | (~x0 & ~x2 & x6))) | (~x4 & (~x1 | (x2 & ~x6)));
  assign n3073 = (~n3074 | n3077) & (~x0 | n3075) & (x0 | n3076);
  assign n3074 = ~x0 & ~x6;
  assign n3075 = (~x1 | x2 | x3 | ~x5 | ~x6) & (x1 | x6 | (x2 ? (~x3 ^ x5) : (x3 | x5)));
  assign n3076 = (~x1 | ~x2 | ~x3 | ~x5 | x6) & (x1 | x2 | x3 | x5 | ~x6);
  assign n3077 = (x1 | ~x2 | x3 | x4 | x5) & (~x1 | ~x4 | ((x3 | x5) & (x2 | ~x3 | ~x5)));
  assign z134 = ~n3097 | ~n3092 | n3089 | n3079 | n3086;
  assign n3079 = ~x0 & (n3080 | n3083);
  assign n3080 = ~x3 & ((~x2 & ~n3081) | (n1133 & ~n3082));
  assign n3081 = (x1 | (x4 ? (x6 | x7) : (~x6 | ~x7))) & (x4 | ((x6 | x7 | ~x1 | x5) & (~x5 | ~x6 | ~x7)));
  assign n3082 = x5 ? (x4 ? (~x6 | x7) : (x6 | ~x7)) : (~x6 | ~x7);
  assign n3083 = x3 & ((n530 & n3084) | (x2 & ~n3085));
  assign n3084 = ~x4 & ~x1 & ~x2;
  assign n3085 = (x1 | x4 | ~x5 | x6 | ~x7) & (~x6 | ((~x1 | ~x4 | x5 | x7) & (x1 | ((x5 | ~x7) & (~x4 | ~x5 | x7)))));
  assign n3086 = n841 & ((~n1198 & ~n3087) | (n597 & ~n3088));
  assign n3087 = (~x2 | ~x3 | ~x4 | x7) & (x2 | (x3 ? (x4 | ~x7) : (~x4 | x7)));
  assign n3088 = (x5 | x7 | ~x2 | x3) & (x2 | ~x3 | (~x5 ^ x7));
  assign n3089 = ~n1097 & ((n733 & n3090) | (~x1 & ~n3091));
  assign n3090 = ~x7 & x3 & x4;
  assign n3091 = (x0 | ~x2 | x3 | ~x4 | x7) & (~x0 | x4 | ~x7 | (~x2 ^ ~x3));
  assign n3092 = ~n3096 & (x2 | (n3094 & (~n543 | ~n3093)));
  assign n3093 = ~x5 & (x3 ? (~x4 & x6) : (x4 & ~x6));
  assign n3094 = (n1408 | n3095) & (~n559 | ~n661);
  assign n3095 = (x0 | x1 | ~x3 | x5) & (~x0 | ~x1 | x3 | ~x5);
  assign n3096 = n1269 & n1228;
  assign n3097 = (n643 | n3099) & (n3098 | n3102);
  assign n3098 = x4 ? (~x6 | ~x7) : (x6 | x7);
  assign n3099 = n3101 & (x2 ? (~n543 | n856) : n3100);
  assign n3100 = (x1 | ((~x0 | (x3 ? (~x4 | x5) : (x4 | ~x5))) & (x4 | x5 | x0 | x3))) & (x0 | ~x1 | (x3 ? (~x4 | x5) : ~x5));
  assign n3101 = x0 ? (x4 | (x1 ? (x2 | x5) : (~x2 | ~x5))) : (x1 | ~x4 | (~x2 ^ x5));
  assign n3102 = (~x0 | x5 | (x2 ? x1 : x3)) & (x1 | ~x5 | (~x2 ^ x3)) & (x0 | ((~x3 | ~x5) & (~x1 | (~x5 & (~x2 | ~x3)))));
  assign z135 = ~n3115 | n3112 | n3110 | n3104 | n3108;
  assign n3104 = x7 & (n3106 | (~n1198 & ~n3105));
  assign n3105 = (x0 | ~x1 | ~x2 | (~x3 ^ x4)) & (x1 | ((~x3 | ~x4 | x0 | ~x2) & (~x0 | (x2 ? (x3 | x4) : (~x3 | ~x4)))));
  assign n3106 = x5 & ((n560 & n744) | (~x0 & ~n3107));
  assign n3107 = (x1 | ~x2 | x3 | x4 | ~x6) & (x2 | ((x3 | x4 | x6) & (~x6 | (x1 ? (~x3 ^ x4) : (~x3 | ~x4)))));
  assign n3108 = n1429 & ((n560 & n1141) | (~x0 & ~n3109));
  assign n3109 = x2 ? (~x6 | (x1 ? (x3 | x4) : (~x3 ^ x4))) : (x1 ? (x3 ? (~x4 | ~x6) : (x4 | x6)) : (x3 ? (x4 | x6) : (~x4 ^ x6)));
  assign n3110 = ~x1 & ((n530 & n549) | (~x3 & ~n3111));
  assign n3111 = (x0 | x2 | ~x6 | (~x5 ^ x7)) & (~x2 | ((x6 | ~x7 | x0 | x5) & (x7 | (x0 ? (~x5 ^ ~x6) : (~x5 | x6)))));
  assign n3112 = ~x2 & (x3 ? ~n3113 : ~n3114);
  assign n3113 = x1 ? ((x5 | x7 | ~x0 | x4) & (~x5 | ~x7 | x0 | ~x4)) : (x0 ? (x4 ? (x5 | x7) : (~x5 | ~x7)) : (~x5 ^ x7));
  assign n3114 = ((x0 ? (x1 | x4) : (~x1 | ~x4)) | (~x5 ^ x7)) & (~x0 | ~x5 | ~x7 | (~x1 & ~x4));
  assign n3115 = ~n3116 & ~n3118 & (n1008 | (~n3121 & ~n3122));
  assign n3116 = x1 & ((n942 & n600) | (n825 & ~n3117));
  assign n3117 = (x2 | x5 | x6 | ~x7) & (x7 | (x2 ? (~x5 ^ ~x6) : (~x5 | x6)));
  assign n3118 = x2 & ((~x1 & ~n3119) | (n543 & ~n3120));
  assign n3119 = (~x7 | (x3 ^ ~x4) | (x0 ^ ~x5)) & (~x3 | x7 | (x0 ? (x4 | ~x5) : (~x4 | x5)));
  assign n3120 = (~x3 | ~x4 | x5 | ~x7) & (x3 | (x4 ? (x5 | x7) : (~x5 | ~x7)));
  assign n3121 = n1044 & ((n543 & n2359) | (~n2208 & n2337));
  assign n3122 = n1209 & n745;
  assign z136 = n3124 | ~n3129 | ~n3136 | (~n643 & ~n3127);
  assign n3124 = ~n640 & ((~n3125 & n2742) | (~x0 & ~n3126));
  assign n3125 = x2 ? (~x3 | x5) : (~x3 ^ ~x5);
  assign n3126 = x4 ? ((~x2 & ~x5) | (x1 ^ ~x3)) : (x5 | (x1 ? (x2 | ~x3) : (~x2 | x3)));
  assign n3127 = x2 ? (~x4 | (n1119 & ~n1600)) : n3128;
  assign n3128 = x1 ? ((~x4 | ~x5 | x0 | ~x3) & (~x0 | x3 | (~x4 ^ x5))) : ((~x3 | x4 | x5) & (~x4 | ~x5 | x0 | x3));
  assign n3129 = ~n3130 & (~x6 | (~n3132 & (~n570 | n3135)));
  assign n3130 = x2 & ((n559 & n712) | (~x4 & ~n3131));
  assign n3131 = (x1 | (~x0 & ~x5) | (~x3 ^ x6)) & (x0 | ~x1 | (x3 ? ~x6 : (~x5 | x6)));
  assign n3132 = ~x2 & ((~n3133 & ~n3134) | (n689 & ~n1591));
  assign n3133 = x3 ? (~x4 | x5) : (x4 | ~x5);
  assign n3134 = x0 ? (x1 | ~x7) : (~x1 | x7);
  assign n3135 = (x0 | x3 | ~x4 | x5 | x7) & (~x0 | ~x3 | x4 | ~x5 | ~x7);
  assign n3136 = ~n3137 & (x6 | (~n3140 & (~n746 | ~n1598)));
  assign n3137 = ~x2 & (x1 ? ~n3139 : ~n3138);
  assign n3138 = x3 ? (x6 | (~x4 ^ x5)) : (x0 ? (x6 | (x4 & ~x5)) : (~x6 | (~x4 ^ x5)));
  assign n3139 = (x4 | ~x6 | ((x3 | x5) & (x0 | ~x3 | ~x5))) & (x6 | ((x0 | x3 | ~x4 | x5) & (~x0 | (x3 ? (x4 | x5) : (~x4 | ~x5)))));
  assign n3140 = ~x1 & ((n547 & n809) | (x2 & ~n3141));
  assign n3141 = (~x0 | x7 | (x3 ? (~x4 | ~x5) : (x4 | x5))) & (x0 | ~x3 | x4 | x5 | ~x7);
  assign z137 = n3148 | (x2 ? (~n3143 | ~n3158) : ~n3154);
  assign n3143 = n3145 & (x1 | (~n3144 & (~n943 | ~n2094)));
  assign n3144 = n1310 & ((x3 & ~x4 & x6 & ~x7) | (~x3 & (x4 ? (x6 ^ ~x7) : (~x6 & x7))));
  assign n3145 = (n2967 | n3146) & (n643 | n3147);
  assign n3146 = x3 ? (~x5 | ~x7) : (x5 | x7);
  assign n3147 = (x0 | ~x1 | x3 | x4 | x5) & (~x0 | x1 | ~x3 | ~x4 | ~x5);
  assign n3148 = ~x2 & (x1 ? ~n3149 : (n3150 | n3153));
  assign n3149 = (~x4 | ~n1070 | x0 | ~x3) & (~x0 | x3 | x4 | ~n658);
  assign n3150 = n3151 & ((n1857 & n566) | (~x4 & ~n3152));
  assign n3151 = ~x3 & x5;
  assign n3152 = x0 ? (~x6 ^ ~x7) : (x6 ^ ~x7);
  assign n3153 = ~x5 & n536 & (n1395 | n2584);
  assign n3154 = ~n3156 & (x3 ? (x5 | n3157) : n3155);
  assign n3155 = (~x1 | (x0 ? (~x5 | (~x4 ^ x7)) : (x5 | x7))) & (x1 | ~x4 | ~x5 | ~x7) & (x0 | x5 | ((~x4 | x7) & (x1 | x4 | ~x7)));
  assign n3156 = ~n1218 & ((x0 & ~x3 & ~x5) | (x5 & (~n1682 | (~x0 & x3))));
  assign n3157 = (x4 | x7 | ~x0 | ~x1) & (x0 | (~x4 ^ x7));
  assign n3158 = n3160 & (x0 | n3159);
  assign n3159 = (~x1 | ~x3 | x4 | x5 | x7) & (~x5 | ((x3 | ~x4 | ~x7) & (x1 | ((~x4 | ~x7) & (x3 | x4 | x7)))));
  assign n3160 = (x0 | ~x1 | n1337) & (x1 | ((~x3 | n1337) & (~x0 | (n1337 & (~x3 | ~n2209)))));
  assign z139 = n638 | ~n648 | n3163 | (~x3 & ~n3162);
  assign n3162 = ~n636 & (x6 | (~n633 & (~n635 | ~n837)));
  assign n3163 = ~n643 & (~n644 | n645 | (n1268 & n733));
  assign z140 = ~n666 | n3165 | (n686 & ~n3168);
  assign n3165 = ~x2 & (n680 | n3166);
  assign n3166 = x4 & (n679 | (~x7 & ~n3167));
  assign n3167 = (~x0 | ((x1 | ~x3 | ~x5 | x6) & (~x1 | x3 | x5 | ~x6))) & (x0 | ~x1 | ~x3 | ~x5 | ~x6) & (x5 | x6 | x1 | x3);
  assign n3168 = ((~x4 ^ ~x7) | ((x1 | ~x6) & (x0 | ~x1 | x6))) & (x4 | ~x7 | ((x1 | x6) & (x0 | ~x1 | ~x6)));
  assign z141 = n3170 | n3177 | ~n3182 | (~x3 & ~n3172);
  assign n3170 = ~n697 & (x0 ? (n1358 & n1188) : ~n3171);
  assign n3171 = (x5 | x6 | x3 | x4) & (~x3 | ((~x1 | ~x4 | ~x5 | x6) & (x5 | ~x6 | x1 | x4)));
  assign n3172 = ~n3173 & ~n3174 & ~n3175 & (~n733 | ~n993);
  assign n3173 = n597 & ((n841 & n2475) | (n543 & n2477));
  assign n3174 = ~x2 & ((n566 & n978) | (x0 & ~n1113));
  assign n3175 = n530 & n3176;
  assign n3176 = x4 & ~x0 & x2;
  assign n3177 = ~x2 & (~n3179 | (~x4 & ~n3178));
  assign n3178 = (~x0 | x1 | ~x3 | ~x5 | x6) & (x0 | ~x1 | (x3 ? (~x5 | x6) : (x5 | ~x6)));
  assign n3179 = ~n3180 & ~n3181 & (~n1358 | ~n699);
  assign n3180 = x3 & x5 & ((~x1 & x6) | (~x0 & (~x1 | x6)));
  assign n3181 = ~x3 & (x0 | ~x1) & (x5 ^ x6);
  assign n3182 = (~n664 | ~n830) & (~x2 | n3183);
  assign n3183 = (x0 | n711) & (x1 | (n711 & (~x0 | x4 | ~n1520)));
  assign z142 = ~n3199 | ~n3195 | ~n3189 | n3185 | n3187;
  assign n3185 = n841 & (x2 ? (n1392 & n658) : ~n3186);
  assign n3186 = (x3 | x4 | x5 | x6 | ~x7) & (~x6 | ((~x3 | ~x4 | ~x5 | x7) & (x3 | (x4 ? (~x5 | ~x7) : (x5 | x7)))));
  assign n3187 = ~n714 & ~n3188;
  assign n3188 = (x1 | ((x2 | x3 | ~x6) & (~x0 | ~x2 | ~x3 | x6))) & (x0 | (x1 ? (~x3 | x6) : (x3 | ~x6)));
  assign n3189 = ~n3191 & ~n3193 & (x2 | n726 | n3190);
  assign n3190 = x0 ? (~x4 | x5) : (x4 | ~x5);
  assign n3191 = ~x0 & ((n943 & n1288) | (n942 & n3192));
  assign n3192 = ~x4 & ~x1 & ~x3;
  assign n3193 = ~n1116 & ((n543 & n1556) | (x0 & n3194));
  assign n3194 = x4 & ~x1 & x3;
  assign n3195 = ~n739 & ~n3196 & ~n3197 & (~n626 | ~n745);
  assign n3196 = n746 & n960;
  assign n3197 = ~n2830 & ~n3198;
  assign n3198 = (~x0 | x1 | ~x2 | ~x4 | ~x6) & (x0 | ((~x1 | x2 | ~x4 | ~x6) & (x1 | ~x2 | x4 | x6)));
  assign n3199 = (n524 | n3200) & (x4 | n3201);
  assign n3200 = (x3 | x6 | ((~x1 | x2) & (x0 | (~x1 & x2)))) & (x0 | ~x3 | ~x6 | (x1 & ~x2));
  assign n3201 = (~x0 | x1 | x2 | ~x3 | x6) & (x3 | ~x6 | (x0 ? (x1 ^ ~x2) : (~x1 | ~x2)));
  assign z143 = n3209 | n3213 | (x7 ? ~n3203 : ~n3216);
  assign n3203 = n3206 & (x5 | (x0 & n3204) | (~x0 & ~n3205));
  assign n3204 = (~x3 | x4 | x6 | ~x1 | x2) & (x1 | ~x2 | x3 | ~x4 | ~x6);
  assign n3205 = x1 & ~x3 & (x2 ? (~x4 & ~x6) : (x4 & x6));
  assign n3206 = (n1353 | n3208) & (~x5 | ~n653 | n3207);
  assign n3207 = (x4 | x6 | ~x1 | x2) & (~x4 | ~x6 | x1 | ~x2);
  assign n3208 = (x0 | x1 | ~x2 | ~x3 | ~x5) & (x5 | ((x0 | ~x1 | x2 | ~x3) & (~x0 | (x1 ? (x2 | x3) : (~x2 | ~x3)))));
  assign n3209 = ~x4 & (~n3211 | (~x2 & ~n3210));
  assign n3210 = ((~x0 ^ x1) | (x3 ? (~x5 | x7) : (x5 | ~x7))) & (x3 | ~x5 | x7 | (~x0 ^ ~x1));
  assign n3211 = ~n3212 & (~n746 | ~n2476) & (~n626 | ~n2477);
  assign n3212 = x2 & ((x0 & ~x1 & x5 & ~x7) | (~x0 & (x1 ? (x5 & ~x7) : (~x5 & x7))));
  assign n3213 = x4 & (n3214 | n3215 | (n733 & n1545));
  assign n3214 = ~x1 & ((x2 & ~n599) | (x0 & n2551));
  assign n3215 = ~n765 & ((~x0 & (x2 ? x1 : x3)) | (~x2 & ~x3 & (x0 | ~x1)));
  assign n3216 = (~n733 | ~n3217) & (~n2925 | n3218);
  assign n3217 = ~x6 & ~x5 & ~x3 & x4;
  assign n3218 = (x0 & x5 & (x2 | x3)) | (~x2 & ~x3 & ~x5) | (~x0 & (~x5 | (~x2 & ~x3)));
  assign z144 = n3220 | n3224 | ~n3228 | (~x0 & ~n3227);
  assign n3220 = ~x2 & (n938 | n3221 | (n699 & n728));
  assign n3221 = ~x3 & ((n943 & n3222) | (n1310 & ~n3223));
  assign n3222 = x4 & x0 & ~x1;
  assign n3223 = (~x4 | x6 | x7) & (~x6 | ~x7 | ~x1 | x4);
  assign n3224 = ~x1 & ((x0 & ~n3225) | (n3074 & ~n3226));
  assign n3225 = x2 ? ((~x6 | ~x7 | ~x3 | ~x5) & (x6 | x7 | x3 | x5)) : (x6 | (x3 ? (~x5 ^ ~x7) : (~x5 ^ x7)));
  assign n3226 = (~x2 | x3 | ~x5 | x7) & (x2 | ((x5 | ~x7) & (~x3 | ~x5 | x7)));
  assign n3227 = (~x1 | ((~x5 | ~x6 | x2 | x3) & (~x2 | ~x3 | x5))) & (x5 | ~x6 | ~x2 | ~x3) & (x1 | ((~x2 | ~x3 | ~x5 | x6) & (x5 | ~x6 | x2 | x3)));
  assign n3228 = ~n3235 & ~n3233 & ~n3231 & ~n3229 & ~n3230;
  assign n3229 = ~n2227 & ((~x0 & ~x5 & (x1 ^ x6)) | (x5 & x6 & x0 & ~x1));
  assign n3230 = ~n753 & ((n653 & n548) | (n536 & n550));
  assign n3231 = ~n3232 & n757 & n596;
  assign n3232 = (~x0 | x1 | ~x4 | x6) & (x0 | (x1 ? (~x4 | ~x6) : (x4 | x6)));
  assign n3233 = n2061 & ((n632 & n1051) | (~x1 & ~n3234));
  assign n3234 = x2 ? (~x3 | x6) : (x3 | ~x6);
  assign n3235 = n3236 & (n3237 | (~x2 & ~n765 & ~n1794));
  assign n3236 = x1 & x6;
  assign n3237 = ~x7 & ~x5 & ~x3 & ~x0 & x2;
  assign z145 = n3239 | ~n3242 | ~n3244 | (x2 & ~n3241);
  assign n3239 = ~n643 & ((n731 & n1209) | (x1 & ~n3240));
  assign n3240 = (x0 | (x3 ? x2 : x4)) & (x2 | ((x4 | x5) & (~x0 | x3)));
  assign n3241 = (x0 | x1 | ~x4 | x6) & ((~x3 ^ x4) | ((x1 | x6) & (x0 | ~x1 | ~x6)));
  assign n3242 = ~n3243 & (~n1250 | (~n2315 & (~x1 | ~n1479)));
  assign n3243 = ~n1744 & ((n841 & n1397) | (n530 & n746));
  assign n3244 = (~x2 | n3245) & (x1 | n640 | n3246);
  assign n3245 = (~n592 | ~n866) & (x6 | ~n841 | n3133);
  assign n3246 = (x0 | (x2 ? (x3 | x4) : ~x3)) & (~x2 | x3 | x4 | x5) & (x2 | ((~x3 | x4) & (~x0 | x3 | ~x4)));
  assign z146 = n3248 | n3252 | ~n3256 | (x2 & ~n3255);
  assign n3248 = x5 & (n3249 | (~x3 & n1283 & n3251));
  assign n3249 = x2 & ((n2320 & ~n2017) | (~x6 & ~n3250));
  assign n3250 = (~x0 | x1 | x3 | x4 | x7) & (x0 | ((~x3 | ~x4 | ~x7) & (~x1 | x3 | x4 | x7)));
  assign n3251 = x7 & (x4 ^ x6);
  assign n3252 = ~x5 & ((x1 & ~n3253) | (n570 & ~n3254));
  assign n3253 = (~x3 | x4 | x7 | ~x0 | x2) & (x0 | ((~x4 | ~x7 | x2 | x3) & (~x2 | (x3 ? (~x4 | ~x7) : (x4 | x7)))));
  assign n3254 = (~x3 | ~x4 | ~x7) & (x4 | x7 | ~x0 | x3);
  assign n3255 = (x0 | x1 | x3 | x4 | x7) & (~x7 | (x0 & x1) | (~x3 ^ x4));
  assign n3256 = (x2 | n3257) & (~x2 | ~x5 | ~n841 | n2017);
  assign n3257 = (x0 | ((~x3 | x7) & (x1 | x3 | ~x7))) & (x7 | (x3 ? x1 : (~x0 & (~x1 | x4))));
  assign z147 = n3259 | n3263 | ~n3267 | (n570 & ~n3265);
  assign n3259 = ~x2 & ((n712 & n2402) | (~x3 & ~n3260));
  assign n3260 = (~n527 | n3262) & (~x5 | ~n543 | ~n3261);
  assign n3261 = x6 & (~x4 ^ x7);
  assign n3262 = (x0 | x4 | x5 | ~x7) & (~x0 | ~x4 | (~x5 ^ ~x7));
  assign n3263 = ~x0 & ((n559 & n2135) | (~x4 & ~n3264));
  assign n3264 = (x1 | ~x2 | ~x3 | x5 | x6) & (x3 | ((x1 | x2 | x5 | ~x6) & (~x1 | ~x5 | (~x2 ^ ~x6))));
  assign n3265 = (~n943 | ~n1908) & (~x6 | ~n825 | n3266);
  assign n3266 = x4 ? (~x5 | ~x7) : (x5 | x7);
  assign n3267 = ~n3268 & ~n3270 & n3271 & (n710 | n2099);
  assign n3268 = ~n1532 & ((n3269 & n543) | (n1746 & n841));
  assign n3269 = ~x6 & x3 & ~x5;
  assign n3270 = ~n2528 & ~x5 & n1181;
  assign n3271 = (~n731 | ~n1209) & (~x0 | ~n1556);
  assign z148 = n3273 | ~n3278 | ~n3282 | (n527 & ~n3277);
  assign n3273 = ~x0 & (n3274 | (~x4 & ~n3276));
  assign n3274 = x4 & ((~n2063 & ~n3275) | (n658 & n676));
  assign n3275 = x1 ? (x2 | x3) : (~x2 | ~x3);
  assign n3276 = (~x3 | ~n1070 | x1 | ~x2) & (~x1 | x2 | x3 | ~n1383);
  assign n3277 = ((~x0 ^ ~x2) | (x3 ? (x4 | ~x5) : (~x4 | x5))) & (x3 | x4 | x5 | (~x0 ^ x2));
  assign n3278 = (n1134 | n3280) & (~x6 | (~n3279 & ~n3281));
  assign n3279 = n560 & n1268;
  assign n3280 = (x0 | ~x1 | ~x2 | ~x3 | ~x6) & (~x0 | x2 | x6 | (~x1 ^ x3));
  assign n3281 = ~n823 & ((n1477 & n902) | (n2332 & n596));
  assign n3282 = ~n3283 & (x3 ? n3285 : n3286);
  assign n3283 = n841 & ((x5 & ~n3284) | (~x2 & ~x5 & ~n1850));
  assign n3284 = (x2 | ~x3 | ~x4 | ~x6 | x7) & (~x2 | x3 | x4 | x6 | ~x7);
  assign n3285 = (x4 | ~x5 | x0 | ~x2) & ((~x4 ^ ~x5) | (x0 ? (x1 | ~x2) : x2));
  assign n3286 = (~x4 | x5 | x0 | ~x2) & (x2 | (x1 ^ ~x5) | (x0 ^ x4));
  assign z149 = ~n3293 | ~n3299 | (~x7 & (n3288 | n3291));
  assign n3288 = ~x3 & ((x6 & ~n3289) | (n706 & ~n3290));
  assign n3289 = x0 ? ((~x1 | x2 | ~x4 | x5) & (x1 | ~x2 | x4 | ~x5)) : (x4 | ((x2 | ~x5) & (~x1 | ~x2 | x5)));
  assign n3290 = x0 ? (x1 ? (x2 | x4) : (~x2 | ~x4)) : (x1 | (~x2 ^ x4));
  assign n3291 = x3 & (x4 ? (n543 & ~n2291) : ~n3292);
  assign n3292 = (x0 | ~x1 | ~x2 | ~x5 | x6) & (x5 | ((x0 | x1 | x2 | ~x6) & (~x0 | (x1 ? (x2 | x6) : (~x2 | ~x6)))));
  assign n3293 = ~n3294 & (n1097 | (n3296 & n3297));
  assign n3294 = ~x0 & (x1 ? ~n3295 : ~n2138);
  assign n3295 = x2 ? ((x3 | ~x4 | ~x5 | x6) & (~x3 | x4 | x5 | ~x6)) : (x4 ? (x5 | ~x6) : (x6 | (~x3 ^ ~x5)));
  assign n3296 = x0 ? ((x1 | ~x2 | ~x3 | x4) & (~x1 | x2 | x3 | ~x4)) : ((x1 | x2 | ~x3 | x4) & (~x2 | (x1 ? (~x3 ^ ~x4) : (x3 | ~x4))));
  assign n3297 = (~n733 | ~n2047) & (~x4 | n3298);
  assign n3298 = (x0 | x1 | ~x3 | (~x2 ^ ~x7)) & ((~x2 ^ x7) | (x0 ? (x1 | ~x3) : (~x1 | x3)));
  assign n3299 = ~n3301 & (~x7 | (~n3303 & (~n733 | ~n3300)));
  assign n3300 = ~x6 & x5 & ~x3 & ~x4;
  assign n3301 = x0 & (x1 ? (n704 & n1044) : ~n3302);
  assign n3302 = (x6 | (x2 ? (x3 ? (~x4 | ~x5) : (x4 | x5)) : (x4 | ~x5))) & (~x4 | ~x6 | ((x3 | x5) & (x2 | (x3 & x5))));
  assign n3303 = ~x1 & ((~n2077 & ~n1998) | (n622 & ~n3304));
  assign n3304 = (~x2 | x4 | ~x5 | x6) & (x2 | x5 | (~x4 ^ x6));
  assign z150 = n3318 | n3321 | (x5 ? ~n3306 : ~n3311);
  assign n3306 = x3 ? n3310 : (~n3308 & (x0 | n3307));
  assign n3307 = (x6 | ~x7 | x1 | ~x4) & (~x1 | x4 | (x2 ? x7 : (x6 | ~x7)));
  assign n3308 = n841 & ((n1518 & n1769) | (~n1408 & ~n3309));
  assign n3309 = x2 ^ x7;
  assign n3310 = (x1 | ~n550) & (x0 | ~n548 | (x1 ^ ~x2));
  assign n3311 = ~n3316 & ~n3312 & ~n3314;
  assign n3312 = x2 & ((n550 & n866) | (~x3 & ~n3313));
  assign n3313 = (x1 | x4 | ~x6 | x7) & (x0 | ~x1 | x6 | ~x7);
  assign n3314 = ~n3315 & ((n626 & n859) | (x0 & ~n913));
  assign n3315 = x3 ? (x6 | ~x7) : (~x6 | x7);
  assign n3316 = ~x2 & (~n1594 | (~x0 & ~n3317));
  assign n3317 = (x1 | ((x3 | x4 | ~x6 | x7) & (x6 | ~x7 | ~x3 | ~x4))) & (~x1 | x3 | ~x4 | x6 | ~x7);
  assign n3318 = ~n3319 & ~n3320;
  assign n3319 = x4 ? (~x6 | x7) : (x6 | ~x7);
  assign n3320 = x1 ? ((x3 | ~x5 | ~x0 | x2) & (x0 | ~x3 | (x2 & ~x5))) : ((~x2 | (~x3 ^ x5)) & (x3 | (x5 ? x0 : x2)));
  assign n3321 = ~n640 & (n3323 | ~n3324 | (x0 & ~n3322));
  assign n3322 = (~x1 | x2 | x3 | ~x4 | x5) & (x1 | ((x4 | x5 | x2 | x3) & (~x2 | ~x3 | (x4 & ~x5))));
  assign n3323 = n626 & ((~x2 & ~x3 & x4 & ~x5) | (x2 & x3 & (~x4 | x5)));
  assign n3324 = (n1566 | n3325) & (n1916 | (~n3222 & ~n2449));
  assign n3325 = (x1 | x2 | x4) & (x0 | ~x1 | ~x4);
  assign z151 = ~n3327 | (x1 ? (n3337 | n3338) : ~n3331);
  assign n3327 = ~n3330 & (n640 | (n3329 & (x2 | n3328)));
  assign n3328 = (~x0 | ~x1 | x3 | ~x4 | ~x5) & (x4 | (x0 ? (x1 ? (x3 | x5) : (~x3 | ~x5)) : (~x3 | (~x1 ^ ~x5))));
  assign n3329 = (~x2 | ((x1 | (~x4 ^ ~x5)) & (x0 | ~x4 | ~x5))) & (x4 | (x0 ? (x1 | x5) : (x1 ? x5 : (x2 | ~x5))));
  assign n3330 = ~n2128 & (n1890 | (~x2 & ~n1794));
  assign n3331 = x3 ? n3332 : (n3336 & (x2 | n3335));
  assign n3332 = x2 ? (~n3333 & (~n525 | ~n943)) : n3334;
  assign n3333 = ~x7 & x6 & ~x5 & ~x0 & ~x4;
  assign n3334 = x4 ? (x5 ? (x6 | ~x7) : (~x6 | x7)) : ((x5 | x6 | ~x7) & (~x0 | ~x5 | ~x6 | x7));
  assign n3335 = (x0 | x4 | x5 | ~x7) & (~x0 | ~x4 | ((x6 | x7) & (~x5 | (x6 & x7))));
  assign n3336 = (~x0 | x4 | (x2 ? ~n530 : n1116)) & (~x4 | n1116 | (x0 & ~x2));
  assign n3337 = ~n1116 & ((~x2 & ~x3 & ~x4) | (~x0 & x4 & (~x2 | ~x3)));
  assign n3338 = ~x4 & ((n530 & n1783) | (~x2 & ~n3339));
  assign n3339 = (~x0 | ~x3 | x5 | ~x6 | x7) & (x0 | ((~x3 | x5 | x6 | ~x7) & (x3 | ~x5 | ~x6)));
  assign z152 = n3353 | ~n3356 | (x2 ? ~n3341 : ~n3346);
  assign n3341 = ~n3344 & (x0 | (~n3343 & (~x6 | n3342)));
  assign n3342 = (~x1 | x4 | x7 | (~x3 ^ ~x5)) & (x5 | ~x7 | (~x3 & ~x4));
  assign n3343 = x7 & n706 & (~n1548 | n3192);
  assign n3344 = n841 & (x3 ? (x7 & ~n1198) : ~n3345);
  assign n3345 = (x4 | x5 | ~x6 | x7) & (~x4 | ~x5 | x6 | ~x7);
  assign n3346 = x0 ? (~n3351 & (x5 | n3350)) : n3347;
  assign n3347 = x4 ? (x7 | n3349) : n3348;
  assign n3348 = (~x1 | x3 | (x5 ? (~x6 | ~x7) : (x6 | x7))) & (~x3 | (x5 ? (x6 | x7) : ((~x6 | x7) & (x1 | x6 | ~x7))));
  assign n3349 = (~x5 | x6) & (~x3 | x5 | ~x6);
  assign n3350 = (x1 | ~x3 | ~x6 | x7) & (x6 | ((x1 | ~x3 | ~x4 | ~x7) & (~x1 | (x3 ? (x4 | ~x7) : (~x4 | x7)))));
  assign n3351 = n551 & (n3352 | (n1300 & n1392));
  assign n3352 = ~x7 & x3 & ~x6;
  assign n3353 = ~n1097 & ((n1044 & ~n3355) | (x3 & ~n3354));
  assign n3354 = x2 ? (x7 | ((x1 | ~x4) & (x0 | (x1 & ~x4)))) : (x4 | ~x7 | (~x0 ^ x1));
  assign n3355 = x0 ? (x4 | x7) : (~x7 | (x1 & ~x4));
  assign n3356 = n3359 & (n823 | n3357) & (~n1044 | n3358);
  assign n3357 = (~x2 | x5 | x7 | (x3 ^ ~x4)) & (~x7 | ((x4 | ~x5 | ~x2 | x3) & (x2 | (x3 ? (~x4 | ~x5) : (x4 | x5)))));
  assign n3358 = (x0 | x4 | ~x5 | x7) & (~x0 | ~x4 | ((~x5 | x7) & (x1 | x5 | ~x7)));
  assign n3359 = (~n1460 | ~n837) & (~n626 | n1546);
  assign z153 = n3370 | ~n3372 | (x2 ? ~n3361 : ~n3365);
  assign n3361 = ~n3362 & (~n661 | ~n817) & (n1097 | n3364);
  assign n3362 = ~x0 & (x6 ? (n681 & ~n1605) : ~n3363);
  assign n3363 = (~x1 | x3 | (x4 ? (~x5 | ~x7) : (x5 | x7))) & (~x3 | ((x4 | ~x5 | x7) & (x5 | ~x7 | x1 | ~x4)));
  assign n3364 = (~x0 | x1 | x3 | x4 | x7) & (x0 | ~x1 | ~x3 | ~x4 | ~x7);
  assign n3365 = x5 ? n3368 : (x0 ? n3366 : n3367);
  assign n3366 = x1 ? (x7 | (x3 ? (x4 | ~x6) : (~x4 | x6))) : (~x4 | ~x7 | (~x3 ^ x6));
  assign n3367 = (x1 | ~x3 | x4 | x6 | ~x7) & (x3 | ((~x4 | ~x6 | x7) & (~x1 | x4 | (~x6 ^ ~x7))));
  assign n3368 = (~n550 | ~n699) & (x1 | n3369);
  assign n3369 = (x0 | ~x3 | ~x6 | (~x4 ^ x7)) & (x6 | (x0 ? (x3 ? (x4 | x7) : (~x4 | ~x7)) : (x3 | (~x4 ^ x7))));
  assign n3370 = ~x2 & ((n548 & n699) | (~x1 & ~n3371));
  assign n3371 = x0 ? ((x3 | ~x4 | ~x6 | x7) & (~x3 | x4 | x6 | ~x7)) : ((~x3 | x4 | x6 | x7) & (x3 | (x4 ? (x6 | ~x7) : (~x6 | x7))));
  assign n3372 = ~n3376 & n3378 & (~x2 | (~n3373 & n3375));
  assign n3373 = ~x1 & ~n3374;
  assign n3374 = (x0 | x3 | ((~x4 | x6 | ~x7) & (~x6 | x7))) & (~x3 | x4 | ((x6 | ~x7) & (~x0 | ~x6 | x7)));
  assign n3375 = (~n699 | ~n1585) & (n671 | n1338);
  assign n3376 = ~n640 & (n3377 | (~x2 & (n936 | ~n1327)));
  assign n3377 = x4 & x3 & x2 & ~x0 & ~x1;
  assign n3378 = (x4 | n1143 | x0 | ~x1) & (~x0 | ~x4 | n2499);
  assign z154 = n3389 | ~n3391 | (x3 ? ~n3380 : ~n3384);
  assign n3380 = x1 ? n3381 : (x4 ? n3383 : n3382);
  assign n3381 = (~x4 | ~n978 | x0 | ~x2) & (~x0 | x2 | x4 | ~n951);
  assign n3382 = (x7 | ((x5 | x6 | ~x0 | x2) & (x0 | (x2 ? (x5 | x6) : (~x5 | ~x6))))) & (~x0 | ~x6 | ~x7 | (~x2 ^ ~x5));
  assign n3383 = (~x0 | x2 | x5 | x6 | ~x7) & (x0 | (x2 ? (x5 | (~x6 ^ x7)) : (~x5 | (~x6 ^ ~x7))));
  assign n3384 = (x1 & n3387) | (~n3385 & ~n3386 & ~x1 & ~n2260);
  assign n3385 = n778 & ((~x0 & x4 & ~x5 & x7) | (x0 & x5 & (x4 ^ x7)));
  assign n3386 = ~n643 & ((n681 & n1181) | (n1121 & n995));
  assign n3387 = x5 ? (~n1181 | (~n1395 & ~n2584)) : n3388;
  assign n3388 = (~x4 | x6 | x7 | ~x0 | x2) & ((~x4 ^ ~x7) | (x0 ? (x2 | ~x6) : (~x2 | x6)));
  assign n3389 = ~n671 & ~n3390;
  assign n3390 = (~x0 | x1 | x2 | ~x3 | ~x5) & (x0 | ((~x1 | (x2 ? (x3 | ~x5) : ~x3)) & (x2 | ~x3 | x5) & (x1 | ~x2 | (~x3 ^ ~x5))));
  assign n3391 = ~n3397 & (n1218 | n3392) & (x3 | n3393);
  assign n3392 = x0 ? ((~x1 | x2 | x3 | ~x5) & (x1 | (x3 ? ~x2 : x5))) : ((~x1 | ~x2 | ~x3 | x5) & (x3 | ~x5 | x1 | x2));
  assign n3393 = (n3395 | ~n3396) & (x4 | n3309 | n3394);
  assign n3394 = x0 ? (x1 | ~x5) : (~x1 | x5);
  assign n3395 = (x2 | x5) & (x1 | ~x2 | ~x5);
  assign n3396 = ~x7 & ~x0 & x4;
  assign n3397 = ~n1090 & n742 & x7 & n774;
  assign z155 = n3404 | ~n3411 | (x2 ? ~n3406 : ~n3399);
  assign n3399 = x0 ? n3400 : (~n3403 & (x1 | n3402));
  assign n3400 = (~x6 | n3401) & (x4 | x6 | n765 | ~n1317);
  assign n3401 = x1 ? ((x3 | ~x4 | ~x5 | ~x7) & (~x3 | x4 | x5 | x7)) : (x7 | (x3 ? (~x4 | x5) : (x4 | ~x5)));
  assign n3402 = (x3 | ~x4 | x5 | ~x6 | x7) & (x6 | ((x3 | x4 | x5 | ~x7) & (~x3 | (x4 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n3403 = n1070 & n945;
  assign n3404 = ~x5 & ((n743 & n761) | (x6 & ~n3405));
  assign n3405 = (x0 | ~x1 | ~x4 | (~x2 ^ ~x3)) & (x1 | ((~x3 | ~x4 | x0 | x2) & (~x0 | x3 | (~x2 ^ ~x4))));
  assign n3406 = ~n3407 & (~n661 | ~n1626) & (n1008 | n3410);
  assign n3407 = ~x0 & ((~n1763 & ~n3409) | (n942 & n3408));
  assign n3408 = x4 & x1 & ~x3;
  assign n3409 = (x6 | x7 | x4 | x5) & (~x6 | ~x7 | ~x4 | ~x5);
  assign n3410 = (~x0 | x1 | ~x3 | x4 | ~x6) & (x0 | ((~x1 | ~x3 | ~x4 | x6) & (x4 | ~x6 | x1 | x3)));
  assign n3411 = ~n3412 & ~n3415 & n3417 & (x0 | n3414);
  assign n3412 = n706 & ~n3413;
  assign n3413 = (x0 | ~x1 | x2 | x3 | ~x4) & (x1 | (x0 ? (x2 ? (~x3 ^ x4) : (x3 | x4)) : (x2 ? (x3 | x4) : (~x3 | ~x4))));
  assign n3414 = (x1 | ~x2 | x3 | ~x4 | ~x5) & (~x3 | x4 | (x1 ? (x2 ^ ~x5) : (x2 | x5)));
  assign n3415 = ~n2259 & (n829 | n3416);
  assign n3416 = (x1 ^ x3) & (~x0 ^ ~x2);
  assign n3417 = (~n560 | ~n959) & (n1920 | n1036);
  assign z156 = ~n3438 | ~n3429 | n3426 | n3419 | n3422;
  assign n3419 = ~n1408 & (x1 ? ~n3421 : ~n3420);
  assign n3420 = (x0 | ~x2 | ~x3 | x5 | ~x7) & ((x0 ? (~x2 | x3) : (x2 | ~x3)) | (~x5 ^ ~x7));
  assign n3421 = (x5 | ~x7 | x2 | x3) & (x0 | (x2 ? (~x3 | x7) : (x3 | ~x5)));
  assign n3422 = ~x0 & (x1 ? ~n3424 : (n3423 | n3425));
  assign n3423 = ~x6 & x5 & ~x4 & ~x2 & ~x3;
  assign n3424 = (x2 | ~x3 | ~x4 | x5 | ~x6) & (~x2 | x3 | x4 | ~x5 | x6);
  assign n3425 = x2 & ((~x3 & x4 & x6) | (x3 & ~x4 & x5 & ~x6));
  assign n3426 = x1 & (n3428 | (~x5 & n742 & ~n3427));
  assign n3427 = x3 ? (~x6 | ~x7) : (x6 | x7);
  assign n3428 = ~x2 & (x0 ? (~x3 & n1857) : (x3 & n530));
  assign n3429 = ~n3433 & (~n841 | (~n3430 & ~n3432 & n3437));
  assign n3430 = ~n647 & ~x7 & n3431;
  assign n3431 = x2 & ~x6;
  assign n3432 = x6 & x7 & n1518 & (~x3 | n1301);
  assign n3433 = ~x1 & ((n3435 & n3436) | (n3434 & n1070));
  assign n3434 = ~x3 & x0 & x2;
  assign n3435 = ~x7 & (x2 ^ x5);
  assign n3436 = ~x6 & ~x0 & x3;
  assign n3437 = (~x2 | ~x3 | ~x4 | ~x6) & (x2 | x4 | x6 | (~x3 & x5));
  assign n3438 = ~n3439 & (x0 | (~x1 & n3443) | (x1 & n3442));
  assign n3439 = ~n643 & (x2 ? ~n3441 : ~n3440);
  assign n3440 = (x3 | ((~x0 | ~x5 | (~x1 ^ ~x4)) & (x1 | ~x4 | (x0 & x5)))) & (~x3 | ~x4 | ~x0 | x1) & (~x1 | x4 | ((~x3 | x5) & (x0 | (~x3 & x5))));
  assign n3441 = (x0 | ~x1 | x3 | ~x4) & (x1 | (x0 ? (~x3 | x4) : (x3 ? (~x4 | ~x5) : x4)));
  assign n3442 = (~x2 | ~x3 | x4 | ~n530) & (x2 | x3 | ~x4 | ~n813);
  assign n3443 = (~n813 | ~n1780) & (~n572 | n3444);
  assign n3444 = (x5 | ~x6 | ~x3 | x4) & (x3 | (x4 ? (~x5 | ~x6) : (x5 | x6)));
  assign z157 = n3454 | ~n3459 | (x2 & (~n3446 | ~n3451));
  assign n3446 = x4 ? n3449 : (~n3448 & (x1 | n3447));
  assign n3447 = (~x0 | ~x3 | x5 | x6 | ~x7) & (x7 | ((x0 | ~x3 | ~x5 | x6) & (~x6 | (x0 ? (x3 ^ ~x5) : (x3 | x5)))));
  assign n3448 = n543 & ((~x3 & ~x5 & x6 & x7) | (x3 & ~x6 & (x5 ^ ~x7)));
  assign n3449 = (~n813 | ~n712) & (~n653 | n3450);
  assign n3450 = (x1 | ~x5 | x6 | ~x7) & (~x1 | x5 | (~x6 ^ x7));
  assign n3451 = n3453 & (x0 | n3452);
  assign n3452 = (x1 | x4 | ~x5 | (~x3 ^ ~x7)) & (~x4 | ((x1 | x3 | x5 | ~x7) & (x7 | (x1 ? (~x3 ^ x5) : (~x3 | ~x5)))));
  assign n3453 = (n1580 | n1775) & (~n2296 | ~n661);
  assign n3454 = ~x2 & (n3457 | (~x3 & (n3455 | n3456)));
  assign n3455 = x5 & ((x0 & x4 & x6 & ~x7) | (~x0 & ~x4 & ~x6 & x7));
  assign n3456 = n1477 & ((n543 & n1857) | (n1300 & n841));
  assign n3457 = x3 & ((n657 & n978) | (~x1 & ~n3458));
  assign n3458 = (~x0 | ((~x6 | ~x7 | ~x4 | ~x5) & (x6 | x7 | x4 | x5))) & (x0 | ~x4 | x5 | ~x6 | ~x7);
  assign n3459 = ~n3460 & ~n3462 & (x2 | (~n3465 & n3467));
  assign n3460 = ~n640 & ((n837 & n1311) | (~x0 & ~n3461));
  assign n3461 = (x1 | x2 | x3 | ~x4 | ~x5) & (~x1 | ((~x4 | ~x5 | ~x2 | ~x3) & (x2 | x4 | (~x3 ^ ~x5))));
  assign n3462 = ~n1218 & (n3463 | n3464);
  assign n3463 = x0 & ((~x1 & x2 & x3 & x5) | (x1 & ~x2 & ~x3 & ~x5));
  assign n3464 = ~x0 & x3 & (x1 ? (~x2 & ~x5) : (x2 ^ x5));
  assign n3465 = ~x1 & ~n3466;
  assign n3466 = (~x0 | x3 | x4 | ~x5 | x7) & (x5 | (x0 & x3) | (~x4 ^ x7));
  assign n3467 = ~n3469 & (~n1234 | ~n2209) & (~n543 | ~n3468);
  assign n3468 = x7 & ~x3 & x4;
  assign n3469 = x0 & ~x1 & x3 & (x4 ^ x7);
  assign z158 = n3471 | ~n3477 | (~n1794 & ~n3474);
  assign n3471 = ~x0 & (x2 ? ~n3472 : ~n3473);
  assign n3472 = x3 ? ((~x5 | x6 | x1 | ~x4) & (x5 | ~x6 | ~x1 | x4)) : (x1 ? (x4 ? (x5 | ~x6) : (~x5 | x6)) : (x5 | (~x4 ^ x6)));
  assign n3473 = (~x5 | (x1 ? (x3 ? (~x4 | ~x6) : (x4 | x6)) : (~x3 | (x4 & x6)))) & (x3 | x5 | ~x6 | (~x1 & x4));
  assign n3474 = x2 ? (x1 | (~n1725 & ~n3476)) : n3475;
  assign n3475 = x1 ? ((x4 | x5 | ~x6 | x7) & (x6 | ~x7 | ~x4 | ~x5)) : (x5 | (x4 ? (~x6 | ~x7) : (x6 | x7)));
  assign n3476 = x4 & ~x7 & (x5 ^ ~x6);
  assign n3477 = n3478 & (x4 ? (~n3485 & ~n3487) : n3481);
  assign n3478 = (n1097 | n3479) & (~n841 | n3480);
  assign n3479 = (x3 | ((x0 | x1 | x2 | ~x4) & (~x0 | (x1 ? x2 : (~x2 | x4))))) & (x0 | ~x3 | (x1 ? (~x2 ^ ~x4) : (~x2 | x4)));
  assign n3480 = x3 ? ((~x2 | ((x5 | ~x6) & (x4 | ~x5 | x6))) & (x5 | ((x4 | ~x6) & (x2 | ~x4 | x6)))) : (~x5 | (x4 ? x6 : x2));
  assign n3481 = (n1097 | n3482 | ~n3483) & (n1008 | n3484);
  assign n3482 = x1 ? (~x2 | ~x3) : (x2 | x3);
  assign n3483 = ~x0 & x7;
  assign n3484 = (~x0 | x1 | x2 | ~x3 | x6) & (x0 | ~x2 | x3 | (~x1 ^ ~x6));
  assign n3485 = ~x1 & ((n549 & n951) | (n702 & ~n3486));
  assign n3486 = x0 ? (x2 | ~x3) : (~x2 | x3);
  assign n3487 = n3488 & ((n750 & n596) | (~x2 & n2980));
  assign n3488 = ~x6 & ~x0 & x1;
  assign z159 = ~n3491 | ~n3501 | ~n3506 | (~n2208 & ~n3490);
  assign n3490 = (x0 | ~x2 | x3 | x5 | x6) & (x2 | (x0 ? (x3 ? (x5 | x6) : (~x5 | ~x6)) : (~x6 | (~x3 ^ ~x5))));
  assign n3491 = ~n3494 & n3496 & n3498 & (x0 | n3492);
  assign n3492 = (~n1241 | ~n1498) & (x6 | ~n1467 | ~n3493);
  assign n3493 = x7 & (x2 ? (x3 & x4) : (~x3 & ~x4));
  assign n3494 = ~n2291 & ~n3495;
  assign n3495 = (x3 | x4 | ~x0 | x1) & (x0 | (x1 ? (x3 | ~x4) : (~x3 | x4)));
  assign n3496 = (~n845 | ~n2144) & (~n733 | ~n3497);
  assign n3497 = ~x7 & ~x6 & x3 & ~x4;
  assign n3498 = (n1040 | n3499) & (n1353 | n3500);
  assign n3499 = (x0 | ~x2 | x3 | (~x1 ^ ~x7)) & (x2 | ((x0 | ~x1 | ~x3 | ~x7) & (~x0 | (x1 ? (x3 | ~x7) : x7))));
  assign n3500 = (x0 | x1 | ~x2 | x3 | ~x7) & (~x0 | x2 | (x1 ? (x3 | x7) : (~x3 | ~x7)));
  assign n3501 = ~n3503 & (~x2 | (~n3502 & (~n1358 | ~n661)));
  assign n3502 = x3 & (x0 ? (~x1 & ~n1040) : (x1 & ~n1100));
  assign n3503 = ~n1097 & ((n1181 & n3505) | (x2 & ~n3504));
  assign n3504 = x0 ? (x1 | (x3 ? (x4 | x7) : (~x4 | ~x7))) : (~x1 | ~x3 | (~x4 ^ x7));
  assign n3505 = ~x3 & ~x7 & (~x1 ^ ~x4);
  assign n3506 = ~n3508 & (n640 | (~n3279 & (x0 | n3507)));
  assign n3507 = (x1 | x2 | ~x3 | ~x4 | x5) & (~x5 | ((x3 | x4 | ~x1 | ~x2) & (x1 | (x2 ? (~x3 | ~x4) : (x3 | x4)))));
  assign n3508 = ~n643 & ((n543 & n3509) | (~x1 & ~n3510));
  assign n3509 = ~x5 & ~x2 & x4;
  assign n3510 = (x0 | x2 | ~x3 | x4 | x5) & (~x2 | ((~x0 | (x3 ? (~x4 | x5) : (x4 | ~x5))) & (x4 | ~x5 | x0 | ~x3)));
  assign z160 = n3523 | ~n3525 | (x3 ? ~n3512 : ~n3518);
  assign n3512 = ~n3513 & ~n3516 & (~n1209 | ~n830);
  assign n3513 = ~x0 & (x2 ? ~n3514 : ~n3515);
  assign n3514 = (x1 | ~x4 | ~x5 | x6 | x7) & (~x6 | ((x1 | ~x4 | x5 | x7) & (~x1 | x4 | (~x5 ^ ~x7))));
  assign n3515 = (x1 | x4 | x5 | x6 | ~x7) & (~x1 | ~x5 | (x4 ? (x6 | ~x7) : (~x6 | x7)));
  assign n3516 = ~n1100 & ((n572 & n841) | (n543 & n3517));
  assign n3517 = x2 & ~x7;
  assign n3518 = ~n3521 & (n1198 | n3519) & (~n551 | n3520);
  assign n3519 = (~x4 | ((x0 | x1 | ~x2 | ~x7) & (~x0 | (x1 ? (x2 | ~x7) : (~x2 | x7))))) & (x0 | ((x1 | x2 | x7) & (x4 | ~x7 | ~x1 | ~x2)));
  assign n3520 = (x0 | ~x2 | x4 | x6 | ~x7) & (~x0 | ~x4 | ~x6 | (~x2 ^ ~x7));
  assign n3521 = n3522 & ((n525 & n1857) | (~x0 & ~n1850));
  assign n3522 = ~x5 & x1 & ~x2;
  assign n3523 = ~n1097 & (x3 ? (~n586 & ~n3309) : ~n3524);
  assign n3524 = (x0 | x1 | ~x2 | x4 | x7) & (x2 | ((x0 | ~x7 | (~x1 ^ x4)) & (~x0 | ~x1 | x4 | x7)));
  assign n3525 = ~n3526 & (n1205 | n3528) & (~n841 | n3529);
  assign n3526 = ~x0 & (~n3527 | (n772 & ~n3088));
  assign n3527 = (~x1 | x2 | (x3 ? (x5 | ~x7) : (~x5 | x7))) & (~x2 | ((x5 | x7 | ~x1 | x3) & (~x5 | ~x7 | x1 | ~x3)));
  assign n3528 = x1 ? ((x4 | x5 | ~x0 | x2) & (~x4 | ~x5 | x0 | ~x2)) : (x0 ? (x2 ? (x4 | ~x5) : (~x4 | x5)) : (x4 | (~x2 ^ x5)));
  assign n3529 = ((x3 ? (~x4 | ~x7) : (x4 | x7)) | (x2 ^ ~x5)) & (~x2 | ~x3 | ~x4 | ~x5 | x7) & (x5 | ~x7 | x2 | x4);
  assign z161 = ~n3550 | ~n3542 | n3539 | n3531 | n3534;
  assign n3531 = x1 & (n2581 | n3532);
  assign n3532 = ~x0 & ((n530 & n1556) | (x4 & ~n3533));
  assign n3533 = (x2 | x3 | x5 | ~x6 | ~x7) & (~x3 | ((x6 | ~x7 | x2 | x5) & (~x2 | ~x5 | (~x6 ^ ~x7))));
  assign n3534 = ~x1 & (n3535 | n3537 | (n547 & n845));
  assign n3535 = x2 & (x0 ? (n828 & n978) : ~n3536);
  assign n3536 = (~x3 | ~x4 | ~x5 | x6 | ~x7) & (x3 | x4 | x5 | ~x6 | x7);
  assign n3537 = ~n640 & ((n639 & n995) | (~x0 & ~n3538));
  assign n3538 = (~x4 | ~x5 | ~x2 | x3) & (x4 | x5 | x2 | ~x3);
  assign n3539 = ~n643 & (~n3540 | (n626 & ~n1150));
  assign n3540 = (n968 | n3541) & (~n1287 | ~n837);
  assign n3541 = (x0 | ~x1 | ~x3 | x4) & (x3 | ~x4 | ~x0 | x1);
  assign n3542 = n3549 & ~n3548 & ~n3547 & ~n3543 & ~n3545;
  assign n3543 = ~x1 & ~n3544;
  assign n3544 = (x0 | x2 | x3 | ~x4 | ~x6) & (~x3 | x6 | (x0 ? (~x2 | ~x4) : (~x2 ^ x4)));
  assign n3545 = ~n714 & ~n3546;
  assign n3546 = (x0 | ~x1 | ~x2 | ~x3 | ~x6) & (~x0 | x2 | x3 | (~x1 ^ ~x6));
  assign n3547 = n873 & ((n1300 & n1156) | (n1518 & n1857));
  assign n3548 = ~n586 & ~n1011;
  assign n3549 = (~n733 | ~n1203) & (~n1029 | ~n560 | ~n1857);
  assign n3550 = ~n3552 & (~x6 | (~n2875 & ~n3551));
  assign n3551 = n570 & (x0 ? ~n647 : (x5 & ~n1744));
  assign n3552 = ~n1353 & ((~x3 & ~n3554) | (~n3553 & n3555));
  assign n3553 = x0 ? (x5 | ~x7) : (~x5 | x7);
  assign n3554 = x0 ? (x2 | (x1 ? (~x5 | ~x7) : (x5 | x7))) : (~x2 | (x1 ? (~x5 | x7) : (x5 | ~x7)));
  assign n3555 = x3 & ~x1 & ~x2;
  assign z162 = n3564 | ~n3568 | (~x0 & (n3557 | n3560));
  assign n3557 = x1 & (x3 ? ~n3558 : ~n3559);
  assign n3558 = (x2 | ~x4 | ~x5 | ~x6 | x7) & (~x2 | x4 | x5 | x6 | ~x7);
  assign n3559 = (x6 | (x2 ? (~x4 | x7) : (x4 ? ~x7 : (~x5 | x7)))) & (~x2 | x4 | ~x7 | (x5 & ~x6));
  assign n3560 = ~x1 & (n3562 | ~n3563 | (~x4 & ~n3561));
  assign n3561 = (x2 | ~x7 | ((x5 | ~x6) & (x3 | ~x5 | x6))) & (~x2 | ~x3 | ~x5 | x7);
  assign n3562 = x4 & ((~x2 & ~x3 & x6 & ~x7) | (x2 & x7 & (x3 ^ x6)));
  assign n3563 = x2 | ((~x4 | ~n658) & (~x3 | x4 | ~n1769));
  assign n3564 = ~n765 & (~n3566 | (~x0 & ~n3565));
  assign n3565 = (x1 | x2 | x3 | x4 | ~x6) & (~x2 | ((x4 | ~x6 | x1 | ~x3) & (x3 | (x1 ? (~x4 ^ ~x6) : (~x4 | x6)))));
  assign n3566 = ~n3567 & (~n560 | ~n1331) & (x4 | n1036);
  assign n3567 = x4 & ((~x2 & ~x3 & x0 & x1) | (~x0 & x3 & (x1 ^ ~x2)));
  assign n3568 = ~n3569 & (~x0 | (n3574 & (x2 | n3571)));
  assign n3569 = ~n1008 & (x0 ? ~n1057 : ~n3570);
  assign n3570 = (~x1 | x2 | ~x4 | (~x3 ^ x6)) & (~x2 | ((x1 | (x3 ? (~x4 | ~x6) : x4)) & (x4 | ~x6 | ~x1 | ~x3)));
  assign n3571 = ~n3572 & ~n3573 & (~x5 | ~n772 | ~n2674);
  assign n3572 = ~x1 & (x4 ? (~x5 & x7) : (x6 & ~x7));
  assign n3573 = x7 & ~x6 & ~x5 & x1 & ~x4;
  assign n3574 = (n671 | n1065) & (~n3576 | (~n1029 & ~n3575));
  assign n3575 = ~x6 & ~x3 & ~x4;
  assign n3576 = ~x7 & x5 & ~x1 & x2;
  assign z163 = x2 ? (~n3585 | ~n3595) : (~n3578 | ~n3590);
  assign n3578 = ~n3580 & ~n3582 & n3584 & (n3579 | n3394);
  assign n3579 = (x4 | x6 | ~x7) & (~x3 | ~x4 | ~x6 | x7);
  assign n3580 = ~x1 & ((n2857 & n978) | (~x3 & ~n3581));
  assign n3581 = (x0 | x4 | x5 | ~x6 | x7) & (x6 | ((~x0 | ~x4 | ~x5 | x7) & (x0 | x5 | (x4 ^ ~x7))));
  assign n3582 = ~n3583 & (x0 ? n1429 : n526);
  assign n3583 = (x1 | x3 | ~x4 | x6) & (~x1 | ~x3 | x4 | ~x6);
  assign n3584 = (x3 | n990 | ~x0 | ~x1) & (x0 | (x1 ? (x3 | ~n993) : (~x3 | n990)));
  assign n3585 = ~n3588 & (x1 | (n3586 & (n2924 | n3098)));
  assign n3586 = (~n942 | ~n2204) & (n1205 | n3587);
  assign n3587 = (x0 | x4 | ~x5 | ~x6) & (x5 | x6 | ~x0 | ~x4);
  assign n3588 = n543 & (n3589 | (~n877 & ~n3098));
  assign n3589 = x7 & ~x6 & x5 & ~x3 & ~x4;
  assign n3590 = ~n3591 & ~n3592 & ~n3593 & (~n696 | ~n841);
  assign n3591 = ~n1566 & ((~x4 & ~x6 & x0 & x1) | (~x0 & x4 & (x1 ^ x6)));
  assign n3592 = ~n1010 & ((~x5 & x6 & x1 & ~x3) | (~x1 & x5 & (x3 ^ x6)));
  assign n3593 = x6 & ~n3594;
  assign n3594 = (x4 | ~x5 | ~x0 | x1) & (x0 | ~x1 | (x3 ? (~x4 ^ ~x5) : (~x4 | x5)));
  assign n3595 = ~n3596 & (~n592 | ~n866) & (x1 | n3597);
  assign n3596 = ~n1408 & ((x3 & x5 & x0 & ~x1) | (~x0 & (x1 ? (x3 ^ x5) : (~x3 & ~x5))));
  assign n3597 = (x5 | ~x6 | ~x0 | x3) & (x0 | ~x3 | ~x5 | x6) & ((~x0 ^ ~x3) | (x4 ? (~x5 | ~x6) : (x5 | x6)));
  assign z164 = n3608 | ~n3613 | (x2 ? ~n3599 : ~n3603);
  assign n3599 = x0 ? (x1 | n3602) : (x1 ? n3601 : n3600);
  assign n3600 = x3 ? (~x4 | x7 | (~x5 ^ x6)) : (x4 | (x5 ? (x6 | ~x7) : ~x6));
  assign n3601 = (x3 | x4 | ~x5 | ~x6 | x7) & (~x3 | ((x6 | ~x7 | x4 | x5) & (~x4 | ~x6 | (~x5 ^ x7))));
  assign n3602 = (~x3 | x4 | ~x5 | x6) & (~x6 | ((~x3 | (x4 ? (~x5 | ~x7) : (x5 | x7))) & (x3 | ~x4 | x5 | x7)));
  assign n3603 = x4 ? (x3 ? n3605 : n3604) : n3606;
  assign n3604 = (x0 | x1 | ~x5 | ~x6 | x7) & (~x0 | ~x1 | x5 | x6 | ~x7);
  assign n3605 = (x0 | ~x1 | x7 | (~x5 ^ x6)) & (x1 | (x0 ? (~x6 | (~x5 ^ x7)) : (x5 | x6)));
  assign n3606 = (~n978 | ~n727) & (~n1051 | n3607);
  assign n3607 = x0 ? (~x1 | ~x7) : (x1 ? (~x5 | x7) : (x5 | ~x7));
  assign n3608 = ~n640 & (n3610 | ~n3611 | (~x1 & ~n3609));
  assign n3609 = (x4 | ((x0 | ~x2 | ~x3 | x5) & (~x0 | (x2 ? (x3 | ~x5) : (~x3 | x5))))) & (x3 | ~x4 | ((x2 | x5) & (x0 | ~x2 | ~x5)));
  assign n3610 = ~x1 & ((x4 & x5 & ~x0 & ~x2) | (x0 & (x2 ? (x4 & ~x5) : (~x4 & x5))));
  assign n3611 = ~n3612 & (~n1392 | ~n632 | (~x0 & ~n1380));
  assign n3612 = ~x0 & x1 & ~x4 & (x2 | ~x5);
  assign n3613 = ~n3616 & (x1 | (~n3614 & ~n3615));
  assign n3614 = ~n1010 & ((n569 & n1966) | (~x2 & ~n1116));
  assign n3615 = n1769 & (x0 ? (~x4 & ~x5) : (x2 & x4));
  assign n3616 = x1 & (x0 ? (n942 & n1084) : ~n3617);
  assign n3617 = (~x4 | ((~x5 | x6 | ~x7) & (~x2 | x5 | ~x6 | x7))) & (x2 | ((x4 | ~x5 | ~x6 | x7) & (~x4 | x6 | ~x7)));
  assign z165 = ~n3630 | (x0 ? ~n3626 : ~n3619);
  assign n3619 = ~n3620 & (x6 | (n3624 & (~x1 | n3623)));
  assign n3620 = x6 & ((~x5 & ~n3621) | (n1301 & ~n3622));
  assign n3621 = (~x3 | (x1 ? (x2 ? (~x4 | ~x7) : x7) : (x2 ? x7 : (~x4 | ~x7)))) & (x4 | ((~x1 | x2 | x7) & (x1 | ~x2 | x3 | ~x7)));
  assign n3622 = x1 ? (x2 ? x7 : (~x4 | ~x7)) : (x2 ? (~x4 | ~x7) : x7);
  assign n3623 = (~x3 | x7 | (x2 ? (x4 | ~x5) : (~x4 | x5))) & (x3 | ~x4 | x5 | ~x7) & (x2 | ~x5 | ((x4 | ~x7) & (x3 | (x4 & ~x7))));
  assign n3624 = (n2017 | n3625) & (~n717 | ~n676);
  assign n3625 = x1 ? (~x2 | ~x5) : (x2 ^ ~x5);
  assign n3626 = (x2 | n3627) & (x1 | ~x2 | n3629);
  assign n3627 = x4 ? n3628 : (x1 | (n1647 & ~n2939));
  assign n3628 = (x3 | ((~x6 | ~x7 | x1 | ~x5) & (~x1 | ((~x6 | x7) & (x5 | x6 | ~x7))))) & (x1 | ~x3 | (~x5 ^ x7));
  assign n3629 = (~x4 | ((~x5 | x6 | ~x7) & (~x3 | x5 | x7))) & (x3 | x4 | x5 | x6 | ~x7) & (~x3 | ~x6 | (~x5 ^ ~x7));
  assign n3630 = ~n3631 & (n3315 | n3634);
  assign n3631 = ~n640 & ((~n1548 & ~n3632) | (~x3 & ~n3633));
  assign n3632 = (x0 | x2 | (~x1 ^ x5)) & (x1 | ~x2 | x5);
  assign n3633 = (~x0 | x1 | x5 | (x2 & x4)) & (~x5 | (x0 ? (~x1 | x2) : (x1 ? ~x2 : (x2 | x4))));
  assign n3634 = (x4 | ((x1 | ~x2 | ~x5) & (~x0 | ~x1 | x2 | x5))) & (x0 | (x1 ? (x2 ? x5 : (~x4 | ~x5)) : (~x2 ^ ~x5)));
  assign z166 = ~n3647 | n3644 | n3636 | n3641;
  assign n3636 = ~x2 & ((~x7 & ~n3638) | (n3637 & ~n3640));
  assign n3637 = x0 & x7;
  assign n3638 = (x5 | n3639) & (~x4 | ~x5 | ~n841 | n1026);
  assign n3639 = (~x0 | x1 | ~x3 | ~x4 | ~x6) & (x0 | ((x4 | ~x6 | x1 | x3) & (~x1 | (x3 ? (~x4 | ~x6) : (x4 | x6)))));
  assign n3640 = (~x1 | x3 | x4 | ~x5 | x6) & (x1 | ((x3 | ~x4 | ~x5 | x6) & (~x3 | ~x6 | (~x4 & ~x5))));
  assign n3641 = x2 & (n3642 | (~n1555 & (n529 | n841)));
  assign n3642 = ~x1 & (x0 ? ~n3643 : (n1029 & n978));
  assign n3643 = (~x6 | ((x3 | x4 | x5 | ~x7) & (~x3 | (x4 ? x5 : (~x5 | x7))))) & (x3 | x6 | ((~x5 | x7) & (~x4 | x5 | ~x7)));
  assign n3644 = x4 & (~n3646 | (~x0 & ~n3645));
  assign n3645 = (x2 | x5 | (x3 ? (~x6 | ~x7) : (x6 | x7))) & (~x2 | ~x3 | ~x5 | ~x6 | ~x7);
  assign n3646 = (~x0 | x2 | x3 | x5 | x6) & (x0 | ((~x5 | ((x3 | x6) & (x2 | ~x3 | ~x6))) & (~x2 | (x3 ? (x5 | ~x6) : x6))));
  assign n3647 = ~n3650 & (n643 | (~n3648 & (~x3 | n3649)));
  assign n3648 = ~n1954 & (n2857 | (x0 & ~n647));
  assign n3649 = (x1 | x2 | x4) & (x0 | (x1 ? (~x2 | x4) : (x2 | x5)));
  assign n3650 = ~x4 & ((n1693 & n813) | (~x3 & ~n3651));
  assign n3651 = (x0 | ((~x6 | ~x7) & (~x5 | x6 | x7))) & (x2 | ((x5 | ~x6 | ~x7) & (~x0 | x6 | x7)));
  assign z167 = ~n3662 | (~x0 & ~n3653) | (x2 & ~n3659);
  assign n3653 = (~x3 & n3657) | (~n3655 & n3656 & x3 & ~n3654);
  assign n3654 = ~n2022 & n3051;
  assign n3655 = ~n671 & ((n904 & n804) | (n1364 & n1133));
  assign n3656 = (~x2 | ~x4 | ~x5 | x6 | ~x7) & (x2 | x4 | x5 | ~x6 | x7);
  assign n3657 = (x5 | n3658) & (~n1769 | ~n859 | ~x1 | ~x5);
  assign n3658 = (x1 | ((x6 | ~x7 | x2 | x4) & (~x2 | x7 | (~x4 ^ x6)))) & (x2 | ~x4 | ((~x6 | ~x7) & (~x1 | x6 | x7)));
  assign n3659 = ~n3661 & (x0 ? (~n1188 | ~n867) : n3660);
  assign n3660 = (x1 | x3 | ~x4 | x5 | ~x7) & (x4 | ~x5 | x7 | (~x1 & ~x3));
  assign n3661 = ~n1218 & (n1600 | (~x5 & (n727 | ~n823)));
  assign n3662 = (~n872 | n3669) & (x2 | (n3663 & n3666));
  assign n3663 = ~n3664 & ~n3665 & (~n727 | ~n809);
  assign n3664 = x0 & ~x1 & (x3 ? (~x4 & ~x7) : (x4 & x7));
  assign n3665 = ~x0 & x1 & (x3 ? (x4 & x7) : (~x4 & ~x7));
  assign n3666 = (n791 | n3667) & (x3 | n3668);
  assign n3667 = x1 ? (x3 ? (x4 | x7) : (~x4 | ~x7)) : (x3 ? (~x4 | ~x7) : (x4 | x7));
  assign n3668 = (~x0 | ~x1 | ~x4 | ~x5 | x7) & ((x0 ? (~x1 | x4) : (x1 | ~x4)) | (~x5 ^ ~x7));
  assign n3669 = x7 ? ((x2 | ((x4 | ~x6) & (~x3 | ~x4 | x6))) & (x3 | ((x4 | ~x6) & (~x2 | ~x4 | x6)))) : ((~x2 | (~x4 ^ ~x6)) & (x3 | x4 | x6));
  assign z168 = ~n3671 | n3678 | (x1 & ~n3681);
  assign n3671 = n3674 & (x0 | (n3673 & (~x1 | n3672)));
  assign n3672 = (x2 | x3 | x4 | x5 | x6) & (~x4 | ((~x2 | (x3 ? (~x5 | ~x6) : (x5 | x6))) & (x2 | x3 | x5 | ~x6)));
  assign n3673 = (x1 | ((~x2 | x3 | x5 | ~x6) & (x2 | ~x5 | x6))) & (~x3 | x5 | ((~x1 | ~x2 | x6) & (x2 | ~x6)));
  assign n3674 = n3677 & (~n841 | n3675) & (~n681 | n3676);
  assign n3675 = (x3 & (x2 ? (x4 & ~x6) : ~x4)) | (~x5 & x6) | (x5 & ~x6) | (~x2 & x4 & (~x3 | x6));
  assign n3676 = (x0 | ~x1 | ~x2 | x3) & (x2 | ~x3 | ~x0 | x1);
  assign n3677 = (x0 | x1 | ~x2 | ~x3 | x5) & (~x0 | ~x1 | x2 | x3 | ~x5);
  assign n3678 = ~x1 & (~n3680 | (~n815 & ~n3679));
  assign n3679 = x0 ? (~x3 | ((~x5 | ~x7) & (~x4 | x5 | x7))) : (x3 | (~x5 ^ x7));
  assign n3680 = (~n662 | ~n2435) & (~n622 | ~n1429 | n1171);
  assign n3681 = x0 ? (~n1044 | ~n588) : (~n3682 & ~n3683);
  assign n3682 = ~n1548 & ((n1857 & n691) | (x2 & n702));
  assign n3683 = n934 & (n684 | n3684);
  assign n3684 = ~x7 & x6 & ~x3 & ~x4;
  assign z169 = n3686 | n3690 | ~n3697 | (~n640 & ~n3693);
  assign n3686 = ~x0 & (n3688 | (n558 & n3687));
  assign n3687 = x7 & x6 & ~x4 & ~x5;
  assign n3688 = x4 & ((n978 & n669) | (x2 & ~n3689));
  assign n3689 = (x1 | x3 | ~x5 | x6 | ~x7) & (~x1 | x5 | (x3 ? (x6 | x7) : (~x6 | ~x7)));
  assign n3690 = ~n643 & (x5 ? ~n3692 : ~n3691);
  assign n3691 = x0 ? ((~x1 | x2 | x3 | x4) & (x1 | ~x4 | (~x2 ^ ~x3))) : (x1 ? (x2 | ~x3) : (~x2 | x3));
  assign n3692 = (~x2 | ~x3 | ~x0 | x1) & (x0 | ((x1 | ~x2 | x3 | x4) & (~x1 | x2 | (~x3 ^ x4))));
  assign n3693 = ~n3694 & ~n3695 & ~n3696 & (~n1287 | ~n1209);
  assign n3694 = x4 & x3 & ~x2 & x0 & ~x1;
  assign n3695 = n1380 & ((n1392 & n1133) | (~x1 & ~n2075));
  assign n3696 = ~x0 & ((x1 & ~x4 & (x2 ^ ~x3)) | (~x3 & x4 & ~x1 & ~x2));
  assign n3697 = ~n3700 & n3702 & (x0 ? n3698 : n3699);
  assign n3698 = (x1 | x2 | ~x3 | x4 | x6) & (x3 | ((~x1 | x2 | ~x4 | x6) & (x1 | ~x6 | (~x2 ^ ~x4))));
  assign n3699 = (x1 | x2 | ~x3 | x4 | ~x6) & (~x2 | ((~x1 | (x3 ? (~x4 | ~x6) : (x4 | x6))) & (x4 | x6 | x1 | ~x3)));
  assign n3700 = n872 & ~n3701;
  assign n3701 = (~x2 | x3 | x4 | x6 | x7) & (x2 | ~x7 | (x3 ? (x4 | ~x6) : (~x4 | x6)));
  assign n3702 = (n1566 | n3703 | ~x0 | x4) & (x0 | ~x4 | n3704);
  assign n3703 = x1 ? (x2 | x6) : (~x2 | ~x6);
  assign n3704 = (~x1 | x2 | ~x3 | ~x5 | x6) & (x5 | (x2 ^ ~x6) | (x1 ^ ~x3));
  assign z170 = n3706 | ~n3712 | n3718 | (~x1 & ~n3717);
  assign n3706 = ~x0 & (n3707 | n3710);
  assign n3707 = x1 & ((n859 & n3709) | (~x6 & ~n3708));
  assign n3708 = (~x4 | x5 | x7 | ~x2 | x3) & (x2 | ~x7 | (x3 ? (~x4 | x5) : (x4 | ~x5)));
  assign n3709 = ~x5 & x6 & (~x3 ^ ~x7);
  assign n3710 = n3711 & ((x2 & ~x3 & (x6 ^ x7)) | (x3 & (x2 ? (~x6 & ~x7) : (x6 & x7))));
  assign n3711 = x5 & ~x1 & x4;
  assign n3712 = ~n3714 & n3716 & (~n872 | n3713);
  assign n3713 = (~x6 | ((x4 | x7 | ~x2 | x3) & (x2 | (x3 ? (x4 | ~x7) : (~x4 | x7))))) & (~x2 | x4 | x6 | (x3 ^ ~x7));
  assign n3714 = x0 & (x4 ? (n757 & n558) : ~n3715);
  assign n3715 = x5 ? ((x1 | ~x2 | ~x3 | ~x7) & (x3 | x7 | ~x1 | x2)) : ((~x1 ^ x2) | (~x3 ^ x7));
  assign n3716 = (n1580 | n1581) & (~n837 | ~n2648);
  assign n3717 = (x4 | x7 | ~x0 | x2) & (x0 | (x2 & x4) | (~x3 ^ x7));
  assign n3718 = ~x0 & ((n2296 & n576) | (x4 & ~n3719));
  assign n3719 = x1 ? (x3 ? (~x5 | x7) : ((~x5 | ~x7) & (x2 | x5 | x7))) : (~x2 | (x3 ? (~x5 ^ ~x7) : (x5 | ~x7)));
  assign z171 = ~n3726 | (~x0 & (n3721 | n3723 | ~n3724));
  assign n3721 = ~x4 & ((n558 & n951) | (~x7 & ~n3722));
  assign n3722 = (~x1 | ~x2 | x3 | x5 | ~x6) & (x1 | ~x3 | ~x5 | (x2 ^ ~x6));
  assign n3723 = ~n2290 & ~n815 & x7 & n1029;
  assign n3724 = (x1 | n3725) & (x5 | n1353 | ~x1 | ~x2);
  assign n3725 = (x2 | x3 | x4 | x5 | ~x6) & (~x5 | ((x2 | ~x3 | x4 | x6) & (~x2 | ((~x4 | ~x6) & (x3 | x4 | x6)))));
  assign n3726 = n3729 & (x2 | n3727) & (~n841 | n3728);
  assign n3727 = (x1 | ((~x4 | ~x5 | ~x0 | x3) & (x0 | x4 | (~x3 ^ x5)))) & (~x0 | ~x1 | x3 | (~x4 ^ x5));
  assign n3728 = (~n813 | ~n1556) & (~n1301 | n671 | n815);
  assign n3729 = n3731 & (~n872 | n3730);
  assign n3730 = (x2 | ~x3 | ~x4 | x6) & (~x2 | ((x4 | ~x6) & (x3 | ~x4 | x6)));
  assign n3731 = (~x0 | x1 | ~x4 | x5) & (x0 | ((x1 | ~x2 | x4 | x5) & (~x1 | ((~x4 | ~x5) & (x2 | x4 | x5)))));
  assign z172 = ~n3738 | (~x0 & ~n3733) | (~x1 & ~n3736);
  assign n3733 = ~n3735 & (~x1 | (~n3734 & (~n1070 | ~n1780)));
  assign n3734 = x3 & ~n815 & ((x5 & ~x7) | (x4 & ~x5 & x7));
  assign n3735 = n669 & n830;
  assign n3736 = (x4 | n3737) & (n765 | n815 | ~x3 | ~x4);
  assign n3737 = x2 ? ((x3 | x5 | ~x6 | x7) & (x6 | ~x7 | ~x3 | ~x5)) : (~x7 | (x3 ? (~x5 | ~x6) : (x5 | x6)));
  assign n3738 = ~n3739 & n3742 & (~n543 | n3741);
  assign n3739 = ~x5 & ((n527 & ~n920) | (x6 & ~n3740));
  assign n3740 = (x0 | ~x1 | ~x2 | x3 | ~x4) & (~x0 | x1 | x2 | ~x3 | x4);
  assign n3741 = (~x2 | (x3 ? (x5 | ~x6) : (~x5 | x6))) & (x2 | ~x3 | ~x5 | x6);
  assign n3742 = ~n3743 & (~n576 | ~n588) & (~n1188 | n1447);
  assign n3743 = ~x3 & (x1 ? (~x2 & x5) : (x2 ? (x5 ^ ~x6) : (~x5 & x6)));
  assign z173 = n3746 | ~n3749 | (~n643 & ~n3745);
  assign n3745 = (x1 & (~x0 ^ x2)) | (~x2 & ~n1287) | (x2 & ~n843);
  assign n3746 = ~x4 & ((n1209 & n3747) | (n1310 & ~n3748));
  assign n3747 = ~x7 & ~x6 & ~x3 & x5;
  assign n3748 = (~x2 | ~x3 | ~x6 | x7) & (x2 | ~x7 | (x1 ? (x3 | x6) : (~x3 | ~x6)));
  assign n3749 = ~n3750 & n3753 & (~n841 | ~n865 | n3752);
  assign n3750 = ~n3751 & ~n640 & ~n710;
  assign n3751 = (x4 | x5 | ~x2 | x3) & (x2 | ~x3 | (~x4 & ~x5));
  assign n3752 = x3 ^ (~x4 & ~x5);
  assign n3753 = (~n878 | n3752) & (~n742 | ~n971 | n3754);
  assign n3754 = ~x4 & ~x5;
  assign z174 = (~x4 | ~n3760) & (x4 | n3756 | n3759 | ~n3761);
  assign n3756 = ~x1 & ((x0 & ~n3757) | (n1310 & ~n3758));
  assign n3757 = (~x2 | x3 | ~x5 | ~x6 | x7) & (x2 | x6 | (x3 ? (~x5 | x7) : (x5 | ~x7)));
  assign n3758 = (~x3 | ~x6 | ~x7) & (~x2 | x6 | (~x3 ^ x7));
  assign n3759 = n1291 & (x2 ? (x3 & n1300) : (~x3 & ~n643));
  assign n3760 = (~x3 & x7) | (x3 & ~x7) | (x0 & x1 & (x2 | x7));
  assign n3761 = (~x3 | n3765) & (x3 | n3763) & (n3762 | n3764);
  assign n3762 = x0 ? (~x1 | x2) : (~x1 ^ ~x2);
  assign n3763 = (x0 | ~x1 | x2 | ~x5 | x7) & (x1 | ((~x5 | x7 | x0 | ~x2) & (~x0 | (x2 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n3764 = x3 ? (x5 | x7) : (x5 ^ ~x7);
  assign n3765 = (x0 | ((~x5 | ~x7) & (~x1 | x2 | x5 | x7))) & (x1 | ((~x5 | ~x7) & (~x0 | x5 | x7)));
  assign z175 = ~n3768 | n3774 | n3776 | (~x1 & ~n3767);
  assign n3767 = (~x0 | ~x4 | x5 | (x2 ^ ~x3)) & (x4 | ~x5 | (x0 & (x2 | x3)));
  assign n3768 = n3772 & (~n689 | n3769) & (n714 | n3771);
  assign n3769 = (~n943 | ~n2057) & (~x6 | ~n1310 | n3770);
  assign n3770 = x2 ? (x4 | ~x7) : (~x4 | x7);
  assign n3771 = (~x2 | ~x3 | ~x0 | x1) & (~x1 | ((x2 | x3) & (x0 | (x2 & x3))));
  assign n3772 = (~n639 | ~n746) & (~x6 | n2227 | ~n3773);
  assign n3773 = x5 & ~x4 & x0 & ~x1;
  assign n3774 = ~x5 & ((n560 & n1331) | (~x0 & ~n3775));
  assign n3775 = (~x2 | ~x3 | ~x4 | x6) & (~x1 | x2 | x3 | x4 | ~x6) & (x1 | ((~x4 | x6) & (x4 | ~x6 | ~x2 | ~x3)));
  assign n3776 = ~n671 & ((~n1446 & n1511) | (x3 & ~n3777));
  assign n3777 = (~x0 | x1 | x2 | ~x5 | x6) & (x0 | x5 | ~x6 | (~x1 ^ ~x2));
  assign z176 = n3779 | ~n3782 | ~n3784 | (~n2227 & ~n3781);
  assign n3779 = n3151 & ((n746 & n2834) | (~x2 & ~n3780));
  assign n3780 = (x0 | ~x1 | ~x4 | ~x6 | x7) & (~x0 | x1 | ~x7 | (~x4 ^ ~x6));
  assign n3781 = (x1 | ((~x7 | ((~x5 | x6) & (x0 | x5 | ~x6))) & (~x0 | (x5 ? ~x6 : (x6 | x7))))) & (x0 | ~x5 | (x6 & (~x1 | x7)));
  assign n3782 = ~n3783 & (~n1322 | ~n1269) & (~n560 | ~n3747);
  assign n3783 = x5 & ((x0 & ~n3275) | (n3074 & (~n3275 | ~n3482)));
  assign n3784 = ~n3785 & (x5 | (~n3787 & ~n3789));
  assign n3785 = x6 & (n3786 | (~n1008 & (n664 | n2144)));
  assign n3786 = ~x0 & ~x2 & x5 & (x1 ^ ~x7);
  assign n3787 = ~n3788 & ~x1 & ~n697;
  assign n3788 = (x0 | x3 | ~x4 | ~x6) & (x4 | x6 | ~x0 | ~x3);
  assign n3789 = n3791 & (n2359 | n3790);
  assign n3790 = ~x7 & x4 & ~x6;
  assign n3791 = ~x3 & ~x2 & ~x0 & x1;
  assign z177 = ~n3793 | (~x7 & ~n3805) | (x2 & ~n3804);
  assign n3793 = n3803 & ~n3801 & ~n3800 & ~n3794 & ~n3798;
  assign n3794 = x7 & ((n3795 & n3796) | (n1084 & ~n3797));
  assign n3795 = x4 & (x5 ^ ~x6);
  assign n3796 = ~x3 & x2 & ~x0 & x1;
  assign n3797 = (x0 | x1 | x3 | x5 | x6) & ((~x1 ^ x5) | (x0 ? (~x3 | x6) : (x3 | ~x6)));
  assign n3798 = ~x1 & ((n1786 & n1783) | (x4 & ~n3799));
  assign n3799 = (x0 | x2 | x3 | x6 | x7) & ((x2 ^ ~x7) | (x0 ? (~x3 | x6) : (x3 | ~x6)));
  assign n3800 = n873 & ((n1156 & n1769) | (~x2 & ~n1850));
  assign n3801 = ~n640 & (n2144 | (~x0 & x3 & ~n3802));
  assign n3802 = x1 ^ x2;
  assign n3803 = ~n1923 & (~n560 | ~n3057) & (~n825 | n3703);
  assign n3804 = (x0 | ~x1 | x3 | x6 | x7) & (x1 | ((~x6 | ~x7 | x0 | x3) & (~x0 | ((x6 | ~x7) & (x3 | ~x6 | x7)))));
  assign n3805 = ~n3806 & (~n1269 | ~n1643) & (n1198 | n3807);
  assign n3806 = ~x2 & (x0 ? ~n897 : (n689 & n728));
  assign n3807 = (x0 | ~x1 | x2 | x3 | ~x4) & (~x0 | x1 | ~x2 | ~x3 | x4);
  assign z178 = n3809 | n3813 | ~n3816 | (~x3 & ~n3815);
  assign n3809 = ~x2 & (n3810 | (n841 & n3812));
  assign n3810 = ~x3 & (x0 ? (n772 & n978) : ~n3811);
  assign n3811 = x1 ? (~x7 | (x4 ? (x5 | x6) : (~x5 | ~x6))) : (x4 | x7 | (~x5 ^ x6));
  assign n3812 = x3 & ~x4 & ~x5 & (x6 ^ ~x7);
  assign n3813 = ~x1 & (x4 ? (n757 & n600) : ~n3814);
  assign n3814 = (x0 | ~x2 | x3 | x5 | ~x7) & (~x5 | ((x0 | x2 | x3 | ~x7) & (~x0 | ~x3 | (x2 ^ ~x7))));
  assign n3815 = (x0 | ~x1 | x4 | x7) & (x1 | ((x4 | ~x7 | ~x0 | x2) & (x0 | ~x4 | (~x2 ^ x7))));
  assign n3816 = n3822 & ~n3821 & ~n3817 & ~n3819;
  assign n3817 = n3818 & (x0 ? (x3 & n951) : (~x3 & n2153));
  assign n3818 = ~x4 & ~x1 & x2;
  assign n3819 = x1 & ((n594 & n2209) | (n539 & ~n3820));
  assign n3820 = x2 ? (~x5 ^ ~x7) : (~x5 | x7);
  assign n3821 = ~x0 & x3 & (x1 ? (x2 ^ ~x7) : (x2 ^ x7));
  assign n3822 = (n697 | ~n936) & (~n622 | n3823);
  assign n3823 = x1 ? (x2 | x7) : (~x2 | ~x7);
  assign z179 = ~n3825 | (n2359 & ~n3834) | (x4 & ~n3833);
  assign n3825 = ~n3829 & ~n3831 & ~n3832 & (x4 | n3826);
  assign n3826 = (~n719 | ~n3828) & (~x6 | ~n2061 | n3827);
  assign n3827 = (x3 | x7 | ~x1 | x2) & (~x3 | ~x7 | x1 | ~x2);
  assign n3828 = ~x2 & ~x0 & ~x1;
  assign n3829 = ~n1954 & ~n3830;
  assign n3830 = (~x0 | x3 | x4 | x5 | x6) & (x0 | (x3 ? (x4 | (x5 & x6)) : (~x4 | ~x5)));
  assign n3831 = n774 & (x0 ? (~x1 & x5) : (x1 ? x2 : (~x2 & ~x5)));
  assign n3832 = n1012 & ((n1044 & n1070) | (n885 & n658));
  assign n3833 = x0 ? (x1 | ~x3) : (x1 ? ((~x2 | x3 | ~x5) & (~x3 | x5)) : (x3 | (x2 & x5)));
  assign n3834 = (~x0 | x1 | x2 | ~x3 | x5) & (x0 | ~x5 | (x1 ? (x2 | ~x3) : x3));
  assign z180 = n3845 | ~n3844 | ~n3841 | n3836 | ~n3839;
  assign n3836 = ~x0 & (n3837 | (n669 & n1725));
  assign n3837 = x4 & ((n978 & n1439) | (n918 & ~n3838));
  assign n3838 = (x2 | x3 | x5 | ~x6) & (~x2 | ~x3 | ~x5 | x6);
  assign n3839 = ~n3840 & (~n993 | ~n2144) & (~n841 | ~n1622);
  assign n3840 = x1 & ((n743 & n1311) | (~x0 & ~n3538));
  assign n3841 = (n671 | n3843) & (~x6 | ~n1145 | n3842);
  assign n3842 = x0 ? (x5 | (x2 ^ ~x3)) : ~x5;
  assign n3843 = (~n1519 | ~n816) & (~x6 | ~n2061 | n3275);
  assign n3844 = (~x0 | x1 | ~x2 | x4 | ~x5) & (x0 | (x1 ? (x2 ? (x4 | x5) : (~x4 | ~x5)) : (~x4 | x5)));
  assign n3845 = x4 & (n3846 | (n527 & ~n791 & ~n2737));
  assign n3846 = x1 & ((n743 & n3848) | (n742 & n3847));
  assign n3847 = x6 & x3 & x5;
  assign n3848 = ~x6 & ~x3 & ~x5;
  assign z181 = n3850 | ~n3856 | (~x0 & ~n3854);
  assign n3850 = ~x2 & (n3851 | (n1511 & n3853));
  assign n3851 = ~x0 & (x6 ? (n1317 & ~n2216) : ~n3852);
  assign n3852 = (x3 | ((~x1 | (~x4 ^ ~x5)) & (x5 | x7 | x1 | ~x4))) & (x1 | ~x3 | ~x7 | (~x4 ^ x5));
  assign n3853 = ~x4 & x5 & (x6 | x7);
  assign n3854 = (~x3 | ~n943 | ~x1 | ~x2) & (x1 | ((x2 | x3 | ~n943) & (~x3 | n3855)));
  assign n3855 = (x6 | x7 | x2 | x5) & (~x6 | ~x7 | ~x2 | ~x5);
  assign n3856 = ~n3861 & ~n3860 & ~n3859 & ~n3857 & ~n3858;
  assign n3857 = ~n2227 & (x0 ? (~x1 & (x5 ^ x6)) : (x5 & (x1 | x6)));
  assign n3858 = x5 & ((n2337 & ~n3275) | (n1686 & ~n3482));
  assign n3859 = ~x6 & ~x5 & x2 & ~x0 & ~x1;
  assign n3860 = x0 & ((n558 & n813) | (n881 & ~n3275));
  assign n3861 = ~n3862 & n742 & n1903;
  assign n3862 = (x1 | x4 | ~x5 | ~x6) & (~x1 | x6 | (x4 ^ ~x5));
  assign z182 = ~n3871 | ~n3868 | n3864 | n3867;
  assign n3864 = x3 & (n3865 | (x2 & n592 & n626));
  assign n3865 = ~x4 & ((~n790 & n1411) | (n2061 & ~n3866));
  assign n3866 = (x6 | x7 | ~x1 | x2) & (~x6 | ~x7 | x1 | ~x2);
  assign n3867 = ~x1 & x6 & ((x2 & ~x3) | (x0 & ~x2 & x3));
  assign n3868 = ~n3869 & n3870 & (n1532 | ~n825 | n682);
  assign n3869 = n662 & n2144;
  assign n3870 = x0 | ~x1 | (x2 ? ~n1051 : ~n3497);
  assign n3871 = x6 ? (x7 ? n3872 : n3873) : (x7 ? n3873 : n3872);
  assign n3872 = ~n576 & ~n2282 & (~x5 | n807 | ~n2343);
  assign n3873 = (x1 | x2 | x3) & (x0 | ((~x3 | ~x4 | ~x1 | ~x2) & (x1 | x2 | x4)));
  assign z183 = ~n3877 | (x0 & (n3875 | (n558 & n1241)));
  assign n3875 = ~x6 & (x1 ? (n2296 & n902) : ~n3876);
  assign n3876 = (~x2 | ~x3 | x4 | x5 | x7) & (x2 | x3 | ~x4 | ~x5 | ~x7);
  assign n3877 = n3879 & (~n825 | (n3878 & n3882 & n3883));
  assign n3878 = (x1 | x4 | (~x2 ^ x7)) & (~x4 | ((x2 | x7) & (~x1 | ~x2 | ~x7)));
  assign n3879 = ~n3880 & ~n3881 & (~n560 | (~n2647 & ~n2992));
  assign n3880 = ~x1 & ((x0 & x3 & (x2 ^ ~x7)) | (~x3 & ((x2 & ~x7) | (~x0 & ~x2 & x7))));
  assign n3881 = x1 & ~x3 & ((~x2 & x7) | (~x0 & x2 & ~x7));
  assign n3882 = (x1 | ~x2 | ~x4 | ~x5 | ~x7) & (x7 | ((x1 | ~x2 | ~x4 | x5) & (~x1 | x4 | (~x2 ^ x5))));
  assign n3883 = (~x4 | ~n1070 | x1 | ~x2) & (~x1 | x4 | n3884);
  assign n3884 = (x2 | x5 | x6 | ~x7) & (~x2 | ~x5 | (~x6 ^ ~x7));
  assign z184 = ~n3897 | ~n3893 | n3891 | n3886 | n3889;
  assign n3886 = ~x7 & (n3887 | (~x2 & n922 & n959));
  assign n3887 = ~x4 & ((n1746 & n746) | (x3 & ~n3888));
  assign n3888 = (~x1 | x2 | x5 | ~x6) & (x1 | ~x2 | (x0 ? (x5 | x6) : (~x5 | ~x6)));
  assign n3889 = n1465 & ((n926 & n746) | (x6 & ~n3890));
  assign n3890 = (x4 | ~x5 | x1 | x2) & (x0 | ((x2 | x4 | ~x5) & (~x1 | ~x2 | ~x4 | x5)));
  assign n3891 = ~n3892 & (x1 ? ~x3 : (x3 & x6));
  assign n3892 = (x0 | ~x2 | (x4 ? (x5 | x7) : (~x5 | ~x7))) & (~x0 | x2 | ~x4 | ~x5 | ~x7);
  assign n3893 = ~n3894 & n3896 & (x4 | ~n825 | ~n3895);
  assign n3894 = ~x0 & ((~x4 & ~x5 & x2 & x3) | (~x3 & x4 & (~x2 | x5)));
  assign n3895 = ~x6 & (x2 ^ ~x5);
  assign n3896 = ~n2030 & (~n743 | ~n1268) & (~n560 | ~n1759);
  assign n3897 = ~n3899 & (x4 | n3898);
  assign n3898 = (x0 | x1 | x2 | ~x3 | ~x5) & (~x0 | x3 | (x1 ? (x2 | ~x5) : ~x2));
  assign n3899 = ~x5 & ((~n627 & ~n3900) | (n1141 & n816));
  assign n3900 = (x0 | x1 | ~x2 | ~x4) & (x2 | x4 | ~x0 | ~x1);
  assign z185 = n3919 | n3917 | ~n3910 | n3902 | n3908;
  assign n3902 = ~x2 & (n3904 | (n3903 & ~n3907));
  assign n3903 = x3 & x6;
  assign n3904 = ~x3 & ((~x1 & ~n3905) | (n3236 & ~n3906));
  assign n3905 = (~x0 | ~x4 | ~x5 | x6 | ~x7) & (x4 | ((~x5 | ~x6 | x7) & (x6 | ~x7 | x0 | x5)));
  assign n3906 = (~x4 | x5 | ~x7) & (x0 | x4 | ~x5 | x7);
  assign n3907 = (~x1 | x4 | x5 | x7) & (~x0 | x1 | ~x5 | (~x4 ^ x7));
  assign n3908 = ~x1 & ~n3909;
  assign n3909 = (~x0 | ~x2 | x3 | ~x4 | x5) & (x2 | (x0 ? (x5 | (~x3 ^ ~x4)) : (~x3 | x4)));
  assign n3910 = n3914 & (~x2 | (~n3911 & ~n3913));
  assign n3911 = ~x6 & ((~n1218 & ~n3912) | (n2296 & n1244));
  assign n3912 = (~x0 | x1 | ~x3 | x5) & (x0 | ~x1 | x3 | ~x5);
  assign n3913 = n852 & ((~x1 & ~x5 & (x4 ^ x7)) | (x5 & x7 & x1 & x4));
  assign n3914 = ~n3915 & ~n3916 & (~n959 | ~n837);
  assign n3915 = x5 & x4 & x2 & x0 & ~x1;
  assign n3916 = ~x0 & ((x1 & (x2 ? (~x4 & ~x5) : (x4 & x5))) | (~x1 & x2 & ~x4 & x5));
  assign n3917 = x2 & (x0 ? (n592 & n1188) : ~n3918);
  assign n3918 = x1 ? (~x5 | (x3 ? (x4 | x6) : (~x4 | ~x6))) : (x5 | ((~x4 | x6) & (x3 | x4 | ~x6)));
  assign n3919 = ~x2 & ((n704 & n1244) | (~x6 & ~n3920));
  assign n3920 = (~x0 | ((x1 | ~x3 | ~x4 | ~x5) & (~x1 | x4 | x5))) & (x4 | ((~x1 | ~x3 | x5) & (x3 | ~x5 | (x0 & x1))));
  assign z186 = n3932 | ~n3935 | (x1 ? ~n3922 : ~n3927);
  assign n3922 = ~n3926 & (x0 | (~n3923 & (~n859 | n3925)));
  assign n3923 = ~x4 & ((n596 & n658) | (n778 & ~n3924));
  assign n3924 = x3 ? (x5 | x7) : (~x5 | ~x7);
  assign n3925 = (x3 | x6 | (~x5 ^ x7)) & (~x3 | ~x5 | ~x6 | x7);
  assign n3926 = n594 & n830;
  assign n3927 = x5 ? (x2 | n3931) : (~n3928 & ~n3930);
  assign n3928 = ~n3929 & (x0 ? n1029 : n828);
  assign n3929 = x2 ? (x6 | x7) : (~x6 | ~x7);
  assign n3930 = x6 & ((n566 & ~n1410) | (n743 & n2647));
  assign n3931 = (x3 | x4 | ~x6 | x7) & (~x3 | ((~x0 | ~x6 | x7) & (x6 | ~x7 | x0 | ~x4)));
  assign n3932 = ~x2 & ((~x5 & ~n3933) | (n551 & ~n3934));
  assign n3933 = (~x3 | ((x0 | ~x1 | ~x4) & (x4 | ~x6 | ~x0 | x1))) & (~x1 | ((x3 | ~x4 | x6) & (x0 | (x6 & (x3 | x4)))));
  assign n3934 = (~x0 & x3 & x4 & ~x6) | (x6 & (x0 | (~x3 & ~x4)));
  assign n3935 = ~n3938 & ~n3939 & (~x2 | (~n3936 & n3937));
  assign n3936 = n1167 & ((~x1 & ~n981) | (n904 & n1317));
  assign n3937 = (x0 | ~x1 | x5 | ~x6) & (~x5 | ((x0 | ~x1 | ~x3 | x6) & (~x0 | x1 | (x3 & ~x6))));
  assign n3938 = ~n3900 & ((~x5 & ~x6) | (~x3 & x5 & x6));
  assign n3939 = ~n765 & ((~n1062 & n1686) | (x0 & ~n3940));
  assign n3940 = (x1 | ~x2 | ~x3 | x4 | x6) & (~x1 | x2 | x3 | ~x4 | ~x6);
  assign z187 = n3947 | n3949 | ~n3953 | (~x1 & ~n3942);
  assign n3942 = x0 ? n3943 : (~n3946 & (n640 | n646));
  assign n3943 = x5 ? n3944 : (~n885 | n3945);
  assign n3944 = (~x3 | x4 | x6 | x7) & (~x7 | ((x2 | x3 | ~x4 | x6) & (~x2 | ~x6 | (x3 ^ ~x4))));
  assign n3945 = (x6 | x7) & (x4 | ~x6 | ~x7);
  assign n3946 = x3 & ((n1518 & n1070) | (x2 & ~n3409));
  assign n3947 = n543 & ((n530 & n949) | (~x3 & ~n3948));
  assign n3948 = (~x4 | ((~x2 | ~x6 | ~x7) & (x5 | x6 | x7))) & (~x5 | ((~x2 | (~x6 ^ ~x7)) & (x2 | x4 | ~x6 | x7)));
  assign n3949 = ~n643 & (n3950 | ~n3952 | (~x2 & ~n3951));
  assign n3950 = ~x0 & ((~x1 & x2 & x3) | (~x2 & (x1 ? (x3 ^ x4) : (~x3 & ~x4))));
  assign n3951 = (x0 | x1 | x3 | ~x4 | x5) & (~x0 | ~x3 | x4 | (x1 ^ ~x5));
  assign n3952 = (~n731 | ~n746) & (~n743 | n3042);
  assign n3953 = ~n3955 & n3957 & (~n551 | n3954);
  assign n3954 = (~x0 | ~x2 | ~x3 | ~x4 | x6) & (x0 | x3 | (x2 ? (x4 | x6) : (~x4 | ~x6)));
  assign n3955 = ~x5 & ((n971 & ~n1580) | (n1005 & ~n3956));
  assign n3956 = (x2 | x4 | ~x0 | x1) & (~x2 | ~x4 | x0 | ~x1);
  assign n3957 = (x4 | n3958) & (x0 | ~x4 | n1332);
  assign n3958 = x0 ? (x3 | (x1 ? (x2 | x6) : (~x2 | ~x6))) : (~x3 | (x1 ? (~x2 | x6) : (x2 | ~x6)));
  assign z188 = n3960 | ~n3965 | ~n3974 | (n543 & ~n3964);
  assign n3960 = ~x4 & ((~n3961 & ~n3962) | (~x3 & ~n3963));
  assign n3961 = x0 ? (x1 | x7) : (~x1 | ~x7);
  assign n3962 = (x5 | x6 | ~x2 | x3) & (~x5 | ~x6 | x2 | ~x3);
  assign n3963 = (~n943 | ~n837) & (x7 | ~n626 | n1446);
  assign n3964 = (x2 | x3 | ~x4 | ~x5 | x7) & (~x2 | ((x3 | x4 | ~x5 | x7) & (~x3 | ~x4 | (~x5 ^ x7))));
  assign n3965 = ~n3973 & ~n3970 & ~n3969 & ~n3966 & ~n3968;
  assign n3966 = ~n1205 & ~n3967;
  assign n3967 = (~x0 | ~x1 | x2 | x4 | x5) & (x0 | x1 | ~x5 | (~x2 ^ x4));
  assign n3968 = ~n1205 & (x0 ? (~x1 & ~n1532) : (x1 & n1084));
  assign n3969 = ~x2 & ~n1164 & (x0 ? n683 : n2438);
  assign n3970 = n742 & (n3971 | (x1 & ~n3972));
  assign n3971 = x7 & x4 & ~x1 & ~x3;
  assign n3972 = x3 ? (x4 | ~x7) : (~x4 | x7);
  assign n3973 = ~n643 & ((n1209 & n959) | (n1310 & ~n1062));
  assign n3974 = x1 | (~n3975 & ~n3976 & (~x4 | n3978));
  assign n3975 = x5 & ((n2492 & n995) | (n1181 & n2765));
  assign n3976 = ~x5 & ~n3977;
  assign n3977 = x0 ? (~x7 | (x2 ? (x3 | ~x4) : (~x3 | x4))) : (x7 | (x2 ? (~x3 ^ ~x4) : (x3 | ~x4)));
  assign n3978 = (x5 | n3979) & (~x3 | ~x5 | ~n742 | n640);
  assign n3979 = (x0 | x2 | ~x3 | ~x6 | x7) & (~x0 | ((x6 | x7 | x2 | x3) & (~x2 | ~x3 | (~x6 ^ ~x7))));
  assign z189 = n3981 | n3984 | ~n3988 | (x2 & ~n3987);
  assign n3981 = ~n1794 & (n3983 | (~x2 & ~n3982));
  assign n3982 = (~x1 & ((x5 & x6 & x7) | (x4 & ~x5 & ~x6 & ~x7))) | (x1 & (~x4 | x5) & (x6 ^ x7)) | (~x4 & x5 & (~x6 | ~x7)) | (x6 & x7 & (x4 ^ ~x5));
  assign n3983 = ~x1 & x2 & ((x5 & x6) | (~x4 & (x5 | x6)));
  assign n3984 = ~x4 & (n3985 | (n1300 & n1451 & n746));
  assign n3985 = ~x6 & ((n733 & n1453) | (n619 & ~n3986));
  assign n3986 = x0 ? (x2 ? (x3 | x5) : (~x3 | ~x5)) : (x3 | (~x2 ^ ~x5));
  assign n3987 = (~x3 | ~n592 | ~x0 | x1) & (x0 | (x1 ? ~n728 : (x3 | ~n592)));
  assign n3988 = n3992 & ~n3991 & ~n3989 & ~n3990;
  assign n3989 = n1250 & (x1 ? (x4 & n1723) : (~x4 & ~n1198));
  assign n3990 = ~n1134 & (n1644 | (~x0 & x1 & ~n2726));
  assign n3991 = ~n2259 & (n1783 | n2534);
  assign n3992 = (~n931 | ~n2534) & (~n959 | ~n816);
  assign z190 = n4000 | ~n4008 | (x3 ? ~n4004 : ~n3994);
  assign n3994 = ~n3995 & ~n3998;
  assign n3995 = ~x1 & ((n942 & n3996) | (~x4 & ~n3997));
  assign n3996 = x4 & x0 & x2;
  assign n3997 = (x0 | x2 | ~x6 | x7) & (~x7 | ((x0 | ~x2 | ~x5 | x6) & (~x0 | x5 | (~x2 ^ x6))));
  assign n3998 = x1 & (x0 ? (n1518 & n943) : ~n3999);
  assign n3999 = (x6 | x7 | ~x4 | ~x5) & (x4 | (x2 ? (~x6 | (~x5 ^ x7)) : (x6 | ~x7)));
  assign n4000 = ~n1097 & ((~x1 & ~n4001) | ~n4003 | (x1 & ~n4002));
  assign n4001 = x0 ? ((~x4 | ~x7 | x2 | x3) & (x4 | x7 | ~x2 | ~x3)) : ((x3 | ~x4 | x7) & (x2 | ~x7 | (~x3 ^ ~x4)));
  assign n4002 = (~x0 | x2 | x3 | x4 | ~x7) & (x0 | ((~x2 | ~x3 | ~x4 | x7) & (x2 | x4 | (~x3 ^ ~x7))));
  assign n4003 = x1 ? ((x3 | ~x4 | ~x0 | x2) & (x0 | ~x3 | (~x2 ^ x4))) : (x0 ? (x2 ? (x3 | ~x4) : (~x3 | x4)) : (~x2 | (~x3 ^ ~x4)));
  assign n4004 = x1 ? (x0 | n4007) : (~n4005 & ~n4006);
  assign n4005 = ~n1100 & (x0 ? n572 : n3517);
  assign n4006 = n1084 & ~x0 & n1070;
  assign n4007 = (x2 | ~x4 | ~x5 | x6 | ~x7) & (~x2 | ~x6 | (x4 ? (~x5 | ~x7) : (x5 | x7)));
  assign n4008 = x0 ? (~n4009 & (x1 | n4013)) : n4010;
  assign n4009 = n704 & n576;
  assign n4010 = x1 ? (x4 ? n4011 : n2511) : (n4012 & (~x4 | n2511));
  assign n4011 = (x3 | x5 | ~x6) & (~x2 | ~x3 | ~x5 | x6);
  assign n4012 = (~x2 | ~x3 | x4 | x5 | ~x6) & (x2 | ~x5 | x6 | (x3 ^ ~x4));
  assign n4013 = x3 ? ((~x4 | ~x5 | x6) & (~x2 | ((~x4 | x5 | ~x6) & (~x5 | x6)))) : ((x2 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (x5 | ~x6 | ~x2 | x4));
  assign z191 = ~n4025 | n4021 | n4017 | n2235 | n4015;
  assign n4015 = ~x5 & (x1 ? ~n4016 : ~n2220);
  assign n4016 = (x2 | ((x3 | ~x4 | ~x6) & (x4 | x6 | ~x0 | ~x3))) & (x0 | ((x2 | ~x4 | ~x6) & (~x2 | x3 | x4 | x6)));
  assign n4017 = ~x0 & (n4018 | (n1044 & ~n4020));
  assign n4018 = x2 & ((n1070 & n3194) | (n2332 & ~n4019));
  assign n4019 = (x1 | ~x3 | ~x6 | x7) & (~x1 | (x3 ? (x6 | x7) : (~x6 | ~x7)));
  assign n4020 = (~x1 | x4 | ~x5 | x6 | ~x7) & (x5 | ((x1 | ~x4 | x6 | ~x7) & (~x1 | x7 | (~x4 ^ x6))));
  assign n4021 = ~n1218 & (~n4023 | (~x2 & ~n4022));
  assign n4022 = (x0 | x1 | ~x3 | ~x5 | ~x6) & (x6 | (~x1 ^ ~x5) | (x0 ^ ~x3));
  assign n4023 = x3 ? (x5 | n1184) : ((~x5 | n1184) & (~n570 | n4024));
  assign n4024 = x0 ? (x5 | ~x6) : (~x5 ^ ~x6);
  assign n4025 = n4028 & (~x5 | (~n4027 & (x0 | n4026)));
  assign n4026 = (x1 | x2 | ((~x4 | x6) & (x3 | x4 | ~x6))) & (~x2 | ~x3 | (x1 ? (~x4 ^ x6) : (~x4 | ~x6)));
  assign n4027 = n841 & ((n902 & n597) | (x2 & n1835));
  assign n4028 = (~n610 | ~n2144) & (n647 | n4029);
  assign n4029 = (~x0 | x1 | ~x2 | ~x6 | x7) & (x0 | x2 | ~x7 | (~x1 ^ x6));
  assign z192 = n4031 | ~n4045 | (x4 ? ~n4043 : ~n4038);
  assign n4031 = ~x2 & (n4036 | (~x0 & (n4032 | ~n4034)));
  assign n4032 = x1 & (n4033 | (x3 & ~n3345));
  assign n4033 = ~x3 & ~x5 & x7 & (x4 ^ x6);
  assign n4034 = (~n530 | ~n944) & (n1097 | n4035);
  assign n4035 = (x4 | x7 | ~x1 | x3) & (x1 | ~x3 | ~x7);
  assign n4036 = x0 & (x1 ? (n1392 & n942) : ~n4037);
  assign n4037 = x3 ? (x5 ? (~x6 | x7) : ((x6 | x7) & (~x4 | ~x6 | ~x7))) : ((x4 | ~x5 | ~x6 | ~x7) & (~x4 | x6 | (~x5 & ~x7)));
  assign n4038 = ~n4041 & (x0 | n4039) & (n3924 | n4040);
  assign n4039 = (x2 | (x1 ? (~x5 | ~x7) : ((~x5 | x7) & (x3 | x5 | ~x7)))) & (~x1 | ~x2 | x5 | (~x3 ^ ~x7));
  assign n4040 = x0 ? (~x1 | x2) : (x1 | ~x2);
  assign n4041 = n841 & (n4042 | (n750 & n885));
  assign n4042 = ~x3 & (~x5 ^ ~x7);
  assign n4043 = n4044 & (n1008 | (~n1270 & ~n2535));
  assign n4044 = x0 ? (~n632 | ~n1545) : (n3924 | (~n570 & ~n632));
  assign n4045 = ~n4046 & (~x2 | (n4051 & (x1 | n4048)));
  assign n4046 = ~n1198 & ((n1317 & ~n4047) | (~x1 & ~n2247));
  assign n4047 = (x4 | x7 | ~x0 | x2) & (x0 | (x2 ? ~x7 : (~x4 | x7)));
  assign n4048 = (x0 | ~x3 | ~n4050) & (x3 | (~n4049 & (~x0 | n3409)));
  assign n4049 = ~x7 & x6 & ~x5 & ~x0 & x4;
  assign n4050 = x5 & (x4 ? (x6 & ~x7) : (~x6 & x7));
  assign n4051 = (~n866 | ~n2402) & (n1097 | n4052);
  assign n4052 = (x0 | ~x1 | x7 | (~x3 ^ x4)) & (~x0 | x1 | ~x3 | ~x7);
  assign z193 = n4069 | n4065 | n4062 | n4054 | n4059;
  assign n4054 = ~n640 & (~n4056 | (~x1 & ~n4055));
  assign n4055 = (x0 | ~x2 | ~x3 | ~x4 | x5) & (~x5 | ((x0 | ~x2 | ~x3 | x4) & (x3 | (x0 ? (~x2 ^ ~x4) : (x2 | ~x4)))));
  assign n4056 = ~n4057 & ~n4058 & (~n731 | ~n733);
  assign n4057 = ~x1 & ((x0 & (x2 ? (x3 & ~x4) : (~x3 & x4))) | (~x0 & ~x2 & x3 & ~x4));
  assign n4058 = ~x4 & ~x3 & x2 & ~x0 & x1;
  assign n4059 = x4 & ((n1269 & n2939) | (~x5 & ~n4060));
  assign n4060 = (x2 | n4061) & (x0 | ~x2 | ~n1769 | n2085);
  assign n4061 = (~x0 | ((x1 | ~x3 | ~x6 | x7) & (~x1 | x3 | x6 | ~x7))) & (x0 | ~x1 | x3 | ~x6 | x7);
  assign n4062 = ~n643 & ((n1156 & ~n4064) | (~x2 & ~n4063));
  assign n4063 = x0 ? ((x1 | ~x3 | ~x4 | ~x5) & (~x1 | x3 | x4)) : ((x4 | x5 | x1 | x3) & (~x1 | (x3 ? (x4 | x5) : (~x4 | ~x5))));
  assign n4064 = (x1 | x3 | x5) & (x0 | (~x1 ^ ~x3));
  assign n4065 = ~x6 & (n4067 | ~n4068 | (~n714 & ~n4066));
  assign n4066 = (~x0 | x1 | ~x2 | x3) & (x0 | x2 | (~x1 ^ ~x3));
  assign n4067 = ~n647 & ~n4040;
  assign n4068 = (~n1287 | ~n560) & (~n731 | ~n746);
  assign n4069 = x6 & (n2294 | n2330 | (~n1685 & ~n1682));
  assign z194 = n4071 | n4073 | ~n4079 | (~n1205 & ~n4078);
  assign n4071 = ~x0 & ((n558 & n809) | (x1 & ~n4072));
  assign n4072 = x2 ? ((x3 | ~x4 | ~x5 | x7) & (~x3 | x4 | x5 | ~x7)) : ((~x4 | ~x5 | ~x7) & (x3 | x4 | x7));
  assign n4073 = ~x6 & (n4074 | ~n4076);
  assign n4074 = x4 & ((n1453 & n816) | (n757 & ~n4075));
  assign n4075 = (x2 | x3 | ~x0 | ~x1) & (x0 | ~x2 | (~x1 ^ ~x3));
  assign n4076 = (n4077 | n2223) & (~n526 | ~n774 | ~n816);
  assign n4077 = x2 ? (x3 | ~x5) : (~x3 | x5);
  assign n4078 = (~x0 | ~x1 | x2 | x4 | x5) & (x1 | ((x4 | x5 | x0 | ~x2) & (~x5 | (x0 ? (~x2 ^ ~x4) : (x2 | ~x4)))));
  assign n4079 = ~n4080 & ~n4083 & n4084 & (~n2570 | n4082);
  assign n4080 = ~n671 & ~n4081;
  assign n4081 = x0 ? ((x1 | ~x2 | ~x3 | x5) & (~x1 | x2 | x3 | ~x5)) : ((x1 | x2 | x5) & (~x2 | (x1 ? (~x3 ^ ~x5) : (x3 | ~x5))));
  assign n4082 = (x0 | ~x1 | ~x2 | ~x3 | x7) & (x2 | ((~x0 | (x1 ? (x3 | x7) : (~x3 | ~x7))) & (x0 | ~x1 | x3 | ~x7)));
  assign n4083 = ~n877 & ((~n3703 & n3396) | (n1209 & n1395));
  assign n4084 = (n714 | n4085) & (~n895 | (n3266 & ~n2992));
  assign n4085 = (~x2 | x3 | x7 | ~x0 | x1) & (x0 | ~x3 | (x1 ? (x2 | x7) : (~x2 | ~x7)));
  assign z195 = n4092 | n4094 | ~n4097 | (x6 & ~n4087);
  assign n4087 = x2 ? (~n4088 & (n814 | n2017)) : n4090;
  assign n4088 = n551 & ((n536 & n4089) | (n653 & n1379));
  assign n4089 = ~x4 & x7;
  assign n4090 = (~n2296 | ~n866) & (~x5 | n4091);
  assign n4091 = (~x1 | x3 | ~x4 | x7) & (x1 | ~x3 | (x0 ? (~x4 | x7) : (x4 | ~x7)));
  assign n4092 = ~x5 & ((n1209 & n745) | (~x4 & ~n4093));
  assign n4093 = x1 ? ((x3 | ~x6 | ~x0 | x2) & (x0 | ~x2 | (~x3 ^ ~x6))) : ((~x3 | (x0 ? (~x2 ^ x6) : (x2 | x6))) & (x3 | ~x6 | x0 | ~x2));
  assign n4094 = n706 & (x1 ? ~n4096 : ~n4095);
  assign n4095 = x0 ? ((~x2 | x3 | ~x4 | ~x7) & (x2 | ~x3 | x4 | x7)) : ((~x4 | ~x7 | x2 | x3) & (~x2 | (x3 ? (~x4 | ~x7) : (x4 | x7))));
  assign n4096 = (~x0 | x2 | x3 | x4 | x7) & (x0 | ~x3 | (x2 ? (x4 | x7) : (~x4 | ~x7)));
  assign n4097 = n4101 & (n4098 | n4099) & (x0 | ~n4100);
  assign n4098 = x4 ? (x5 ^ ~x6) : (x5 | x6);
  assign n4099 = (x0 | ~x2 | (~x1 ^ ~x3)) & (x2 | ((~x1 | x3) & (~x0 | x1 | ~x3)));
  assign n4100 = x1 & ((x2 & ~x3 & x4 & ~x5) | (~x2 & x3 & ~x4 & x5));
  assign n4101 = (x1 | n4102) & (~x6 | ~n1121 | n4103);
  assign n4102 = (x0 | ~x3 | (x2 ? (x4 | ~x5) : (~x4 | x5))) & (x3 | x4 | ~x5 | (~x0 & x2));
  assign n4103 = (x0 | ~x1 | x2 | ~x3) & (x1 | (x0 ? (~x2 | x3) : (~x2 ^ ~x3)));
  assign z196 = n4113 | ~n4115 | (x0 ? ~n4109 : ~n4105);
  assign n4105 = ~n4108 & (~n1498 | ~n2402) & (~x3 | n4106);
  assign n4106 = (~x6 | n4107) & (~x1 | ~n813 | ~n1084);
  assign n4107 = x1 ? ((~x5 | ~x7 | ~x2 | ~x4) & (x2 | (x4 ? (~x5 | x7) : (x5 | ~x7)))) : ((~x5 | ~x7 | x2 | x4) & (x5 | x7 | ~x2 | ~x4));
  assign n4108 = ~n1532 & ((n942 & n927) | (n689 & n943));
  assign n4109 = ~n4110 & (~n1467 | n4112);
  assign n4110 = x5 & ((~n643 & ~n2137) | (x7 & ~n4111));
  assign n4111 = (~x1 | x2 | x3 | ~x4 | ~x6) & (x1 | ((x2 | ~x4 | (~x3 ^ ~x6)) & (x4 | ~x6 | ~x2 | ~x3)));
  assign n4112 = (x6 | x7 | x3 | x4) & (~x6 | (x2 ? (~x7 | (~x3 ^ ~x4)) : (x7 | (x3 ^ ~x4))));
  assign n4113 = x6 & (x0 ? (n1716 & n570) : ~n4114);
  assign n4114 = (x3 | x5 | ~x1 | x2) & (x4 | (x1 ? ((x3 | x5) & (~x2 | ~x3 | ~x5)) : (x2 ? (x3 | ~x5) : (~x3 | x5))));
  assign n4115 = ~n4118 & ((x6 & (x3 | n4120)) | (n4116 & (n4120 | (~x3 & ~x6))));
  assign n4116 = (~x4 & (~x5 | (~n661 & ~n802))) | (n4117 & ((~n661 & ~n802) | (x4 & x5)));
  assign n4117 = (~x0 | x1 | ~x2 | ~x3 | ~x5) & (x0 | ((~x2 | (x1 ? (x3 | ~x5) : (~x3 | x5))) & (x1 | x2 | (~x3 ^ ~x5))));
  assign n4118 = ~n1353 & (x5 ? (n626 & ~n2726) : ~n4119);
  assign n4119 = x0 ? (x2 | (~x1 ^ x3)) : (~x2 | (~x1 ^ ~x3));
  assign n4120 = (x5 | x7 | n3290) & (x0 | ~x5 | ~x7 | n4121);
  assign n4121 = x1 ? (x2 ^ ~x4) : (~x2 | ~x4);
  assign z197 = ~n4136 | ~n4134 | n4130 | n4123 | n4125;
  assign n4123 = ~x1 & ((n600 & n1241) | (n1769 & ~n4124));
  assign n4124 = (x2 | x3 | x5 | (~x0 & ~x4)) & (x0 | ((~x2 | x3 | x4 | ~x5) & (~x3 | ((~x4 | x5) & (x2 | x4 | ~x5)))));
  assign n4125 = ~n640 & (n4126 | n4128 | (~n1134 & ~n4119));
  assign n4126 = ~x1 & ~n4127;
  assign n4127 = (~x0 | ((x3 | ~x4 | x5) & (x4 | ~x5 | ~x2 | ~x3))) & (x2 | x3 | ~x4 | x5) & (x0 | ~x3 | (x2 ? (~x4 | x5) : (x4 | ~x5)));
  assign n4128 = n543 & ((n2332 & n596) | (~x2 & ~n4129));
  assign n4129 = x3 ? (~x4 | x5) : ~x5;
  assign n4130 = ~n1134 & (n4132 | n4133 | (n543 & ~n4131));
  assign n4131 = x2 ? (x3 | x7) : (~x3 | ~x7);
  assign n4132 = ~x1 & ((~x0 & ~x2 & x3 & ~x7) | (x0 & x2 & (x3 ^ x7)));
  assign n4133 = n1910 & (x3 ? x2 : ~x1);
  assign n4134 = (n1934 | n4135) & (~n526 | ~n828 | ~n837);
  assign n4135 = (~x3 | ~x7 | ~x0 | x1) & (x0 | x7 | (~x1 ^ ~x3));
  assign n4136 = x7 ? (~n4137 | n4140) : n4138;
  assign n4137 = x1 & ~x6;
  assign n4138 = (x1 | n4139) & (~n1195 | (x0 & ~x4));
  assign n4139 = (x0 | ~x2 | ~x3 | x4 | ~x5) & (~x0 | ((x3 | x4 | ~x5) & (x2 | ~x3 | ~x4 | x5)));
  assign n4140 = (~x3 | x4 | x5 | ~x0 | x2) & (x0 | ((~x2 | (x3 ? (x4 | ~x5) : (~x4 | x5))) & (x4 | ~x5 | x2 | x3)));
  assign z198 = (x2 & ~n4154) | (~x2 & ~n4142) | (~n643 & ~n4151);
  assign n4142 = n4148 & n4147 & ~n4146 & ~n4143 & ~n4145;
  assign n4143 = ~x3 & ((n841 & ~n3409) | (n543 & ~n4144));
  assign n4144 = (~x6 | ~x7 | ~x4 | x5) & (x4 | x7 | (x5 ^ ~x6));
  assign n4145 = ~n1134 & ((n626 & n3903) | (x0 & n3050));
  assign n4146 = ~x0 & ((n689 & n3790) | (x1 & n2834));
  assign n4147 = (~n662 | ~n866) & (~n661 | (~n577 & ~n3790));
  assign n4148 = (x0 | n4149) & (n714 | n4150);
  assign n4149 = (x1 | x3 | x4 | ~x5 | ~x6) & (~x1 | ~x4 | x6 | (~x3 ^ x5));
  assign n4150 = (~x0 | ~x6 | ~x7 | (x1 ^ ~x3)) & (x0 | x1 | ~x3 | x6 | x7);
  assign n4151 = ~n4153 & (n1566 | n3290) & (x4 | n4152);
  assign n4152 = (x0 | ~x1 | ~x3 | (~x2 ^ ~x5)) & (x1 | ((x2 | x3 | x5) & (~x0 | ((x3 | x5) & (x2 | ~x3 | ~x5)))));
  assign n4153 = n566 & ((n1301 & n570) | (x1 & ~n1916));
  assign n4154 = (x1 | n4155) & (x0 | ~x1 | n4157);
  assign n4155 = (x3 & ((~x4 & x5 & n2341) | (~x5 & n4156))) | (n4156 & (x4 ^ ~x5)) | (~x3 & ((x5 & n4156) | (x4 & ~x5 & n2341)));
  assign n4156 = x0 ? (~x6 | ~x7) : (x6 | x7);
  assign n4157 = x6 ? (x3 ? (~x4 | x5) : (x4 ? ~x5 : (x5 | ~x7))) : (x3 ? (x7 | (x4 & ~x5)) : (x4 | ~x5));
  assign z199 = n4168 | ~n4171 | (x0 ? ~n4159 : ~n4163);
  assign n4159 = ~n4160 & (~n576 | ~n610);
  assign n4160 = ~x1 & (x3 ? ~n4161 : ~n4162);
  assign n4161 = (x5 | ((~x2 | ~x4 | ~x6 | ~x7) & (x2 | (x4 ? (~x6 | x7) : (x6 | ~x7))))) & (x4 | ~x5 | ((x6 | x7) & (x2 | ~x6 | ~x7)));
  assign n4162 = (~x2 | x4 | x5 | ~x6 | ~x7) & (x2 | (x4 ? (x5 ? (~x6 | x7) : (~x6 ^ ~x7)) : (x5 ? (x6 | ~x7) : (~x6 | x7))));
  assign n4163 = x2 ? n4166 : (x1 ? n4164 : n4165);
  assign n4164 = (x3 | ~x4 | ~x5 | x6 | x7) & (~x3 | x4 | x5 | ~x6 | ~x7);
  assign n4165 = ((~x3 ^ ~x4) | (x5 ? (x6 | ~x7) : (~x6 | x7))) & (x3 | ~x4 | ~x5 | ~x6 | x7) & (~x3 | x4 | x5 | x6 | ~x7) & ((~x6 ^ ~x7) | (x3 ? (x4 | ~x5) : (~x4 | x5)));
  assign n4166 = (n990 | n2085) & (n1218 | n4167);
  assign n4167 = (~x1 | x3 | ~x5 | x6) & (x1 | ~x3 | x5 | ~x6) & ((~x5 ^ ~x6) | (~x1 ^ ~x3));
  assign n4168 = ~n643 & (x0 ? ~n4170 : ~n4169);
  assign n4169 = (~x1 | x2 | (x3 ? (x4 | ~x5) : (~x4 | x5))) & (~x2 | ((x4 | x5 | ~x1 | x3) & (~x4 | ~x5 | x1 | ~x3)));
  assign n4170 = (~x1 | x2 | x3 | ~x4 | x5) & (x1 | ~x2 | (x3 ? (~x4 ^ ~x5) : (x4 | ~x5)));
  assign n4171 = (n2063 | n4176) & (x2 | n4172) & (~x2 | n4175);
  assign n4172 = x0 ? n4173 : (~x1 | n4174);
  assign n4173 = (~x3 | ((x5 | x7 | ~x1 | x4) & (~x5 | ~x7 | x1 | ~x4))) & (~x1 | x3 | (x4 ? (~x5 | ~x7) : (~x5 ^ x7)));
  assign n4174 = (x5 | x7 | ~x3 | x4) & (~x5 | ~x7 | x3 | ~x4) & ((~x3 ^ ~x4) | (~x5 ^ x7));
  assign n4175 = (x3 | n1014 | x0 | ~x1) & (x1 | ((~x3 | n1014) & (~x0 | x3 | n2216)));
  assign n4176 = (~x0 | x1 | ~x2 | x3 | ~x4) & (~x1 | x2 | ((x3 | x4) & (x0 | ~x3 | ~x4)));
  assign z200 = n4182 | ~n4184 | ~n4192 | (~x1 & ~n4178);
  assign n4178 = x5 ? (x7 | n4181) : (~n4179 & ~n4180);
  assign n4179 = ~x6 & ((n743 & n2647) | (~n2466 & ~n1218));
  assign n4180 = n1300 & ((~x0 & x2 & ~x3 & x4) | (x0 & (x2 ? (x3 ^ ~x4) : (x3 & ~x4))));
  assign n4181 = (x0 | x2 | ~x3 | x4 | ~x6) & (~x0 | ~x2 | ((~x4 | x6) & (x3 | x4 | ~x6)));
  assign n4182 = ~x2 & ((n852 & n2712) | (~x3 & ~n4183));
  assign n4183 = x6 ? ((x0 | ~x4 | x5 | x7) & (x4 | ~x5 | ~x7)) : ((x0 | x4 | (~x5 ^ x7)) & (~x4 | (x0 ? (x5 | x7) : (~x5 | ~x7))));
  assign n4184 = ~n4185 & ~n4188 & n4190 & (n1408 | n4187);
  assign n4185 = ~x6 & ((n1209 & n1641) | (~x2 & ~n4186));
  assign n4186 = (x0 | ~x3 | (x1 ? (x4 | x5) : (~x4 | ~x5))) & (x4 | ~x5 | ~x0 | x3);
  assign n4187 = (~x0 | x1 | x2 | ~x3 | ~x5) & (x0 | ((~x2 | x3 | x5) & (~x1 | x2 | ~x3 | ~x5)));
  assign n4188 = ~n643 & ((~n2185 & ~n4189) | (~n1327 & n3522));
  assign n4189 = (x3 | ~x5) & (x1 | ~x3 | x5);
  assign n4190 = (n752 | n4191) & (~n1364 | ~n1029 | ~n1209);
  assign n4191 = (x0 | x1 | ~x2 | ~x5) & (~x0 | x2 | x5);
  assign n4192 = ~n4194 & (~n742 | n4193);
  assign n4193 = (~x3 | ~x4 | x5 | ~x6 | ~x7) & (x7 | ((x5 | x6 | x3 | x4) & (~x4 | (x3 ? (~x5 ^ ~x6) : (~x5 | x6)))));
  assign n4194 = ~n823 & (x2 ? ~n4195 : (n774 & n658));
  assign n4195 = (x3 | ~x4 | ~x5 | ~x6 | ~x7) & (~x3 | x4 | (x5 ? (x6 | ~x7) : (~x6 | x7)));
  assign z201 = n4208 | ~n4211 | (x0 ? ~n4197 : ~n4202);
  assign n4197 = x1 ? (~n1044 | ~n610) : (~n4198 & n4200);
  assign n4198 = ~x2 & (x3 ? (~x5 & ~n2803) : (x5 & n4199));
  assign n4199 = ~x6 & (~x4 ^ x7);
  assign n4200 = ~n4201 & (~n942 | (~n1044 & ~n1489));
  assign n4201 = x2 & ((x3 & ~x5 & x6 & x7) | (~x3 & x5 & ~x6 & ~x7));
  assign n4202 = x5 ? n4206 : (n4204 & (~x4 | n4203));
  assign n4203 = (x1 | x2 | ~x3 | ~x6 | x7) & (~x1 | ((~x6 | ~x7 | x2 | x3) & (x6 | x7 | ~x2 | ~x3)));
  assign n4204 = ~n4205 & (~n550 | ~n576) & (~n689 | ~n1668);
  assign n4205 = ~x4 & ((x1 & x3 & x6 & x7) | (~x1 & ~x7 & (x3 ^ x6)));
  assign n4206 = (x6 | x7 | n2528) & (~x7 | n4207);
  assign n4207 = x1 ? (~x2 | ~x4 | (~x3 ^ ~x6)) : (x4 | ((x3 | x6) & (x2 | ~x3 | ~x6)));
  assign n4208 = ~n1097 & (x1 ? ~n4210 : ~n4209);
  assign n4209 = x0 ? ((x3 | x4 | ~x7) & (~x2 | ~x3 | ~x4 | x7)) : (~x4 | ((~x3 | ~x7) & (x2 | x3 | x7)));
  assign n4210 = (~x0 | x2 | x3 | x4 | ~x7) & (x0 | ~x3 | ((x4 | x7) & (x2 | ~x4 | ~x7)));
  assign n4211 = ~n4212 & ~n4214 & ~n4218 & (~n1317 | n4217);
  assign n4212 = ~n1954 & ((n653 & n670) | (x0 & ~n4213));
  assign n4213 = (x5 | x7 | ~x3 | x4) & (~x5 | ~x7 | x3 | ~x4);
  assign n4214 = x3 & ((~n1008 & ~n4215) | (n1080 & ~n4216));
  assign n4215 = (x0 | (x1 ? (~x2 | ~x4) : x4)) & (x2 | ~x4 | ~x0 | x1);
  assign n4216 = (x4 | x5 | ~x0 | x1) & (~x4 | ~x5 | x0 | ~x1);
  assign n4217 = (~x0 | x2 | x4 | ~x5 | x7) & (x0 | ((x4 | ~x5 | ~x7) & (x5 | x7 | ~x2 | ~x4)));
  assign n4218 = ~n643 & (x5 ? ~n4219 : (n1317 & ~n2185));
  assign n4219 = (~x0 | x1 | ~x3 | x4) & (x0 | x3 | ~x4 | (x1 ^ ~x2));
  assign z202 = ~n4231 | n4229 | n4221 | n4225;
  assign n4221 = ~n1218 & (n4223 | ~n4224 | (x0 & ~n4222));
  assign n4222 = (~x1 | x2 | x3 | ~x5 | x6) & (x1 | ((~x5 | ~x6 | x2 | x3) & (~x2 | x6 | (~x3 ^ ~x5))));
  assign n4223 = ~x0 & x6 & (x1 ? (x2 ^ ~x5) : (x2 & ~x5));
  assign n4224 = x1 | x2 | (x0 ? ~n904 : ~n1519);
  assign n4225 = ~n671 & ((~n4226 & ~n4227) | (~x0 & ~n4228));
  assign n4226 = x0 ^ x6;
  assign n4227 = x1 ? (x2 | x3) : (x5 | (~x2 & ~x3));
  assign n4228 = (x1 | x2 | x3 | x5 | x6) & (~x5 | (x1 ? (x6 | (~x2 & ~x3)) : (x2 | ~x6)));
  assign n4229 = ~x2 & (x0 ? (n704 & n689) : ~n4230);
  assign n4230 = (x1 | ~x3 | x4 | ~x5 | x6) & (~x1 | ~x4 | (x3 ? (x5 | x6) : (~x5 | ~x6)));
  assign n4231 = ~n4234 & ~n4236 & n4238 & (~n596 | n4232);
  assign n4232 = (~n943 | ~n3222) & (~x6 | ~n1167 | n4233);
  assign n4233 = x1 ? (x5 | x7) : (~x5 | ~x7);
  assign n4234 = x3 & ((n610 & n1269) | (~n538 & ~n4235));
  assign n4235 = (x4 | x7 | ~x0 | x1) & (~x4 | ~x7 | x0 | ~x1);
  assign n4236 = ~x2 & ~n4237;
  assign n4237 = (x0 | x1 | ~x4 | x5 | ~x6) & (~x0 | x6 | (x1 ? (x4 | x5) : (~x4 | ~x5)));
  assign n4238 = (~n2940 | ~n3093) & (n4239 | ~n4240);
  assign n4239 = x0 ? (x4 | ~x6) : (~x4 ^ ~x6);
  assign n4240 = x5 & ~x1 & x2;
  assign z203 = n4249 | ~n4254 | (x0 ? ~n4252 : ~n4242);
  assign n4242 = x4 ? n4246 : n4243;
  assign n4243 = (n1097 | n4245) & (x1 | ~n4244) & (~x1 | ~n2907);
  assign n4244 = ~x2 & x6 & (x3 ? (x5 & x7) : (~x5 & ~x7));
  assign n4245 = (x1 | ~x2 | x3 | ~x7) & (~x1 | x2 | x7);
  assign n4246 = (x1 | n4247) & (~n4248 | (~n813 & ~n2153));
  assign n4247 = x2 ? ((~x3 | ~x5 | ~x6 | x7) & (x6 | ~x7 | x3 | x5)) : (~x3 | ~x7 | (~x5 ^ ~x6));
  assign n4248 = ~x3 & x1 & ~x2;
  assign n4249 = ~n1198 & ((n1084 & n4250) | (x4 & ~n4251));
  assign n4250 = (x1 ^ ~x7) & (~x0 ^ ~x3);
  assign n4251 = x7 ? ((x0 | ~x1 | x2 | ~x3) & (~x0 | (x1 ? (x2 | x3) : (~x2 | ~x3)))) : ((x1 | x2 | x3) & (x0 | (x1 ? (~x2 | ~x3) : x2)));
  assign n4252 = ~n1505 & (x1 | (~n4253 & (~x4 | n1635)));
  assign n4253 = ~n1097 & (~n1410 | (n902 & n4089));
  assign n4254 = ~n4257 & (~n543 | n4255) & (n1548 | n4256);
  assign n4255 = (x5 | ((x4 | x7 | ~x2 | x3) & (x2 | (x3 ? (~x4 | x7) : ~x7)))) & (~x2 | ~x5 | ~x7 | (~x3 ^ ~x4));
  assign n4256 = (x0 | ~x2 | ~x5 | (~x1 ^ ~x7)) & (x5 | ((x0 | ~x1 | ~x2 | x7) & (~x0 | (x1 ? (x2 | x7) : (~x2 | ~x7)))));
  assign n4257 = ~x1 & (~n4259 | (x2 & n4258));
  assign n4258 = ~x3 & ~x4 & ((x5 & ~x7) | (x0 & ~x5 & x7));
  assign n4259 = (~x0 | x2 | ~x3 | ~x5 | x7) & (x0 | ~x7 | (x2 ? (~x3 | x5) : (x3 | ~x5)));
  assign z204 = n4268 | ~n4271 | (x7 ? ~n4266 : ~n4261);
  assign n4261 = x3 ? n4264 : (~n4263 & (x4 | n4262));
  assign n4262 = (~x0 | ~x1 | x2 | x5 | ~x6) & (x0 | ~x5 | (x1 ? (~x2 | x6) : x2));
  assign n4263 = x4 & n570 & (x0 ? (x5 ^ ~x6) : (x5 & ~x6));
  assign n4264 = (~n577 | ~n746) & (x6 | n4265);
  assign n4265 = x0 ? (x2 | (x1 ? (x4 | x5) : (~x4 | ~x5))) : (~x2 | x5 | (~x1 ^ x4));
  assign n4266 = (~n3074 | n4267) & (~n774 | ~n1723 | ~n560);
  assign n4267 = (x1 | x2 | ~x3 | x4 | x5) & (x3 | ((x1 | ~x2 | ~x4 | ~x5) & (~x1 | (x2 ? (x4 | ~x5) : (~x4 | x5)))));
  assign n4268 = ~n640 & (n2369 | n4270 | n1265 | n4269);
  assign n4269 = n1287 & n746;
  assign n4270 = ~x1 & (x0 ? (~x2 & n1909) : (x2 & n1268));
  assign n4271 = n4272 & ~n4275 & (n643 | n4274);
  assign n4272 = (~x2 | x6 | n3495) & (~x6 | n4273);
  assign n4273 = (x1 | (x0 ? (x2 ? (~x3 | ~x4) : x3) : (x2 | ~x3))) & (x0 | x2 | ((~x3 | x4) & (~x1 | x3 | ~x4)));
  assign n4274 = (x0 | ((~x2 | ~x3 | ~x4) & (~x1 | x2 | x3 | x4))) & (x1 | ((~x0 | ~x2 | ~x3 | x4) & (x3 | ~x4 | x0 | x2)));
  assign n4275 = x7 & ((n761 & n746) | (~x3 & ~n4276));
  assign n4276 = (~x0 | ((x1 | ~x2 | ~x4 | x6) & (~x1 | x2 | x4 | ~x6))) & (x0 | x1 | x2 | x4 | x6);
  assign z205 = ~n4284 | (x4 ? ~n4278 : ~n4280);
  assign n4278 = (~n1188 | n4279) & (~n1769 | ~n1451 | ~n733);
  assign n4279 = x0 ? ((~x2 | x5 | ~x6 | x7) & (x2 | ~x5 | x6 | ~x7)) : ((x2 | ~x5 | ~x6 | ~x7) & (~x2 | x5 | (~x6 ^ ~x7)));
  assign n4280 = ~n4281 & (x2 | (~n4283 & (~n626 | ~n942)));
  assign n4281 = ~n1558 & ((n922 & n878) | (~x0 & ~n4282));
  assign n4282 = x1 ? (~x2 | ~x6) : (x2 | x6);
  assign n4283 = x0 & ((n813 & n1188) | (n530 & n1317));
  assign n4284 = ~n4285 & ~n4288 & n4292 & (x2 | n4291);
  assign n4285 = x5 & ((~x1 & ~n4286) | (~x0 & n4287));
  assign n4286 = (x0 | ~x2 | ~x4 | (~x3 ^ ~x7)) & ((~x3 ^ x7) | (x0 ? (~x2 | ~x4) : (x2 | x4)));
  assign n4287 = x1 & ((~x2 & ~x3 & x4 & ~x7) | (~x4 & x7 & x2 & x3));
  assign n4288 = ~x5 & ((x0 & ~n4289) | (n742 & ~n4290));
  assign n4289 = (~x1 | x2 | x3 | x4 | x7) & (x1 | ~x4 | (x2 ? (x3 | x7) : (~x3 | ~x7)));
  assign n4290 = (x1 | x3 | ~x4 | ~x7) & (~x1 | x4 | (~x3 ^ x7));
  assign n4291 = (x0 | ~x1 | x4 | (~x3 ^ x7)) & (~x4 | ((x0 | x1 | x3 | ~x7) & ((~x1 ^ ~x7) | (x0 ^ ~x3))));
  assign n4292 = (n835 | n4294) & (~x2 | ~n626 | ~n4293);
  assign n4293 = ~x4 & (~x3 ^ ~x7);
  assign n4294 = (~x0 | x1 | x4) & (~x2 | ~x4 | x0 | ~x1);
  assign z206 = n4301 | ~n4308 | (x1 ? ~n4304 : ~n4296);
  assign n4296 = x6 ? n4299 : (~n4298 & (~x0 | n4297));
  assign n4297 = (x2 | ~x3 | x4 | x5 | x7) & (~x2 | ((~x5 | ~x7 | x3 | x4) & (x5 | x7 | ~x3 | ~x4)));
  assign n4298 = n1181 & ((n757 & n1029) | (~x3 & n2317));
  assign n4299 = (~n2296 | ~n2435) & (x2 | n4300);
  assign n4300 = (~x3 | ~x4 | ~x5 | x7) & (x3 | ~x7 | (x0 ? (x4 | ~x5) : (~x4 | x5)));
  assign n4301 = ~x0 & ((~x2 & ~n4303) | (~x1 & x2 & ~n4302));
  assign n4302 = (x3 | x4 | ~x5 | ~x6) & (x5 | x6 | ~x3 | ~x4);
  assign n4303 = (x1 | ~x3 | ~x4 | ~x5 | x6) & (x5 | ((x1 | x3 | x4 | ~x6) & (~x1 | (x3 ? (x4 | ~x6) : (~x4 | x6)))));
  assign n4304 = ~n4305 & (~n742 | n4307);
  assign n4305 = ~x2 & ((n566 & n4306) | (x0 & ~n985));
  assign n4306 = x6 & (x3 ? (x5 & x7) : (~x5 & ~x7));
  assign n4307 = (x3 | x4 | ~x5 | x6 | x7) & (~x3 | x5 | (x4 ? (x6 | ~x7) : (~x6 | x7)));
  assign n4308 = ~n4309 & ~n4312 & (x1 ? n4311 : n4314);
  assign n4309 = x0 & (x1 ? (n902 & n696) : ~n4310);
  assign n4310 = (x2 | ~x3 | ~x4 | ~x5 | x6) & (~x2 | x4 | ~x6 | (~x3 ^ x5));
  assign n4311 = (x0 | ~x2 | ~x4 | ~x5) & (x4 | ((x2 | x3 | x5) & (x0 | (x5 ? x2 : x3))));
  assign n4312 = ~n1353 & (n4313 | (~x5 & n825 & ~n3802));
  assign n4313 = x5 & ~x3 & ~x2 & x0 & x1;
  assign n4314 = x2 ? (x3 ? (x4 | ~x5) : (~x4 | x5)) : (~x4 | (x5 ? x3 : ~x0));
  assign z207 = n4316 | ~n4325 | (~x3 & ~n4322);
  assign n4316 = ~x2 & (n4319 | (~n4317 & ~n4318));
  assign n4317 = x0 ? (~x3 | x5) : (x3 | ~x5);
  assign n4318 = (~x1 | x4 | ~x6 | x7) & (x1 | (x4 ? (~x6 | ~x7) : (x6 | x7)));
  assign n4319 = ~x1 & (x6 ? (n1875 & n4321) : ~n4320);
  assign n4320 = (~x0 | ~x3 | x4 | ~x5 | ~x7) & (x0 | x5 | (x3 ? (~x4 | x7) : (x4 | ~x7)));
  assign n4321 = ~x7 & (x3 ^ ~x4);
  assign n4322 = ~n4324 & (n1100 | n4040) & (x5 | n4323);
  assign n4323 = (~x0 | x1 | x2 | ~x4 | ~x6) & (x0 | ((x1 | x4 | ~x6) & (x2 | ~x4 | x6)));
  assign n4324 = ~n823 & (x2 ? (~x5 & x6) : (x5 & (x4 ^ ~x6)));
  assign n4325 = ~n4328 & ~n4332 & (x2 ? n4326 : n4331);
  assign n4326 = (~n661 | ~n1626) & (n823 | n4327);
  assign n4327 = (~x3 | ~x4 | x5 | x6 | x7) & (x3 | ~x5 | (x4 ? (~x6 | ~x7) : (x6 | x7)));
  assign n4328 = x3 & (x4 ? ~n4330 : ~n4329);
  assign n4329 = (~x5 & x6) | (x5 & ~x6) | (x0 & (x1 ^ (~x2 & ~x6)));
  assign n4330 = (x0 | x1 | ~x2 | x5 | x6) & (~x5 | ((x0 | (~x2 ^ ~x6)) & (x1 | (x6 ? ~x2 : ~x0))));
  assign n4331 = (x0 | ~x3 | ~n4050) & (x3 | (~n4049 & (~x0 | n990)));
  assign n4332 = n742 & ((n1392 & n951) | (x3 & ~n3345));
  assign z208 = n4339 | n4342 | ~n4346 | (~x1 & ~n4334);
  assign n4334 = x0 ? (~n4338 & (~x5 | n4337)) : n4335;
  assign n4335 = (n1850 | n4336) & (~n1070 | ~n1556);
  assign n4336 = x2 ? (~x3 | x5) : (x3 | ~x5);
  assign n4337 = (x2 | x3 | x4 | x6 | ~x7) & (~x4 | ((x2 | x7 | (~x3 ^ ~x6)) & (~x2 | ~x3 | ~x6 | ~x7)));
  assign n4338 = n1429 & ((x4 & x6 & ~x2 & x3) | (~x3 & (x2 ? (x4 ^ ~x6) : (~x4 & x6))));
  assign n4339 = n632 & ((n1285 & n4341) | (~x0 & ~n4340));
  assign n4340 = (x3 | x4 | ~x5 | x6 | ~x7) & (~x3 | ~x4 | ~x6 | (~x5 ^ x7));
  assign n4341 = x7 & (~x4 | ~x5);
  assign n4342 = ~n640 & (n4343 | ~n4344);
  assign n4343 = ~n714 & (x0 ? (~x1 & x2) : ((x2 & ~x3) | (~x1 & ~x2 & x3)));
  assign n4344 = ~n4345 & (~n816 | ~n1311) & (x0 | ~n2003);
  assign n4345 = ~x2 & ((~x0 & x1 & x3 & ~x4) | (x0 & (x1 ? (~x3 & x4) : (x3 & ~x4))));
  assign n4346 = n4355 & ~n4353 & ~n4351 & ~n4347 & ~n4350;
  assign n4347 = ~x0 & ((~x1 & ~n4348) | (n1445 & ~n4349));
  assign n4348 = (x2 | ~x3 | x4 | x5 | x6) & (~x2 | x3 | ~x4 | ~x5 | ~x6);
  assign n4349 = (~x2 | ~x3 | ~x5 | x6) & (x2 | x3 | ~x6);
  assign n4350 = ~n1548 & ((n1209 & n943) | (n1291 & ~n790));
  assign n4351 = ~n823 & (n4352 | (x2 & ~n1113));
  assign n4352 = x7 & ~x6 & x5 & ~x2 & x4;
  assign n4353 = ~n4354 & ~x7 & n778;
  assign n4354 = (~x4 & (~x0 | (~x1 & ~x5))) | (x0 & x4) | (x1 & x5);
  assign n4355 = (~n1395 | ~n1885) & (~n560 | ~n3217);
  assign z209 = ~n4362 | ~n4375 | (x1 ? ~n4371 : ~n4357);
  assign n4357 = x3 ? n4358 : (x2 ? n4360 : n4361);
  assign n4358 = (~x5 | x6 | ~n564 | n3309) & (x5 | n4359);
  assign n4359 = (~x0 | ~x2 | x4 | x6 | x7) & (~x6 | ((x0 | x2 | ~x4 | ~x7) & (x7 | (x0 ? (~x2 ^ ~x4) : (~x2 | x4)))));
  assign n4360 = (~x4 | ~x6 | (x0 ? (~x5 ^ x7) : (x5 | x7))) & (x0 | x4 | x6 | (~x5 ^ ~x7));
  assign n4361 = (x0 | x5 | (x4 ? (x6 | ~x7) : (~x6 | x7))) & (~x5 | ((x4 | x6 | x7) & (~x0 | ~x4 | ~x6 | ~x7)));
  assign n4362 = ~n4368 & ~n4363 & ~n4366;
  assign n4363 = ~x2 & ((~x5 & ~n4364) | (~n1164 & n4365));
  assign n4364 = (x0 | ~x3 | ~x7 | (~x1 ^ ~x4)) & (x3 | ((~x0 | (x1 ? (x4 | x7) : (~x4 | ~x7))) & (x0 | ~x1 | x4 | ~x7)));
  assign n4365 = ~x7 & x5 & ~x0 & x3;
  assign n4366 = ~n643 & ((n1269 & n1641) | (~x2 & ~n4367));
  assign n4367 = (~x0 | x3 | x5 | (~x1 ^ ~x4)) & (~x3 | ((~x0 | x1 | ~x4 | x5) & (x0 | (x1 ? (x4 | x5) : (~x4 | ~x5)))));
  assign n4368 = ~x0 & ((~x6 & ~n4369) | (n1364 & ~n4370));
  assign n4369 = (x1 | x2 | ~x3 | ~x4 | x5) & (~x2 | ((~x1 | (x3 ? (~x4 | ~x5) : (x4 | x5))) & (x4 | ~x5 | x1 | ~x3)));
  assign n4370 = x1 ? (x2 | x4) : (~x4 | (~x2 ^ ~x3));
  assign n4371 = ~n4374 & (x0 | (~n4373 & (~x4 | n4372)));
  assign n4372 = (~x6 | ((~x2 | x3 | x5 | ~x7) & ((~x5 ^ ~x7) | (~x2 ^ ~x3)))) & (x3 | ~x5 | x6 | (~x2 ^ ~x7));
  assign n4373 = ~x7 & n2332 & (n1146 | n878);
  assign n4374 = n594 & n845;
  assign n4375 = ~n4378 & (n2803 | n4380) & (~x2 | n4376);
  assign n4376 = (x4 | n4377) & (x1 | ~x4 | ~n526 | n2129);
  assign n4377 = x0 ? (x1 | x3 | (~x5 ^ x7)) : (~x1 | ~x3 | (~x5 ^ ~x7));
  assign n4378 = x0 & ((n926 & n676) | (n691 & ~n4379));
  assign n4379 = (~x4 | ~x6 | x1 | ~x3) & (x3 | (x1 ? (~x4 ^ ~x6) : (~x4 ^ x6)));
  assign n4380 = x2 ? ((~x0 | x1 | ~x3 | x5) & (x0 | ((x3 | x5) & (x1 | ~x3 | ~x5)))) : (~x5 | (x0 ? (~x1 ^ x3) : (x1 | x3)));
  assign z210 = n4382 | n4386 | ~n4390 | (~n1701 & ~n4389);
  assign n4382 = ~x5 & (n4383 | n4385 | (n560 & n3497));
  assign n4383 = ~x0 & ((n1786 & n1439) | (x4 & ~n4384));
  assign n4384 = (x1 | ((x2 | x6 | x7) & (~x2 | x3 | ~x6 | ~x7))) & (x6 | x7 | ((x2 | x3) & (~x1 | ~x2 | ~x3)));
  assign n4385 = ~n1580 & ((n1300 & n1044) | (x2 & ~n3427));
  assign n4386 = ~n643 & (n4387 | n4388 | (n543 & n1622));
  assign n4387 = ~x1 & (x0 ? (x2 & n1909) : (~x2 & n1392));
  assign n4388 = ~n1998 & (x1 ? (x3 ? (~x4 & ~x5) : (x4 & x5)) : (x3 ? (x4 & x5) : (x4 ^ x5)));
  assign n4389 = x1 ? ((x3 | x4 | ~x0 | x2) & (x0 | (x2 ? (~x3 ^ ~x4) : (x3 | ~x4)))) : (x0 ? (x2 ? (x3 | ~x4) : (~x3 | x4)) : (x2 ? (~x3 | x4) : (~x3 ^ ~x4)));
  assign n4390 = ~n4395 & (x0 ? n4391 : (~n4393 & n4394));
  assign n4391 = x1 ? (~n1044 | ~n926) : n4392;
  assign n4392 = ((~x2 ^ ~x3) | (x4 ? (~x5 | ~x6) : (x5 | x6))) & (x2 | ~x3 | ~x4 | x5 | x6) & (~x2 | x3 | x4 | ~x6);
  assign n4393 = n3903 & ((n681 & n804) | (x1 & ~n2652));
  assign n4394 = x1 ? ((x3 | n2760) & (x2 | ~x3 | n2819)) : ((~x2 | x3 | n2819) & (~x3 | n2760));
  assign n4395 = ~n4396 & ~x6 & n691;
  assign n4396 = (x1 | ~x3 | ~x7 | (x0 ^ ~x4)) & (x3 | (~x1 ^ ~x4) | (~x0 ^ x7));
  assign z211 = x2 ? (~n4404 | ~n4411) : (~n4398 | ~n4407);
  assign n4398 = n4401 & (x3 | (~n4400 & (~x4 | n4399)));
  assign n4399 = x0 ? (~x5 | (x1 ? (~x6 | x7) : (x6 | ~x7))) : (x1 | x5 | (~x6 ^ x7));
  assign n4400 = n1445 & ((n1769 & n1380) | (x0 & n702));
  assign n4401 = (n627 | n4402) & (~n3436 | n4403);
  assign n4402 = (x0 | ~x1 | x4 | x5 | ~x7) & (x1 | ((x5 | x7 | x0 | x4) & (~x0 | (x4 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n4403 = (x1 | x4 | ~x5 | ~x7) & (~x4 | (x1 ? (~x5 ^ ~x7) : (~x5 | x7)));
  assign n4404 = ~n4406 & (~n588 | ~n661) & (n640 | n4405);
  assign n4405 = (x0 | x1 | (x3 ? (x4 | ~x5) : (~x4 | x5))) & ((~x3 ^ x5) | (x0 ? (x1 | ~x4) : (~x1 | x4)));
  assign n4406 = n3483 & ((n689 & n696) | (n559 & n927));
  assign n4407 = ~n4408 & ~n4409 & ~n4410 & (~n712 | ~n2209);
  assign n4408 = ~n1794 & (x1 ? ~n1337 : (~x5 & ~n671));
  assign n4409 = ~n2129 & ((~x5 & ~x7 & x1 & ~x4) | (~x1 & x5 & (x4 ^ x7)));
  assign n4410 = n566 & (x1 ? (~x3 & ~n765) : (x3 & n526));
  assign n4411 = ~n4412 & ~n4415 & n4417 & (n3146 | n1580);
  assign n4412 = n626 & (n4413 | n4414);
  assign n4413 = ~x7 & ~x5 & x3 & ~x4;
  assign n4414 = ~x3 & x5 & (x4 ^ ~x7);
  assign n4415 = ~n1008 & ((n774 & n841) | (~x0 & n4416));
  assign n4416 = x4 & (x1 ^ x3);
  assign n4417 = (x0 | ~x1 | ~x3 | ~x4 | x7) & (~x0 | x1 | x3 | x4 | ~x7);
  assign z212 = n4429 | ~n4432 | (x0 ? ~n4425 : ~n4419);
  assign n4419 = x1 ? n4420 : (~n4424 & (~x2 | n4423));
  assign n4420 = (~x3 | n4421) & (~n608 | ~n4422);
  assign n4421 = (x2 | x4 | x5 | ~x6 | ~x7) & (~x2 | x7 | (x4 ? x5 : (~x5 | x6)));
  assign n4422 = x7 & (~x4 | x5);
  assign n4423 = (x3 | ~x4 | ~x5 | x6 | x7) & (~x6 | ((~x3 | (x4 ? (~x5 | ~x7) : (x5 | x7))) & (x3 | x4 | x5 | ~x7)));
  assign n4424 = n691 & ((x3 & x4 & ~x6 & x7) | (~x3 & ~x7 & (~x4 ^ ~x6)));
  assign n4425 = ~n4428 & (x1 | n4426);
  assign n4426 = (x2 | ~x7 | n1100) & (x3 | (n4427 & (~x2 | x7 | n1100)));
  assign n4427 = (~x2 | x4 | x5 | x6 | ~x7) & (x2 | ~x4 | ~x5 | (~x6 ^ ~x7));
  assign n4428 = n576 & n1621;
  assign n4429 = x2 & ((~x0 & ~n4430) | (n841 & ~n4431));
  assign n4430 = x1 ? ((x3 | ~x4 | ~x5 | x6) & (~x3 | x4 | x5 | ~x6)) : ((~x3 | ~x4 | ~x5 | x6) & (x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))));
  assign n4431 = (x3 | x4 | x5 | ~x6) & (~x3 | ((~x5 | x6) & (~x4 | x5 | ~x6)));
  assign n4432 = ~n4437 & (n1097 | (n4434 & (x1 | n4433)));
  assign n4433 = x0 ? (x2 ? (x3 | ~x4) : (x4 | (x3 & ~x7))) : (~x3 | (x2 ? (x4 | x7) : (~x4 | ~x7)));
  assign n4434 = ~n4435 & (~n841 | ~n2047) & (~n1317 | n4436);
  assign n4435 = ~x0 & ((~x1 & x3 & ~x4 & x7) | (x4 & (x1 ? (x3 ^ ~x7) : (x3 & ~x7))));
  assign n4436 = x0 ? (x2 | (~x4 & ~x7)) : (~x2 | x4);
  assign n4437 = ~x2 & (x0 ? ~n4438 : ~n4439);
  assign n4438 = (x1 | ~x3 | ~x4 | ~x5 | x6) & (~x1 | x3 | x4 | x5 | ~x6);
  assign n4439 = x5 ? (x6 | ((x3 | x4) & (~x1 | (x3 & x4)))) : (~x6 | (x1 ? (~x3 | ~x4) : (x3 ^ ~x4)));
  assign z213 = ~n4455 | n4451 | n4447 | n4441 | n4444;
  assign n4441 = ~x2 & (x3 ? ~n4443 : ~n4442);
  assign n4442 = (x0 | ~x4 | (x1 ? (~x5 | x6) : (x5 | ~x6))) & ((~x1 ^ ~x6) | (x0 ? (~x4 | x5) : (x4 | ~x5)));
  assign n4443 = (~x0 | ~x1 | x4 | x5 | x6) & (~x4 | ((x0 | ~x1 | ~x5 | x6) & (x1 | (x0 ? (~x5 ^ ~x6) : (x5 | ~x6)))));
  assign n4444 = x2 & ((~x1 & ~n4445) | (n1291 & ~n4446));
  assign n4445 = (~x3 | ((~x5 | x6 | x0 | ~x4) & (~x0 | (x4 ? (x5 | ~x6) : (~x5 | x6))))) & (x0 | x4 | ((~x5 | ~x6) & (x3 | x5 | x6)));
  assign n4446 = (~x3 | ~x4 | x6) & (x4 | ~x6);
  assign n4447 = x2 & (n4448 | (n841 & ~n4450));
  assign n4448 = ~x0 & (x1 ? n4449 : (n774 & n658));
  assign n4449 = x4 & ((x6 & x7 & x3 & ~x5) | (~x6 & ~x7 & ~x3 & x5));
  assign n4450 = (~x3 | x4 | x5 | ~x6 | x7) & (x3 | ~x5 | (x4 ? (~x6 | x7) : (x6 | ~x7)));
  assign n4451 = ~n1218 & (n4453 | ~n4454 | (~x3 & ~n4452));
  assign n4452 = x0 ? ((~x1 | x2 | ~x5 | x6) & (x1 | ~x2 | x5 | ~x6)) : (~x2 | x6 | (~x1 ^ x5));
  assign n4453 = n825 & ((n1364 & n632) | (n527 & ~n968));
  assign n4454 = (~x0 | x1 | x2 | x5 | ~x6) & (x0 | ~x1 | (x2 ? (~x5 | ~x6) : (x5 | x6)));
  assign n4455 = ~n4463 & (n671 | (~n4456 & ~n4458 & n4459));
  assign n4456 = ~n1097 & (n829 | n4457);
  assign n4457 = x0 & (x1 ? (~x2 & ~x3) : (x2 & x3));
  assign n4458 = ~x0 & ~x5 & x6 & (~x1 ^ ~x2);
  assign n4459 = ~n4461 & (~n3848 | ~n1209) & (n4460 | ~n4462);
  assign n4460 = x1 ? (~x2 | x6) : (x2 | ~x6);
  assign n4461 = ~x6 & x5 & ~x2 & x0 & ~x1;
  assign n4462 = x5 & ~x0 & x3;
  assign n4463 = n4464 & ((n559 & n622) | (~x0 & n2851));
  assign n4464 = x7 & ~x1 & ~x2;
  assign z214 = ~n4479 | n4476 | ~n4472 | n4466 | n4468;
  assign n4466 = n632 & (x0 ? (n1392 & n942) : ~n4467);
  assign n4467 = x3 ? (~x5 | (x4 ? (x6 | x7) : (~x6 | ~x7))) : (x5 | x6 | (x4 ^ ~x7));
  assign n4468 = ~x1 & (n4469 | (~x6 & n1518 & ~n4471));
  assign n4469 = x6 & ((n594 & n809) | (~n4077 & ~n4470));
  assign n4470 = x0 ? (~x4 | ~x7) : (x4 | x7);
  assign n4471 = (x5 | x7 | ~x0 | x3) & (x0 | ~x7 | (~x3 ^ ~x5));
  assign n4472 = n4474 & (n1548 | n4473);
  assign n4473 = (~x0 | x1 | ~x2 | ~x5 | x7) & (x0 | ~x7 | (x1 ? (~x2 ^ ~x5) : (x2 | ~x5)));
  assign n4474 = (~x3 | x5 | ~n742 | n1543) & (x3 | n4475);
  assign n4475 = (x0 | ~x1 | x2 | ~x5 | x7) & (~x0 | ~x7 | (x1 ? (x2 | ~x5) : (~x2 | x5)));
  assign n4476 = ~n1097 & ((~n4477 & ~n3961) | (~x1 & ~n4478));
  assign n4477 = x2 ? (x3 | x4) : (~x3 | ~x4);
  assign n4478 = x0 ? ((x4 | x7 | x2 | x3) & (~x2 | ~x3 | ~x7)) : ((x4 | ~x7 | x2 | x3) & (~x2 | x7 | (~x3 ^ x4)));
  assign n4479 = ~n4480 & (n1198 | (~x1 & n4482) | (x1 & n4483));
  assign n4480 = ~x7 & ((n1287 & n1269) | (x3 & ~n4481));
  assign n4481 = (x4 | x5 | ~x0 | x2) & (x0 | ((~x1 | x2 | x4 | ~x5) & (x1 | ~x4 | (~x2 ^ ~x5))));
  assign n4482 = (x3 | (x0 ? (x2 | ~x7) : (~x2 ^ ~x7))) & (~x0 | ((x2 | x4 | ~x7) & (~x2 | ~x3 | ~x4 | x7)));
  assign n4483 = (~x0 | x2 | x3 | x4 | x7) & (x0 | ~x2 | (x3 ? (~x4 | ~x7) : x7));
  assign z216 = ~n4489 | n4485 | n4486;
  assign n4485 = ~x0 & ((n558 & n670) | (x1 & ~n668));
  assign n4486 = ~x3 & ((~n2996 & n4487) | (~n1218 & ~n4488));
  assign n4487 = x7 & ~x6 & ~x1 & ~x4;
  assign n4488 = x1 ? (x6 | ((x2 | x5) & (x0 | ~x2 | ~x5))) : (~x6 | (~x2 ^ ~x5));
  assign n4489 = n673 & ~n4490 & ~n4492 & (~n610 | ~n2534);
  assign n4490 = ~n1312 & ((n600 & n670) | (n1380 & ~n4491));
  assign n4491 = (x2 | ~x3 | ~x4 | x7) & (x4 | ~x7 | ~x2 | x3);
  assign n4492 = ~n671 & ((n570 & ~n4493) | (~x2 & ~n4494));
  assign n4493 = ~x3 & x5;
  assign n4494 = x1 ? (x3 | ~x5) : (~x3 | x5);
  assign z217 = n4500 | ~n4501 | (~x1 & ~n4496);
  assign n4496 = x0 ? (~n4499 & (~n1562 | ~n813)) : n4497;
  assign n4497 = x3 ? (~n4352 & (~n1156 | ~n942)) : n4498;
  assign n4498 = x2 ? ((~x6 | ~x7 | ~x4 | ~x5) & (x6 | x7 | x4 | x5)) : (~x4 | ~x6 | (~x5 ^ x7));
  assign n4499 = ~x3 & (x2 ? (x4 & n702) : (~x4 & n951));
  assign n4500 = ~n697 & ((n696 & n699) | (x4 & ~n3178));
  assign n4501 = ~n4504 & ~n4506 & (x2 | (~n4502 & n4503));
  assign n4502 = n551 & ((~x4 & ~x6 & ~x0 & ~x3) | (x0 & (x4 ? x6 : x3)));
  assign n4503 = (x3 | ((~x4 | ~x5 | x6) & (x4 | x5 | ~x6) & (~x0 | (~x5 ^ x6)))) & (x0 | ~x3 | ~x5 | (x4 & ~x6));
  assign n4504 = x2 & ((~n710 & ~n711) | (n681 & ~n4505));
  assign n4505 = (~x3 | ~x6 | x0 | ~x1) & (~x0 | x1 | (~x3 ^ ~x6));
  assign n4506 = n1317 & ((n530 & n3176) | (~x2 & ~n4507));
  assign n4507 = (~x4 | ~x5 | ~x6 | x7) & (x4 | x6 | (x0 ? (x5 | ~x7) : (~x5 | x7)));
  assign z218 = n4513 | ~n4517 | ~n4522 | (~x0 & ~n4509);
  assign n4509 = x1 ? (~n4511 & (x5 | n4510)) : n4512;
  assign n4510 = (x3 | ~x4 | ~x6 | ~x7) & (x7 | ((x2 | x3 | (~x4 ^ x6)) & (~x3 | (x2 ? (x4 | x6) : (~x4 | ~x6)))));
  assign n4511 = x7 & n3151 & ((x4 & x6) | (~x2 & ~x4 & ~x6));
  assign n4512 = n740 & (~x4 | ~n1044 | n1701);
  assign n4513 = ~x1 & ((x3 & ~n4514) | n4515 | ~n4516);
  assign n4514 = (~x0 | ~x2 | ~x4 | x5 | x6) & (x2 | (x0 ? (x4 ? (~x5 | ~x6) : (x5 | x6)) : (x6 | (~x4 ^ x5))));
  assign n4515 = ~n1998 & (n747 | (~x3 & x6 & ~n714));
  assign n4516 = (x0 | x2 | x3 | x4 | ~x6) & (~x2 | ((~x4 | x6 | x0 | ~x3) & (~x0 | x4 | (~x3 ^ x6))));
  assign n4517 = ~n4519 & (n524 | n4518);
  assign n4518 = (~x1 | x2 | x3 | x6) & (x0 | ((x1 | ~x2 | ~x3 | ~x6) & (~x1 | x3 | x6)));
  assign n4519 = x1 & ((~x4 & ~n4520) | (n1477 & ~n4521));
  assign n4520 = (x2 | x3 | ~x6 | (~x0 & ~x5)) & (x0 | ((~x2 | x3 | ~x6) & (~x3 | x6 | (x2 & ~x5))));
  assign n4521 = (x3 | ~x6 | ~x0 | x2) & (x0 | ~x3 | x6);
  assign n4522 = ~n4523 & (~x0 | (~n4526 & ~n4527));
  assign n4523 = ~n643 & ((n1029 & ~n4525) | (~x1 & n4524));
  assign n4524 = ~x3 & ~x4 & ~x5 & (x0 ^ x2);
  assign n4525 = x0 ? (x1 | (~x2 ^ ~x5)) : (~x5 | (~x1 & x2));
  assign n4526 = ~x2 & (x1 ? ~n740 : (n1029 & n943));
  assign n4527 = x4 & n570 & (n2888 | n2302);
  assign z219 = n4543 | ~n4529 | n4539;
  assign n4529 = ~n4530 & ~n4533 & n4536 & (n1218 | n4535);
  assign n4530 = ~n1408 & ((n746 & n4531) | (~x1 & ~n4532));
  assign n4531 = ~x7 & ~x3 & ~x5;
  assign n4532 = (x0 | x2 | x3 | x5 | x7) & (~x3 | ((x0 | ~x2 | ~x5 | x7) & (~x0 | (x2 ? (x5 | x7) : (~x5 | ~x7)))));
  assign n4533 = ~x2 & ((n712 & n809) | (~x3 & ~n4534));
  assign n4534 = (~x7 | ((x4 | x5 | ~x0 | x1) & (x0 | ~x1 | (~x4 & x5)))) & (~x0 | x1 | x7 | (~x4 & ~x5));
  assign n4535 = x0 ? (x1 | (~x2 ^ (x3 & ~x5))) : ((x3 | ~x5 | x1 | x2) & (~x1 | (x2 ? (x3 | ~x5) : ~x3)));
  assign n4536 = (n1176 | n4537) & (x5 | ~n570 | n4538);
  assign n4537 = (x0 | x1 | (~x2 ^ x3)) & (~x1 | (x0 ? (x2 | x3) : (~x2 | ~x3)));
  assign n4538 = (~x4 | ~x7 | ~x0 | ~x3) & (x0 | ((x4 | ~x7) & (~x3 | ~x4 | x7)));
  assign n4539 = ~x0 & (n4540 | (x7 & n1835 & ~n4542));
  assign n4540 = x4 & (x5 ? (n570 & ~n3427) : ~n4541);
  assign n4541 = (~x1 | ((~x2 | x3 | ~x6 | ~x7) & (x2 | ~x3 | x6 | x7))) & (x1 | x2 | ~x6 | ~x7);
  assign n4542 = (x1 | x2 | ~x3 | x5) & (~x1 | (x2 ? x5 : (x3 | ~x5)));
  assign n4543 = n743 & ((n945 & n951) | (~x3 & ~n4544));
  assign n4544 = (~x1 | x4 | x5 | ~x6 | x7) & (~x7 | ((x1 | ~x4 | ~x5 | x6) & (~x1 | x5 | (~x4 ^ ~x6))));
  assign z220 = ~n4558 | ~n4553 | n4546 | n4551;
  assign n4546 = ~x2 & (n4547 | (n774 & ~n4550));
  assign n4547 = x4 & ((x0 & ~n4548) | (n825 & ~n4549));
  assign n4548 = (~x1 | x3 | ~x5 | ~x6 | ~x7) & (x1 | ((x6 | ~x7 | x3 | x5) & (~x3 | ~x6 | (~x5 ^ x7))));
  assign n4549 = (x1 | x5 | ~x6 | x7) & (~x1 | x6 | (~x5 ^ ~x7));
  assign n4550 = (~x0 | x1 | ~x5 | ~x6 | x7) & (x0 | ((x1 | ~x6 | (~x5 ^ ~x7)) & (x6 | ~x7 | ~x1 | ~x5)));
  assign n4551 = n885 & ((n813 & n3222) | (~x4 & ~n4552));
  assign n4552 = (x0 | ~x1 | x5 | ~x6 | x7) & (x1 | x6 | (x0 ? (~x5 ^ ~x7) : (x5 | ~x7)));
  assign n4553 = ~n4556 & (x1 ? n4555 : n4554);
  assign n4554 = (x2 | x3 | ~x6 | (x0 ^ ~x5)) & ((x0 ^ x5) | (~x2 ^ (x3 & ~x6)));
  assign n4555 = (x0 | ~x2 | x5 | x6) & (x2 | ((x5 | x6 | ~x0 | x3) & (x0 | ~x5 | (x3 & ~x6))));
  assign n4556 = ~n1548 & ((n742 & n4557) | (n942 & n837));
  assign n4557 = x5 & (x1 ? (x6 & x7) : (~x6 & ~x7));
  assign n4558 = x0 ? (x2 | n4561) : (~n4559 & ~n4560);
  assign n4559 = x4 & ((n1133 & n1322) | (n527 & ~n1515));
  assign n4560 = ~n605 & n828 & x1 & x6;
  assign n4561 = (x1 | x3 | ~x4 | ~x5 | x6) & (x4 | (x1 ? (x3 ? (x5 | x6) : (~x5 | ~x6)) : (x5 | (~x3 ^ ~x6))));
  assign z221 = ~n4574 | n4573 | n4570 | n4563 | n4567;
  assign n4563 = ~n643 & (~n4565 | (~x2 & ~n4564));
  assign n4564 = (x0 | ~x1 | x3 | x4 | ~x5) & (~x3 | ((~x0 | x4 | (x1 ^ ~x5)) & (x0 | x1 | ~x4 | x5)));
  assign n4565 = ~n932 & ~n4566 & (~n959 | ~n746);
  assign n4566 = ~x2 & ((~x0 & ~x1 & x3 & ~x4) | (x0 & x4 & (x1 ^ x3)));
  assign n4567 = ~n640 & ((x3 & ~n4568) | (~n2267 & n4569));
  assign n4568 = (x0 | ~x1 | x2 | (~x4 ^ x5)) & (x1 | ~x2 | x4 | (~x0 & x5));
  assign n4569 = x4 & ~x1 & ~x3;
  assign n4570 = x1 & (n4571 | n4572 | (n743 & n3575));
  assign n4571 = ~x0 & ((x4 & x6 & ~x2 & ~x3) | (x2 & (x3 ? (x4 & x6) : (~x4 & ~x6))));
  assign n4572 = ~n1685 & n653 & ~x5 & ~x6;
  assign n4573 = n1283 & (n2202 | (n530 & n828));
  assign n4574 = x1 | (n4575 & ~n4578 & (~n600 | ~n601));
  assign n4575 = x6 ? n4577 : n4576;
  assign n4576 = (~x4 | (~x2 ^ ~x3) | (x0 & ~x5)) & (x2 | ((x4 | x5 | ~x0 | ~x3) & (x0 | x3 | ~x5)));
  assign n4577 = (x0 | x2 | ~x3 | ~x4 | ~x5) & (x3 | ((~x2 | x4) & (~x0 | x5 | (~x2 & x4))));
  assign n4578 = x2 & ((n2857 & n658) | (x4 & ~n4579));
  assign n4579 = (~x0 | ((x3 | ~x5 | ~x6 | ~x7) & (~x3 | x5 | x6 | x7))) & (x0 | x3 | x5 | ~x6 | ~x7);
  assign z222 = n4592 | n4590 | n4581 | ~n4584;
  assign n4581 = ~x1 & (x4 ? ~n4582 : ~n4583);
  assign n4582 = x7 ? ((x3 | ~x5 | ~x0 | x2) & ((~x3 ^ ~x5) | (~x0 ^ ~x2))) : ((x3 | x5 | ~x0 | x2) & (x0 | (x2 ? (x3 | ~x5) : (~x3 | x5))));
  assign n4583 = (x0 | ~x2 | ~x3 | x5 | x7) & (x2 | ((~x5 | ~x7 | x0 | x3) & (~x0 | (x3 ? (~x5 | x7) : (x5 | ~x7)))));
  assign n4584 = ~n4585 & (x2 ? n4588 : n4589);
  assign n4585 = x3 & ((~n640 & ~n4586) | (n1632 & ~n4587));
  assign n4586 = (~x0 | x1 | ~x2 | ~x4 | x5) & (x0 | ~x5 | (x1 ? (x2 | ~x4) : (~x2 | x4)));
  assign n4587 = (x0 | ~x1 | ~x6 | x7) & (x6 | ~x7 | ~x0 | x1);
  assign n4588 = (~x4 | ~x7 | x0 | ~x3) & (x4 | ((x0 | ((x3 | ~x7) & (~x1 | ~x3 | x7))) & (x1 | ((x3 | ~x7) & (~x0 | ~x3 | x7)))));
  assign n4589 = (x0 | x1 | ~x3 | x4 | x7) & (~x4 | ((~x0 | x7 | (x1 ^ ~x3)) & (x0 | ~x1 | x3 | ~x7)));
  assign n4590 = x1 & ((n674 & n1783) | (~x2 & ~n4591));
  assign n4591 = (x0 | ~x3 | ~x4 | x5 | x7) & (x4 | (x0 ? (x5 | (x3 ^ ~x7)) : (~x5 | x7)));
  assign n4592 = ~x3 & (~n4594 | (~x1 & (n4006 | n4593)));
  assign n4593 = n1121 & ((n1769 & n1181) | (x0 & n2753));
  assign n4594 = (n4595 | n4596) & (~n601 | ~n733);
  assign n4595 = x1 ? (x6 | ~x7) : (~x6 | x7);
  assign n4596 = (x4 | ~x5 | ~x0 | x2) & (x0 | x5 | (~x2 ^ ~x4));
  assign z223 = n2806 | (~x2 & (~n2792 | ~n2802 | n4598));
  assign n4598 = ~x5 & (x4 ? ~n2800 : (n1769 & n866));
  assign z224 = n4600 | ~n4603 | ~n4606 | (~n765 & ~n4601);
  assign n4600 = x1 & (n2563 | n2833);
  assign n4601 = ~n4602 & (n1408 | n2457) & (~n560 | ~n3575);
  assign n4602 = ~x0 & ((n1133 & n3575) | (x4 & n1614));
  assign n4603 = (~n1931 | ~n4604) & (n1566 | n4605);
  assign n4604 = ~x6 & (x3 ^ ~x5);
  assign n4605 = (~x4 | ~x6 | ~x0 | x1) & (x0 | (x1 ? ((~x2 | x4 | ~x6) & (~x4 | x6)) : (x4 | x6)));
  assign n4606 = (x2 | n4607) & (x1 | (~n2831 & ~n4609));
  assign n4607 = (x4 | n4608) & (~x4 | ~x5 | ~n622 | n1312);
  assign n4608 = (~x0 | x1 | ~x5 | (~x3 ^ x6)) & (~x1 | ((x5 | x6 | ~x0 | x3) & (x0 | (x3 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n4609 = ~n2830 & ((x4 & ~x6 & n995) | (~x0 & (x4 | x6)));
  assign z225 = ~n4611 | (~x2 & n2839);
  assign n4611 = ~n2842 & ~n2848 & n4614 & (n671 | n4612);
  assign n4612 = (x2 | n4613) & (~n1723 | ~n626) & (~x2 | n2357);
  assign n4613 = (~x1 | (x0 ? (x3 | ~x6) : (~x3 | x6))) & (~x0 | x1 | (x3 ? ~x6 : (x5 | x6)));
  assign n4614 = (~n2851 | ~n895) & (~n543 | ~n559);
  assign z226 = ~n4621 | n4620 | n4618 | n2865 | n4616;
  assign n4616 = x0 & (n4617 | (n558 & n2402));
  assign n4617 = x7 & ((~n1198 & ~n1226) | (n558 & n1358));
  assign n4618 = ~n1097 & ((n560 & n2765) | (~x0 & ~n4619));
  assign n4619 = x7 ? x1 : (~x1 | (~x2 & ~x3 & ~x4));
  assign n4620 = n934 & ((x0 & ~x1 & (x3 ^ x7)) | (x1 & (x0 ? (~x3 & ~x7) : (x3 & x7))));
  assign n4621 = ~n4622 & ~n4623 & (~n845 | ~n3791);
  assign n4622 = ~x7 & ~x5 & x2 & x0 & ~x1;
  assign n4623 = ~x0 & ((~x1 & x5 & ~x7) | (~x5 & x7 & x1 & x2));
  assign z227 = n2876 | n4625 | (~n640 & ~n4626);
  assign n4625 = ~x2 & (n2869 | (n939 & ~n1935));
  assign n4626 = n4627 & (x0 | x4 | ~n1044 | n2290);
  assign n4627 = (x2 | x3 | ~x0 | ~x1) & (x1 | (~x2 & ~x3 & (x0 | ~x4)));
  assign z228 = x7 & (~n2732 | (n837 & n1203));
  assign z229 = ~n4631 | (x1 & ~n2373) | (n1093 & ~n4630);
  assign n4630 = (~x3 | x4 | x6 | ~x0 | x2) & (x0 | ~x2 | x3 | ~x4 | ~x6);
  assign n4631 = ~n841 & (~n830 | ~n4632) & (~n959 | ~n746);
  assign n4632 = x3 & ~x2 & x0 & x1;
  assign z230 = n4634 | n4635 | ~n4636 | (n742 & ~n2528);
  assign n4634 = x3 & ((n577 & n1269) | (n743 & ~n1335));
  assign n4635 = n774 & ((n943 & n1269) | (n942 & n837));
  assign n4636 = ~n880 & n1036 & (~n746 | ~n3217);
  assign z231 = ~n4638 | ~n4644 | (x3 & (n4641 | n4643));
  assign n4638 = n4640 & (x1 | n4639);
  assign n4639 = (~x0 | x2 | x3 | x4 | ~x5) & (~x3 | ((x0 | ~x2 | x4 | x5) & (~x4 | (x0 ? (~x2 ^ ~x5) : (x2 | ~x5)))));
  assign n4640 = (x0 | ~x2 | x3 | (x1 & x4)) & (x2 | ((~x1 | (x0 ^ ~x3)) & (~x0 | ((x3 | ~x4) & (x1 | ~x3 | x4)))));
  assign n4641 = ~x5 & ((n816 & n1668) | (x0 & ~n4642));
  assign n4642 = (x1 | ~x2 | ~x4 | x6 | ~x7) & (~x1 | x2 | x4 | ~x6 | x7);
  assign n4643 = n1269 & n993;
  assign n4644 = ~n4645 & (~n560 | ~n2145) & (~n662 | ~n3791);
  assign n4645 = ~x5 & ((n1331 & n746) | (n536 & ~n3207));
  assign z232 = ~n4648 | (x2 & (~n4647 | (n926 & n699)));
  assign n4647 = (x0 | (x1 ? (~x3 ^ ~x4) : (x3 | ~x4))) & (x1 | (x3 ? (x4 | (~x0 & x5)) : (~x4 | ~x5)));
  assign n4648 = ~n4656 & (x2 | (n4649 & n4651 & n4653));
  assign n4649 = n4650 & (~n1287 | ~n841) & (~n559 | ~n866);
  assign n4650 = (x0 | x1 | ~x3 | x4) & (~x0 | ~x1 | x3 | ~x4);
  assign n4651 = (n981 | n4652) & (n1682 | (n714 & n1040));
  assign n4652 = x0 ? (~x1 | x4) : (x1 | ~x4);
  assign n4653 = (n2786 | n4654) & (~n2446 | n4655);
  assign n4654 = x1 ? (~x6 | x7) : (x6 | ~x7);
  assign n4655 = (x1 | x5 | ~x6 | x7) & (~x1 | ~x5 | x6 | ~x7);
  assign n4656 = n885 & ((n4557 & n1167) | (n813 & n3222));
  assign z233 = ~n4666 | n4663 | n4658 | n4660;
  assign n4658 = ~x1 & ((~n1143 & ~n3190) | (~x4 & ~n4659));
  assign n4659 = (x0 | ~x2 | x3 | x5 | ~x6) & (~x0 | (x2 ? (~x6 | (~x3 ^ x5)) : (x3 | x5)));
  assign n4660 = x2 & (n4661 | (~x4 & n543 & n1293));
  assign n4661 = ~x1 & ((n530 & n1074) | (~x6 & ~n4662));
  assign n4662 = x0 ? ((~x5 | ~x7 | x3 | x4) & (x5 | x7 | ~x3 | ~x4)) : (x4 | (x3 ? (~x5 | x7) : (x5 | ~x7)));
  assign n4663 = ~x2 & ((~x7 & ~n4664) | (n1465 & ~n4665));
  assign n4664 = (~x4 | ~n825 | n899) & (n1312 | n2786);
  assign n4665 = (x0 | x1 | x4 | ~x5 | ~x6) & (~x4 | ((x0 | ~x1 | x5 | x6) & (~x0 | (x1 ? (~x5 | x6) : (x5 | ~x6)))));
  assign n4666 = ~n4667 & ~n4669 & ~n4670 & (n1011 | n4672);
  assign n4667 = ~n4668 & (x2 ? ~x4 : (x4 & ~x6));
  assign n4668 = (~x3 | ~x5 | ~x0 | x1) & (x0 | ((~x3 | x5) & (~x1 | x3 | ~x5)));
  assign n4669 = n1017 & ((x5 & x6 & ~x0 & x3) | (x0 & ~x5 & (~x3 | ~x6)));
  assign n4670 = ~n4671 & ((x1 & ~x4 & ~x6) | (x4 & (~x1 | x6)));
  assign n4671 = (x3 | ~x5 | ~x0 | x2) & (x0 | (x2 ? (~x3 | ~x5) : (x3 | x5)));
  assign n4672 = (~x0 | x1 | ~x4 | x5) & (x0 | (x1 ? (~x4 | x5) : (x4 | ~x5)));
  assign z234 = ~n4678 | n4682 | (x2 ? ~n4674 : ~n4685);
  assign n4674 = (x1 | n4676) & (x0 | (x1 ? n4677 : ~n4675));
  assign n4675 = ~x3 & x5 & (x4 ? (x6 & ~x7) : (~x6 & x7));
  assign n4676 = (n1035 | n3098) & (~x0 | ~n1029 | ~n813);
  assign n4677 = (~x3 | x4 | ~x5 | ~x6 | x7) & (x3 | ((x4 | ~x6 | (~x5 ^ ~x7)) & (x6 | ~x7 | ~x4 | ~x5)));
  assign n4678 = ~n4679 & (~x3 | (~n4681 & (x6 | n4680)));
  assign n4679 = ~n1100 & (n880 | (~x0 & (n558 | n927)));
  assign n4680 = (~x0 | x4 | x5 | (x1 ^ ~x2)) & (~x4 | (x0 ? (x1 | ~x5) : (x1 ? (~x2 | ~x5) : x5)));
  assign n4681 = n2315 & ((~x0 & ~x2 & x4 & x5) | ((x2 | ~x4) & (~x0 ^ x5)));
  assign n4682 = ~x3 & (x5 ? ~n4684 : ~n4683);
  assign n4683 = (~x0 | x1 | ~x4 | x6) & ((~x2 & x4) | (x0 ? (x1 | ~x6) : (~x1 | x6)));
  assign n4684 = (~x0 | x1 | x2 | ~x4 | ~x6) & (x0 | ((~x4 | ~x6 | ~x1 | ~x2) & ((x1 ^ ~x2) | (~x4 ^ x6))));
  assign n4685 = n4688 & (x0 | (n4686 & (~n772 | ~n2660)));
  assign n4686 = (~n1070 | ~n945) & (n1008 | n4687);
  assign n4687 = (x1 | x3 | x4 | ~x6) & (~x1 | ~x3 | ~x4 | x6);
  assign n4688 = x0 ? (x5 ? (x6 | n4689) : n4690) : (n4689 | (~x5 ^ ~x6));
  assign n4689 = (~x1 | x3 | ~x4 | x7) & (x1 | ~x3 | x4 | ~x7);
  assign n4690 = (x1 | ~x4 | ~x6 | (~x3 ^ ~x7)) & (x4 | (x3 ^ ~x7) | (x1 ^ x6));
  assign z235 = n4701 | ~n4706 | (x7 ? ~n4692 : ~n4697);
  assign n4692 = x2 ? n4693 : n4695;
  assign n4693 = (x3 | ~x4 | ~n841 | n1198) & (~x3 | n4694);
  assign n4694 = (x0 | ~x1 | (x4 ? (~x5 | x6) : (x5 | ~x6))) & (x1 | (~x4 ^ ~x6) | (x0 ^ x5));
  assign n4695 = (~n577 | ~n661) & (x6 | n4696);
  assign n4696 = (x0 | x1 | ~x3 | ~x4 | ~x5) & (x3 | ((x0 | x1 | x4 | ~x5) & (~x0 | (x4 ? x5 : ~x1))));
  assign n4697 = ~n4700 & (x0 | (~n4699 & (x1 | n4698)));
  assign n4698 = x2 ? (x4 | (x3 ? (x5 | x6) : (~x5 | ~x6))) : (~x4 | (x3 ? (~x5 ^ x6) : (x5 | x6)));
  assign n4699 = n632 & (n960 | (x3 & ~x4 & ~n1198));
  assign n4700 = n1209 & n960;
  assign n4701 = ~n640 & (~n4703 | ~n4704 | (~x0 & ~n4702));
  assign n4702 = (x1 | x2 | x3 | ~x4 | ~x5) & (~x3 | ((x1 | x4 | (~x2 ^ ~x5)) & (~x1 | ~x2 | ~x4 | ~x5)));
  assign n4703 = (n586 | n2227) & (~n1287 | ~n560);
  assign n4704 = ~n4705 & (n714 | (~n1644 & ~n3791));
  assign n4705 = ~x3 & ((~x0 & ~x1 & x2 & ~x4) | (x0 & x1 & ~x2 & x4));
  assign n4706 = ~n4707 & ~n4710 & ~n4711 & (n1113 | n1036);
  assign n4707 = ~x2 & ((n4708 & n951) | (~x4 & ~n4709));
  assign n4708 = x4 & ~x0 & ~x1;
  assign n4709 = (x0 | ((x1 | ~x6 | x7) & (x6 | ~x7 | ~x1 | ~x5))) & (~x6 | x7 | ((~x0 | ~x1 | x5) & (x1 | ~x5)));
  assign n4710 = n742 & ((n772 & n978) | (x1 & ~n2128));
  assign n4711 = ~n1116 & ((n742 & ~n2208) | (n1518 & n841));
  assign z236 = ~n4729 | n4726 | n4724 | n4713 | ~n4717;
  assign n4713 = x1 & (n4374 | n4714);
  assign n4714 = ~x0 & (x2 ? ~n4715 : ~n4716);
  assign n4715 = (~x3 | x6 | ~x7 | (~x4 ^ ~x5)) & ((x4 ? (x5 | ~x7) : (~x5 | x7)) | (x3 ^ x6));
  assign n4716 = (x6 | x7 | x4 | x5) & (~x7 | ((~x5 | ~x6 | ~x3 | ~x4) & (x3 | (x4 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n4717 = ~n4722 & (x1 | n4718) & (n2803 | n4721);
  assign n4718 = (n882 | n4719) & (~x6 | ~n1121 | n4720);
  assign n4719 = (x3 | ~x4 | ~x5 | ~x6 | x7) & (x4 | x6 | (x3 ? (~x5 ^ ~x7) : (x5 | ~x7)));
  assign n4720 = (x0 | ~x2 | ~x3 | x7) & (~x0 | x2 | ~x7);
  assign n4721 = x1 ? ((x3 | ~x5 | ~x0 | x2) & (x0 | x5 | (~x2 ^ ~x3))) : ((~x3 | (x0 ? (~x2 ^ x5) : (x2 | x5))) & (x3 | ~x5 | x0 | ~x2));
  assign n4722 = x2 & ((n674 & n699) | (~x1 & ~n4723));
  assign n4723 = ((~x3 ^ ~x5) | (x0 ? (~x4 | ~x7) : (x4 | x7))) & (~x0 | x3 | x4 | ~x5 | x7) & (x0 | ~x3 | x5 | ~x7);
  assign n4724 = ~n643 & ((n1287 & n746) | (x4 & ~n4725));
  assign n4725 = (x0 | x1 | ~x2 | x3 | x5) & (x2 | ((x0 | ~x1 | x3 | ~x5) & (~x0 | x5 | (~x1 ^ x3))));
  assign n4726 = ~x2 & (~n4728 | (~x1 & ~n4727));
  assign n4727 = (x5 | x7 | ~x0 | x4) & (x0 | ((~x5 | ~x7 | ~x3 | ~x4) & (x3 | (x4 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n4728 = (n1014 | n1119) & (~n2209 | ~n1734);
  assign n4729 = ~n4730 & (~n561 | ~n1209) & (n2208 | n4732);
  assign n4730 = x5 & ((n3575 & n1269) | (~x2 & ~n4731));
  assign n4731 = (x0 | ~x1 | ~x3 | ~x4 | x6) & (~x0 | ((~x1 | x3 | ~x4 | ~x6) & (x1 | ~x3 | x4 | x6)));
  assign n4732 = (~x0 | x2 | x3 | ~x5 | x6) & (x0 | ~x6 | (x2 ? (x3 | ~x5) : (~x3 | x5)));
  assign z237 = n4748 | n4743 | n4734 | ~n4737;
  assign n4734 = ~n643 & (n4067 | n4735 | (~x1 & ~n4736));
  assign n4735 = n543 & ((x2 & x4 & (x3 ^ ~x5)) | (~x4 & ((~x3 & x5) | (~x2 & x3 & ~x5))));
  assign n4736 = x3 ? ((~x0 ^ ~x2) | (~x4 ^ x5)) : ((x2 | x4 | x5) & (~x0 | ((x4 | x5) & (x2 | ~x4 | ~x5))));
  assign n4737 = x1 ? n4741 : (n4739 & (~x7 | n4738));
  assign n4738 = (x0 | ~x2 | ~x3 | x4 | ~x6) & (~x0 | x2 | (x3 ? (~x4 | x6) : ~x6));
  assign n4739 = (n2099 | n4156) & (n1532 | n4740);
  assign n4740 = (x0 | x3 | ~x6 | ~x7) & (x6 | x7 | ~x0 | ~x3);
  assign n4741 = (n2373 | n2803) & (x0 | n4742);
  assign n4742 = (x6 | x7 | x3 | x4) & (x2 | ~x4 | (x3 ? (~x6 | ~x7) : x6));
  assign n4743 = ~x1 & (n4744 | n4747 | (~n882 & ~n4746));
  assign n4744 = ~n4745 & ~x7 & n743;
  assign n4745 = (x3 | ~x4 | ~x5 | x6) & (x4 | (x3 ? (~x5 ^ x6) : (~x5 | ~x6)));
  assign n4746 = x3 ? ((~x4 | ~x5 | ~x6) & (x6 | ~x7 | x4 | x5)) : (x4 ? (x7 | (~x5 ^ x6)) : (~x5 | ~x6));
  assign n4747 = n742 & ((~n1026 & ~n1337) | (n1029 & n658));
  assign n4748 = x1 & (n4749 | (n1686 & ~n4751));
  assign n4749 = ~x6 & ((~n2373 & ~n1337) | (~x0 & ~n4750));
  assign n4750 = (x2 | ~x3 | ~x4 | ~x5 | x7) & (x5 | ~x7 | x3 | x4);
  assign n4751 = (~x4 | ~x5 | ~x2 | x3) & (x2 | ((~x3 | (x4 ? (x5 | x7) : ~x5)) & (x4 | ~x5 | ~x7)));
  assign z238 = ~n4756 | ~n4763 | (x6 ? ~n4761 : ~n4753);
  assign n4753 = ~n4755 & (~n895 | n4754) & (n1337 | n4066);
  assign n4754 = (x3 | ~x4 | ~x5 | x7) & (x5 | ~x7 | ~x3 | x4);
  assign n4755 = ~n1682 & ((n1156 & n1429) | (~x2 & n2316));
  assign n4756 = ~n4759 & (~x1 | (~n4757 & (~n2296 | ~n1783)));
  assign n4757 = ~x2 & ((~x0 & n1460) | (n1903 & ~n4758));
  assign n4758 = x0 ? (x4 | x5) : (~x4 | ~x5);
  assign n4759 = ~n643 & ((~n1134 & ~n4075) | (n2332 & ~n4760));
  assign n4760 = (x0 | (x1 ? (~x2 | x3) : (x2 | ~x3))) & (~x2 | ~x3 | ~x0 | x1);
  assign n4761 = (~n750 | ~n828 | ~n733) & (x1 | n4762);
  assign n4762 = (x4 | x5 | x7 | ~n547) & (n2373 | (x4 ? (~x5 ^ ~x7) : (x5 | ~x7)));
  assign n4763 = ~n4765 & (n1337 | n4119) & (n765 | n4764);
  assign n4764 = (x0 | ~x1 | (x2 ? (x3 | ~x4) : (~x3 | x4))) & (x1 | (x0 ? ((x3 | x4) & (~x2 | ~x3 | ~x4)) : (~x3 | (~x2 ^ x4))));
  assign n4765 = ~x1 & ((~n882 & ~n4754) | (n1380 & ~n3036));
  assign z239 = n4778 | ~n4783 | (x2 ? ~n4774 : ~n4767);
  assign n4767 = x0 ? n4768 : (~n4772 & (x5 | n4771));
  assign n4768 = x5 ? n4769 : n4770;
  assign n4769 = (~x1 | x3 | x4 | x6 | x7) & (x1 | ~x3 | ~x4 | ~x6 | ~x7);
  assign n4770 = x4 ? ((~x1 | x3 | ~x6 | x7) & (x1 | x6 | ~x7)) : ((~x3 | x6 | x7) & (x1 | (~x6 ^ ~x7)));
  assign n4771 = (x1 | x4 | (x3 ? (~x6 | x7) : (x6 | ~x7))) & (~x4 | ((x1 | ~x3 | x6 | x7) & (~x7 | (x1 ? (~x3 ^ ~x6) : (x3 | ~x6)))));
  assign n4772 = n2074 & ((n774 & n1769) | (~x3 & ~n4773));
  assign n4773 = x4 ? (~x6 | ~x7) : (x6 ^ ~x7);
  assign n4774 = ~n4777 & (x1 | (~n4776 & (x0 | n4775)));
  assign n4775 = (x7 | ((x5 | x6 | ~x3 | x4) & (x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))))) & (~x3 | ~x7 | (x4 ? (~x5 ^ ~x6) : (x5 | ~x6)));
  assign n4776 = n2061 & ((x3 & ~x4 & (x6 ^ x7)) | (x4 & (x3 ? (~x6 & ~x7) : (x6 & x7))));
  assign n4777 = ~x7 & n543 & (n747 | (~x3 & ~n2982));
  assign n4778 = ~x0 & (n4780 | n4782 | (~x1 & ~n4779));
  assign n4779 = (x2 | x3 | x4 | ~x5 | ~x6) & (~x3 | ((~x5 | x6 | x2 | ~x4) & (~x2 | (x4 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n4780 = ~n2085 & ~n4781;
  assign n4781 = (x2 | ~x4 | ~x5 | x6) & (x5 | ~x6 | ~x2 | x4);
  assign n4782 = n1317 & (x2 ? (x5 & ~n1408) : (~x5 & ~n1353));
  assign n4783 = ~n4784 & (n1898 | n4787) & (n1097 | n4786);
  assign n4784 = x0 & (x1 ? (n704 & n1044) : ~n4785);
  assign n4785 = (~x5 | (x2 ? ((~x4 | x6) & (~x3 | x4 | ~x6)) : (x4 | x6))) & (x2 | ~x4 | ~x6 | (x3 & x5));
  assign n4786 = (x3 | ((x0 | x1 | ~x2 | ~x4) & (~x0 | (x1 ? (x2 | ~x4) : (~x2 | x4))))) & (x0 | ~x3 | ((x2 | x4) & (~x1 | ~x2 | ~x4)));
  assign n4787 = (x0 | (x1 ? (~x2 | x5) : (x2 | ~x5))) & (~x2 | ~x5 | ~x0 | x1);
  assign z240 = ~n4797 | (x6 ? ~n4793 : ~n4789);
  assign n4789 = x1 ? n4791 : (~n2492 & (~x0 | ~n4790));
  assign n4790 = ~x3 & ((~x5 & ~x7 & x2 & ~x4) | (~x2 & x4 & (x5 ^ x7)));
  assign n4791 = (x2 | ~n4792) & (x0 | (~n3468 & (~x2 | ~n4413)));
  assign n4792 = ~x4 & ((~x0 & ((~x5 & ~x7) | (~x3 & x5 & x7))) | (~x5 & ((~x3 & ~x7) | (x0 & x3 & x7))));
  assign n4793 = (x7 | n4794) & (x4 | ~x7 | n4796);
  assign n4794 = (x2 | x3 | n3394) & (x4 | (n4795 & (~x3 | n3394)));
  assign n4795 = (x0 | x1 | ~x3 | ~x5) & (x3 | ((x0 | (x1 ? (~x2 | ~x5) : x5)) & (x5 | ((~x0 | ~x1 | x2) & (x1 | ~x2)))));
  assign n4796 = (x0 | ~x1 | x3 | (~x2 ^ x5)) & (x1 | x5 | (x2 ? ~x3 : ~x0));
  assign n4797 = (n3319 | n4798) & (n640 | n4799);
  assign n4798 = (~x0 | x2 | (x1 ? (x3 | ~x5) : x5)) & (x1 | ((~x2 | x3 | ~x5) & (~x3 | x5))) & (x0 | (x1 ? ((~x3 | ~x5) & (~x2 | x3 | x5)) : (x3 | ~x5)));
  assign n4799 = n4801 & (x4 ? (~n622 | ~n2849) : n4800);
  assign n4800 = (~x0 | x1 | x2 | x3 | ~x5) & (x0 | ((x1 | x2 | ~x3 | x5) & (x3 | ~x5 | ~x1 | ~x2)));
  assign n4801 = (x1 | ~x3 | ~x5) & (x0 | ~x4 | (x1 ? (~x3 ^ x5) : (x3 | x5)));
  assign z241 = n4811 | (~x5 & ~n4803) | (~n640 & ~n4809);
  assign n4803 = ~n4804 & n4806 & (n1408 | (n823 & n1766));
  assign n4804 = n626 & ~n4805;
  assign n4805 = (~x2 | x3 | x4 | ~x6 | x7) & (x2 | ((~x4 | x6 | ~x7) & (~x3 | x4 | ~x6 | x7)));
  assign n4806 = (n4807 | ~n4808) & (~n774 | ~n569 | ~n837);
  assign n4807 = x2 ? (~x4 | x6) : (x4 | ~x6);
  assign n4808 = ~x3 & ~x0 & ~x1;
  assign n4809 = ~n4810 & (~n1121 | (~n880 & (n710 | n2726)));
  assign n4810 = ~n2227 & ((~x1 & x4 & x5) | (~x0 & ((x4 & x5) | (~x1 & ~x4 & ~x5))));
  assign n4811 = ~n2732 & n2332 & ~n643;
  assign z242 = ~n4814 | (~x7 & n626 & ~n4813);
  assign n4813 = (~x2 | x3 | x4 | x5 | x6) & (x2 | (x5 ? ~x6 : (x6 | (~x3 & ~x4))));
  assign n4814 = ~n2507 & (n1008 | n2881) & (~n626 | ~n2477);
  assign z243 = n4816 | ~n4820 | (x6 & ~n4819);
  assign n4816 = n4817 & ((~n4818 & n4808) | (n1322 & n837));
  assign n4817 = ~x4 & ~x7;
  assign n4818 = x2 ? (~x5 ^ ~x6) : (~x5 | x6);
  assign n4819 = x0 ? (x1 & (x2 | x3)) : (~x1 & ~x7 & (~x2 | ~x3));
  assign n4820 = (~n816 | ~n3352) & (~x4 | ~n2753 | ~n4808);
  assign z244 = ~n4825 | n4824 | n4822 | n4823;
  assign n4822 = n939 & ((n757 & n632) | (~x1 & ~n3820));
  assign n4823 = n1084 & ((n951 & n1234) | (n653 & ~n4655));
  assign n4824 = x7 & ((x0 & (~x1 | (~x2 & ~x3))) | (~x1 & x2 & x3) | (~x0 & x1 & (x2 | x3)));
  assign n4825 = ~n4826 & (~n539 | (x1 & ~n572) | (~x1 & n3309));
  assign n4826 = ~x7 & x3 & ~x2 & ~x0 & ~x1;
  assign z245 = n4836 | ~n4834 | n4832 | n4828 | n4829;
  assign n4828 = x0 & (x1 ? (~x2 & ~x3) : x2);
  assign n4829 = ~x2 & ((n939 & n4831) | (n898 & ~n4830));
  assign n4830 = (x1 | x3 | ~x4 | ~x5 | x6) & (~x1 | ~x3 | x4 | x5 | ~x6);
  assign n4831 = x7 & (x1 ? (x5 & x6) : (~x5 & ~x6));
  assign n4832 = ~x0 & ~n4833;
  assign n4833 = (~x1 | ~x2 | ~x3 | ~x4 | ~x5) & (x1 | x3 | x4 | (x2 ^ ~x5));
  assign n4834 = ~n4835 & (~n902 | ~n626) & (~n560 | ~n1268);
  assign n4835 = ~x1 & ~x2 & ~x3 & (x0 ^ x4);
  assign n4836 = n1632 & ((n1005 & n922) | (n626 & n971));
  assign z246 = n4838 | ~n4841 | (x1 & ~n4840);
  assign n4838 = x6 & ((n1287 & n746) | (n772 & ~n4839));
  assign n4839 = (~x3 | ~x5 | x0 | ~x2) & (~x0 | (x2 ? (~x3 | x5) : (x3 | ~x5)));
  assign n4840 = (x2 & (x0 | (~x3 & ~x4 & ~x5))) | (x3 & x4 & x5) | (~x2 & (x3 | (~x0 & x4)));
  assign n4841 = n4842 & (x2 | (~n941 & (~n817 | ~n1244)));
  assign n4842 = (~n837 | ~n1203) & (x1 | n4843);
  assign n4843 = (x0 | ((x2 | ~x4 | ~x5) & (~x2 | x3 | x4 | x5))) & (~x3 | (x2 & (~x0 | ~x4 | ~x5)));
  assign z247 = n4849 | ~n4852 | (x7 & (n4845 | n4847));
  assign n4845 = ~x0 & ((n559 & n1498) | (~x4 & ~n4846));
  assign n4846 = (x1 | ~x2 | ~x3 | x5 | x6) & (x2 | ((x5 | x6 | x1 | x3) & (~x1 | ~x5 | (~x3 ^ x6))));
  assign n4847 = x0 & ((n576 & n577) | (~x1 & ~n4848));
  assign n4848 = (~x2 | x3 | ~x4 | ~x5 | x6) & (x2 | x5 | (x3 ? (x4 | ~x6) : (~x4 | x6)));
  assign n4849 = ~x1 & (x4 ? ~n4850 : ~n4851);
  assign n4850 = (x2 & ((x0 & (x5 ^ x6)) | (~x3 & ~x6) | (x3 & x5 & x6))) | (~x3 & ((~x2 & x5) | (~x0 & x6) | (x0 & ~x6)));
  assign n4851 = (x3 & ((~x2 & ~x5) | (~x0 & (~x2 | (~x5 & ~x6))))) | (~x2 & ~x5 & ~x6) | (~x3 & (x0 | (x2 & x5)));
  assign n4852 = ~n4855 & (~x1 | (n4854 & (x4 | n4853)));
  assign n4853 = (~x3 | x5 | x6 | ~x0 | x2) & (x0 | ((x2 | ~x3 | ~x5 | ~x6) & (~x2 | x3 | x5 | x6)));
  assign n4854 = (x0 | ~x2 | ~x3 | x4) & (~x4 | (x0 ? (x2 | x3) : (~x3 | (x2 & x5))));
  assign n4855 = n1080 & (x0 ? ~n4830 : (n689 & n592));
  assign z248 = n4871 | n4868 | n4857 | ~n4861;
  assign n4857 = x1 & (n4858 | (n902 & n4817 & ~n4860));
  assign n4858 = ~x3 & ((n951 & n3176) | (x5 & ~n4859));
  assign n4859 = (x0 | ~x2 | ~x4 | ~x6 | x7) & (x2 | (x0 ? (x4 ? (x6 | ~x7) : (~x6 | x7)) : (~x7 | (~x4 ^ ~x6))));
  assign n4860 = x0 ? (x5 | ~x6) : (~x5 | x6);
  assign n4861 = n4864 & (~x0 | (~n4862 & (x1 | n4863)));
  assign n4862 = n696 & n979;
  assign n4863 = (x3 | x4 | ~x6 | (x2 & ~x5)) & (~x2 | ~x3 | ~x4 | x5 | x6);
  assign n4864 = (~x1 | n4867) & (x1 | n4865) & (n1353 | n4866);
  assign n4865 = (~x5 | (x0 ? (~x3 | (~x2 ^ x4)) : (x3 | (~x2 ^ ~x4)))) & (~x2 | x5 | (x0 ? (x3 | ~x4) : (~x3 ^ ~x4)));
  assign n4866 = (x0 | ~x1 | ~x2 | x3 | x5) & (x2 | ((x0 | x1 | ~x3 | ~x5) & (~x0 | ((x3 | ~x5) & (x1 | ~x3 | x5)))));
  assign n4867 = (~x0 | x2 | x3 | x4 | x5) & (x0 | ~x3 | (x2 ? (~x4 | x5) : (~x4 ^ ~x5)));
  assign n4868 = ~x0 & ((~n615 & ~n4869) | (x5 & ~n4870));
  assign n4869 = x1 ? (~x2 | ~x5) : (x2 | x5);
  assign n4870 = (~x1 | x2 | x3 | x4 | ~x6) & (x1 | ~x3 | (x2 ? (~x4 | x6) : (x4 | ~x6)));
  assign n4871 = ~x1 & (n4872 | (n1723 & ~n3309 & ~n1433));
  assign n4872 = ~x6 & ((~n697 & ~n2628) | (n743 & n4873));
  assign n4873 = x4 & ~x5 & (~x3 ^ x7);
  assign z249 = n4875 | n4882 | ~n4888 | (x2 & ~n4878);
  assign n4875 = ~x0 & (x2 ? ~n4877 : ~n4876);
  assign n4876 = (~x1 | ((x3 | ~x4 | ~x5 | x6) & (~x3 | x5 | ~x6))) & (x5 | ~x6 | x3 | x4) & (x1 | ((x3 | ~x4 | x5 | x6) & (~x5 | (~x3 ^ (x4 & x6)))));
  assign n4877 = ((~x4 ^ x6) | (x1 ? (x3 | ~x5) : (~x3 ^ ~x5))) & (x1 | x3 | ~x4 | ~x5 | ~x6) & (~x1 | x4 | x5 | (~x3 ^ ~x6));
  assign n4878 = ~n4879 & (~n543 | (~n3589 & (n835 | ~n3795)));
  assign n4879 = ~x1 & (x4 ? (~n835 & ~n4880) : ~n4881);
  assign n4880 = x0 ? (~x5 | x6) : (x5 | ~x6);
  assign n4881 = (x0 | ~x3 | ~x5 | x6 | ~x7) & (x5 | (x3 ^ ~x7) | (x0 ^ x6));
  assign n4882 = ~x2 & (n4883 | (~x0 & (n4885 | ~n4886)));
  assign n4883 = x0 & (x7 ? ~n4438 : ~n4884);
  assign n4884 = (x3 | ~x5 | ((~x4 | x6) & (~x1 | x4 | ~x6))) & (x5 | ((x1 | ~x4 | x6) & (~x3 | x4 | ~x6)));
  assign n4885 = ~n1090 & ((n1392 & n569) | (x3 & ~n3098));
  assign n4886 = (~n1288 | ~n951) & (~n828 | n4887);
  assign n4887 = x5 ? ((~x6 | ~x7) & (~x1 | x6 | x7)) : (x6 | ~x7);
  assign n4888 = ~n4889 & (n1100 | (~n664 & ~n1101));
  assign n4889 = x0 & (x1 ? (n902 & n696) : ~n4890);
  assign n4890 = (x2 | x4 | (~x5 ^ ~x6)) & (~x3 | ((~x5 | ~x6) & (~x2 | x5 | x6)));
  assign z250 = n4898 | n4902 | ~n4904 | (~x2 & ~n4892);
  assign n4892 = ~n4896 & (n2063 | n4650) & (x3 | n4893);
  assign n4893 = (~x5 | n4895) & (~n1769 | ~n4894 | ~x0 | x5);
  assign n4894 = x1 & x4;
  assign n4895 = (x0 | x1 | ~x4 | ~x6 | ~x7) & (x7 | ((x0 | ~x1 | x4 | ~x6) & (~x0 | x6 | (~x1 ^ ~x4))));
  assign n4896 = ~n3394 & (n4897 | (n1029 & n1857));
  assign n4897 = x7 & x6 & ~x3 & ~x4;
  assign n4898 = ~x0 & ((n551 & ~n1171) | n4899 | ~n4901);
  assign n4899 = ~x1 & ((n943 & n859) | (~x2 & n4900));
  assign n4900 = ~x4 & x6 & (x5 ^ x7);
  assign n4901 = ~x1 | x2 | (x4 ? ~n1723 : ~n813);
  assign n4902 = x0 & (x6 ? ~n4903 : (n570 & n886));
  assign n4903 = (~x1 | x2 | x4 | x5 | x7) & (x1 | ((x2 | ~x4 | ~x5 | ~x7) & (~x2 | x4 | x5 | x7)));
  assign n4904 = n4908 & (x6 ? (x7 ? n4905 : n4906) : (x7 ? n4906 : n4905));
  assign n4905 = (x0 | ~x1 | ((x4 | ~x5) & (~x2 | ~x4 | x5))) & (x1 | ((x4 | x5 | x0 | ~x2) & (~x0 | ~x4 | (~x2 & x5))));
  assign n4906 = (~x0 | ~n1084 | n4494) & (~n566 | (n4494 & n4907));
  assign n4907 = (~x3 | ~x5 | ~x1 | x2) & (x1 | x3 | x5);
  assign n4908 = (n4910 | n4911) & (n3319 | (n2485 & n4909));
  assign n4909 = (~x0 | x1 | x2 | x3 | x5) & (x0 | ~x1 | ~x2 | ~x3 | ~x5);
  assign n4910 = (~x4 | ~x6 | ~x0 | x3) & (x4 | x6 | x0 | ~x3);
  assign n4911 = (x1 | ~x2 | ~x5 | x7) & (x5 | ~x7 | ~x1 | x2);
  assign z251 = n4913 | n4916 | ~n4920 | (~n765 & ~n4919);
  assign n4913 = x7 & ((n746 & n1203) | (~x2 & ~n4914));
  assign n4914 = (~n873 | (~n1477 & ~n728)) & (~x0 | n4915);
  assign n4915 = (~x1 | ~x3 | x4 | x5 | x6) & (x1 | ~x5 | (x3 ? (x4 | x6) : (~x4 | ~x6)));
  assign n4916 = ~x7 & ((x6 & ~n4917) | (n3074 & ~n4918));
  assign n4917 = (~n560 | ~n1311) & (n1134 | (~n1644 & ~n3791));
  assign n4918 = (x1 | ~x2 | x3 | ~x4 | ~x5) & (x2 | ((x1 | x3 | ~x4 | x5) & (~x1 | ~x3 | (~x4 ^ x5))));
  assign n4919 = (x6 | ((x2 | x3 | ~x0 | x1) & (~x2 | ~x3 | x0 | ~x1))) & (x1 | ((x0 | ~x3 | ~x6) & ((~x2 ^ x3) | (x0 & ~x6))));
  assign n4920 = ~n4921 & ~n4924 & n4926 & (x3 | n4923);
  assign n4921 = ~x2 & ((n543 & n1741) | (~x1 & ~n4922));
  assign n4922 = (x0 | x3 | ~x5 | x6 | ~x7) & (~x0 | ((~x6 | ~x7 | x3 | x5) & (x6 | x7 | ~x3 | ~x5)));
  assign n4923 = (~x0 | ~x1 | x2 | ~x5 | ~x6) & (x0 | x5 | (x1 ? (~x2 | x6) : (x2 | ~x6)));
  assign n4924 = ~n1008 & ((x2 & ~n800) | (n632 & ~n4925));
  assign n4925 = x0 ? (x3 | x6) : (~x3 | ~x6);
  assign n4926 = ~n570 | (x0 ? (~n1300 | ~n1301) : ~n624);
  assign z252 = n4928 | ~n4933 | ~n4937 | (~n877 & ~n4932);
  assign n4928 = ~x1 & (n4930 | (x4 & n743 & n4929));
  assign n4929 = ~x6 & x7 & (x3 ^ ~x5);
  assign n4930 = x2 & ((n564 & n4929) | (~x7 & ~n4931));
  assign n4931 = (x0 | x3 | ~x4 | x5 | ~x6) & (x6 | ((~x4 | ~x5 | x0 | ~x3) & (~x0 | x4 | (~x3 ^ ~x5))));
  assign n4932 = (~x0 | x1 | x2 | x6 | x7) & (x0 | ((x1 | ~x2 | ~x6 | ~x7) & (~x1 | (x2 ? (x6 | x7) : (~x6 | ~x7)))));
  assign n4933 = ~n4935 & (~n543 | (n4934 & (~n885 | ~n1725)));
  assign n4934 = x2 ? (~x7 | (x3 ? (~x4 | x6) : ~x6)) : (x7 | (x3 ? (~x4 ^ x6) : (~x4 ^ ~x6)));
  assign n4935 = ~n643 & (~n4936 | (n1716 & n837));
  assign n4936 = (x2 | x3 | x0 | x1) & (~x0 | ((x1 | ~x2 | ~x3 | ~x4) & (~x1 | x2 | x3)));
  assign n4937 = (n1566 | n4932) & (x1 | (n4939 & (n1566 | n4938)));
  assign n4938 = (x0 | ~x2 | ~x4 | x6 | x7) & (~x0 | ((x2 | ~x4 | ~x6 | ~x7) & (~x2 | x4 | x6)));
  assign n4939 = n4941 & (x4 | n4940);
  assign n4940 = x0 ? (x2 | ~x7 | (~x3 ^ ~x6)) : (~x2 | x7 | (~x3 ^ x6));
  assign n4941 = (~x0 | ~x2 | x3 | ~x4 | x6) & (x0 | x2 | ~x3 | ~x6);
  assign z253 = ~n4943 | n4946 | ~n4948 | (n743 & ~n4947);
  assign n4943 = n4944 & (~n2940 | ~n3812) & (x2 | n4945);
  assign n4944 = (x0 | x1 | ~x3 | (~x2 ^ x7)) & (x3 | ((x0 | ~x1 | ~x2 | x7) & (~x0 | (x1 ? (x2 | x7) : (~x2 | ~x7)))));
  assign n4945 = (~n830 | ~n1244) & (~x5 | n627 | n2223);
  assign n4946 = n543 & ((~x4 & ~x7 & ~x2 & ~x3) | (x4 & (x2 ? (x3 & x7) : (x3 ^ x7))));
  assign n4947 = (~x1 | ~x3 | x4 | x5 | x7) & (x1 | ~x4 | (x3 ? (~x5 ^ ~x7) : (x5 | ~x7)));
  assign n4948 = (x1 | n4949) & (x0 | n4950);
  assign n4949 = (x3 | ((x4 | ~x7 | ~x0 | x2) & (x0 | (x2 ? (x4 | ~x7) : (~x4 | x7))))) & (~x0 | ~x3 | (x2 ? (~x4 ^ x7) : (x4 | x7)));
  assign n4950 = (x4 | n4951) & (x3 | ~x4 | ~n570 | n1008);
  assign n4951 = (x1 | x2 | x3 | ~x5 | x7) & (~x1 | ~x3 | ~x7 | (~x2 ^ ~x5));
  assign z255 = ~n4960 | (x1 ? ~n4953 : (n4956 | n4958));
  assign n4953 = ~n609 & ~n4954;
  assign n4954 = ~x0 & ((n530 & n949) | (x4 & ~n4955));
  assign n4955 = (x2 | ~x3 | ~x5 | x6 | x7) & (x5 | ((x2 | x3 | x6 | ~x7) & (~x2 | x7 | (~x3 ^ x6))));
  assign n4956 = x2 & ((~x6 & ~n4957) | (x0 & n2836));
  assign n4957 = (~x0 | ~x3 | x4 | x5 | x7) & (x0 | ((x3 | x4 | ~x5 | x7) & (x5 | ~x7 | ~x3 | ~x4)));
  assign n4958 = ~x2 & ((x4 & ~n4959) | (~x0 & ~x4 & n1293));
  assign n4959 = (x0 | x3 | x5 | x6 | x7) & (~x0 | ~x5 | ~x7 | (~x3 ^ x6));
  assign n4960 = n1305 & ~n4961 & (~n1875 | n4963);
  assign n4961 = ~x0 & (x5 ? (~n1353 & n3555) : ~n4962);
  assign n4962 = (~x1 | x2 | x3 | ~x4 | ~x6) & (~x2 | (x1 ? (x3 ? (x4 | ~x6) : (~x4 | x6)) : (~x3 | (~x4 ^ ~x6))));
  assign n4963 = (~x1 | x2 | x3 | x4 | ~x6) & (x1 | ((~x2 | ~x3 | ~x4 | x6) & (x2 | ((x4 | x6) & (~x3 | ~x4 | ~x6)))));
  assign z256 = ~n4974 | n4971 | n4969 | n1319 | n4965;
  assign n4965 = ~x2 & ((x1 & ~n4966) | n4967 | (~x1 & ~n4968));
  assign n4966 = (~x0 | x3 | ~x4 | ~x5 | ~x6) & (x0 | x5 | ((x4 | x6) & (x3 | ~x4 | ~x6)));
  assign n4967 = ~n1097 & (~n1327 | (n774 & n841));
  assign n4968 = (~x4 | ((~x0 | (x3 ? (~x5 | ~x6) : (x5 | x6))) & (x0 | x3 | x5 | ~x6))) & (x0 | x4 | (x3 ? x5 : (~x5 | x6)));
  assign n4969 = ~n765 & ((n3575 & n1269) | (~x2 & ~n4970));
  assign n4970 = (x0 | ~x1 | ~x3 | x4 | ~x6) & (~x0 | ~x4 | x6 | (x1 ^ ~x3));
  assign n4971 = ~n4973 & (x2 ? n4817 : n4972);
  assign n4972 = x4 & x7;
  assign n4973 = (~x0 | x1 | x3 | ~x5 | ~x6) & (x0 | ~x1 | x6 | (~x3 ^ ~x5));
  assign n4974 = x0 ? (x1 | n4980) : (~n4975 & ~n4978);
  assign n4975 = x4 & ((n804 & n4976) | (x2 & ~n4977));
  assign n4976 = ~x3 & ~x6 & (x5 ^ x7);
  assign n4977 = (x5 | ~x7 | ((~x3 | x6) & (~x1 | x3 | ~x6))) & (x1 | ~x5 | x7 | (~x3 ^ x6));
  assign n4978 = ~n4979 & x6 & n1084;
  assign n4979 = (x5 | x7 | ~x1 | x3) & (x1 | ~x7 | (~x3 ^ ~x5));
  assign n4980 = (x4 | n4982) & (~x6 | ~n4981 | ~x2 | ~x4);
  assign n4981 = x7 & (x3 ^ ~x5);
  assign n4982 = (x2 | x5 | ~x6 | x7) & (~x2 | ~x3 | x6 | (~x5 ^ x7));
  assign z257 = ~n4994 | (x5 ? (n4990 | n4993) : ~n4984);
  assign n4984 = x7 ? n4985 : (n4989 & (x1 | n4988));
  assign n4985 = x3 ? n4986 : n4987;
  assign n4986 = (x0 | ~x1 | ~x2 | ~x4 | x6) & (~x0 | x1 | x2 | x4 | ~x6);
  assign n4987 = (x0 | ~x1 | x6 | (~x2 ^ x4)) & (~x6 | ((x0 | ((x2 | x4) & (~x1 | ~x2 | ~x4))) & (x1 | ((x2 | x4) & (~x0 | ~x2 | ~x4)))));
  assign n4988 = (x0 | ((x2 | ~x3 | ~x4 | x6) & (~x2 | x3 | x4 | ~x6))) & (~x4 | ~x6 | x2 | x3) & (~x0 | ((~x2 | (x3 ? (x4 | ~x6) : (~x4 | x6))) & (x2 | ~x3 | x4 | x6)));
  assign n4989 = (~n733 | ~n2352) & (n1353 | n1766);
  assign n4990 = ~x1 & ((~n640 & ~n4991) | (x6 & ~n4992));
  assign n4991 = (x0 | x2 | ~x3 | x4) & (~x2 | (x0 ? (~x3 ^ ~x4) : (x3 | ~x4)));
  assign n4992 = (x0 | ~x2 | ~x3 | x4 | x7) & (~x0 | x2 | x3 | ~x4 | ~x7);
  assign n4993 = n543 & ((n1044 & n1786) | (~n643 & n1619));
  assign n4994 = n5003 & ~n5000 & ~n4995 & ~n4997;
  assign n4995 = ~x6 & ((n731 & n746) | (~x3 & ~n4996));
  assign n4996 = (x0 | ~x1 | x2 | (~x4 ^ ~x5)) & (~x2 | ((x4 | x5 | ~x0 | x1) & (x0 | (x1 ? (x4 | ~x5) : (~x4 | x5)))));
  assign n4997 = ~x2 & ((x3 & ~n4998) | (n1051 & ~n4999));
  assign n4998 = x0 ? (x1 | ~x4 | (~x6 ^ x7)) : (~x1 | x4 | (~x6 ^ ~x7));
  assign n4999 = (~x0 | (x1 ? (~x4 | ~x7) : (x4 | x7))) & (x0 | x1 | ~x4 | ~x7);
  assign n5000 = x6 & ((~x2 & ~n5001) | (n742 & ~n5002));
  assign n5001 = x0 ? (x4 | (x1 ? (x3 | x5) : ~x5)) : (~x3 | ~x4 | (x1 & x5));
  assign n5002 = (~x3 | x4 | x5) & (~x4 | ~x5 | ~x1 | x3);
  assign n5003 = (n981 | n1350) & (~n3431 | n5004);
  assign n5004 = (x0 | ~x1 | x3 | ~x4 | x7) & (x1 | ~x7 | (x0 ? (~x3 | x4) : (~x3 ^ ~x4)));
  assign z258 = n5011 | ~n5014 | (x3 ? ~n5009 : ~n5006);
  assign n5006 = (~x2 | x6 | ~n841 | n1337) & (x2 | n5007);
  assign n5007 = (x0 | ~x1 | x5 | ~n3251) & (x1 | n5008);
  assign n5008 = x0 ? (~x6 | (x4 ? (x5 | ~x7) : (~x5 | x7))) : (x5 | x6 | (x4 ^ ~x7));
  assign n5009 = (x1 | n3381) & (n765 | n5010);
  assign n5010 = (~x0 | x1 | x2 | ~x4 | x6) & (x0 | x4 | (x1 ? (x2 | x6) : (~x2 | ~x6)));
  assign n5011 = ~n643 & (x3 ? ~n5013 : ~n5012);
  assign n5012 = (x0 | x1 | ~x5 | (~x2 ^ x4)) & (~x1 | (~x4 ^ ~x5) | (x0 ^ ~x2));
  assign n5013 = (~x0 | x1 | ~x2 | x4 | ~x5) & (x0 | ~x4 | x5 | (~x1 ^ ~x2));
  assign n5014 = ~n5016 & ~n5018 & n5020 & (n765 | n5015);
  assign n5015 = ((~x3 ^ ~x4) | (x0 ? (x1 | ~x2) : (~x1 | x2))) & (~x0 | x1 | x2 | x3 | ~x4) & (x0 | ((~x1 | ~x2 | ~x3 | x4) & (x1 | (x2 ? (x3 | ~x4) : (~x3 | x4)))));
  assign n5016 = ~x2 & ((~n1605 & n5017) | (n674 & n727));
  assign n5017 = ~x5 & x0 & ~x4;
  assign n5018 = n742 & (n5019 | (n674 & n927));
  assign n5019 = x7 & ~x5 & ~x4 & ~x1 & ~x3;
  assign n5020 = (n1036 | n4754) & (n1337 | (~n829 & ~n3416));
  assign z259 = ~n5026 | n5030 | (x3 ? ~n5022 : ~n5032);
  assign n5022 = ~n5025 & (x0 ? (~n632 | ~n588) : n5023);
  assign n5023 = (x5 | x6 | ~n1145 | n3309) & (~x5 | (~n5024 & (~x6 | ~n1145 | n3309)));
  assign n5024 = x4 & ((~x7 & (x1 ? (x2 ^ x6) : (~x2 & ~x6))) | (~x1 & x2 & ~x6 & x7));
  assign n5025 = ~n697 & ((n704 & n841) | (~n1097 & ~n1580));
  assign n5026 = x5 ? (n5028 & (~x6 | n5027)) : (x6 | n5027);
  assign n5027 = (~x0 | x3 | (x1 ? (x2 | ~x4) : x4)) & (~x2 | ((x0 | ~x4 | (~x1 ^ x3)) & (x1 | x4 | (~x0 & x3))));
  assign n5028 = (x1 | n5029) & (~n3488 | (~n1044 & ~n1619));
  assign n5029 = (~x4 | ~x6 | x2 | x3) & (x6 | ((~x4 | ((~x2 | x3) & (~x0 | (~x2 & x3)))) & (x2 | x4 | (x0 & ~x3))));
  assign n5030 = ~x5 & ((n745 & n733) | (x6 & ~n5031));
  assign n5031 = (~x3 | ((x1 | x2 | ~x4) & (x0 | (x1 ? (~x2 ^ ~x4) : (~x2 | x4))))) & (~x1 | x3 | x4 | (x0 ^ ~x2));
  assign n5032 = ~n5035 & (x0 | (~n5034 & (~x1 | n5033)));
  assign n5033 = x2 ? (x7 | (x4 ? (x5 | ~x6) : (~x5 | x6))) : (~x6 | ~x7 | (x4 & x5));
  assign n5034 = n1467 & ((n1518 & n569) | (~n697 & ~n1408));
  assign n5035 = n5036 & (x1 ? (~x2 & ~x7) : x7);
  assign n5036 = x0 & (x4 ? (~x5 & x6) : (x5 & ~x6));
  assign z260 = n5038 | n5044 | n5049 | (~n3319 & ~n5048);
  assign n5038 = ~x2 & (n5039 | n5042 | (n1188 & ~n5043));
  assign n5039 = ~x3 & ((~x4 & ~n5040) | (n772 & ~n5041));
  assign n5040 = (~x0 | ~x1 | x5 | x6 | x7) & (~x6 | ((x1 | ~x5 | x7) & (x0 | ((~x5 | x7) & (x1 | x5 | ~x7)))));
  assign n5041 = (~x0 & x5) | (x0 & x6) | (~x5 & ~x7);
  assign n5042 = ~n4758 & ((n569 & n689) | (x1 & ~n3315));
  assign n5043 = x0 ? ((x4 | ~x5 | ~x6 | x7) & (~x4 | x5 | x6 | ~x7)) : (x5 ? (x6 | ~x7) : (x7 | (~x4 ^ x6)));
  assign n5044 = ~n640 & ((~x1 & ~n5045) | ~n5047 | (x1 & ~n5046));
  assign n5045 = (x0 | ~x5 | (~x3 ^ x4)) & (x5 | (x0 ? ((~x3 | x4) & (~x2 | x3 | ~x4)) : (~x2 | (~x3 ^ ~x4))));
  assign n5046 = (x0 | ~x2 | ~x3 | x4 | ~x5) & (~x0 | x2 | x3 | ~x4 | x5);
  assign n5047 = x0 ? (x1 | ((~x3 | ~x5) & (x2 | x3 | x5))) : (~x1 | ((x3 | x5) & (x2 | ~x3 | ~x5)));
  assign n5048 = x3 ? ((x1 | x5) & (x0 | (x5 & (x1 | ~x2)))) : (~x5 | (~x0 ^ (x1 & x2)));
  assign n5049 = x2 & ((n1986 & ~n5050) | n5051 | ~n5052);
  assign n5050 = (~x1 | x3 | ~x4 | ~x5 | x6) & (x1 | ~x6 | (x3 ? (x4 | x5) : ~x5));
  assign n5051 = ~n877 & ((n550 & n841) | (~x0 & n548));
  assign n5052 = (~n550 | ~n699) & (~n548 | ~n712);
  assign z261 = ~n5062 | (x2 ? (n5059 | n5061) : ~n5054);
  assign n5054 = x0 ? (~n5056 & (~x3 | n5055)) : n5057;
  assign n5055 = (~x1 | x4 | x5 | ~x6 | x7) & (x1 | ((x4 | ~x5 | ~x6 | x7) & (~x4 | x6 | ~x7)));
  assign n5056 = n526 & n689 & (x4 | ~x6);
  assign n5057 = x1 ? n5058 : (~n828 | ~n951);
  assign n5058 = (x3 | ((x5 | x6 | ~x7) & (x4 | ~x5 | x7))) & (~x5 | ((~x4 | ~x6 | x7) & (x6 | ~x7 | ~x3 | x4)));
  assign n5059 = ~x0 & (x1 ? (n1029 & n978) : ~n5060);
  assign n5060 = (x5 | (x4 ? (~x6 | x7) : (x6 | ~x7))) & (~x3 | ~x5 | (x4 ? (x6 | ~x7) : (~x6 | x7)));
  assign n5061 = n841 & (x5 ? (n828 & n569) : ~n1850);
  assign n5062 = ~n5066 & ~n5069 & ~n5071 & (n643 | n5063);
  assign n5063 = (x4 | n5065) & (~x4 | ~x5 | ~n626 | n5064);
  assign n5064 = x2 & x3;
  assign n5065 = (~x0 | x1 | (x2 ? (~x3 | ~x5) : (x3 | x5))) & (~x1 | ((x3 | ~x5 | ~x0 | x2) & (x0 | x5 | (~x2 & ~x3))));
  assign n5066 = ~n640 & (~n5068 | (~x2 & ~n5067));
  assign n5067 = (x3 | ((~x1 | (x0 ? (~x4 | ~x5) : (x4 | x5))) & (~x0 | x1 | (~x4 ^ x5)))) & (~x0 | x1 | ~x3 | (~x4 ^ ~x5));
  assign n5068 = (x0 | (x1 ? (~x4 | (x2 & x5)) : (x4 | ~x5))) & (x1 | ~x2 | ((x4 | x5) & (~x0 | ~x4 | ~x5)));
  assign n5069 = x1 & ((n728 & n2435) | (~x3 & ~n5070));
  assign n5070 = x0 ? (x2 | x5 | (~x4 ^ x6)) : (~x2 | ~x5 | (~x4 ^ ~x6));
  assign n5071 = n626 & n934 & (n2352 | n5072);
  assign n5072 = x3 & (x4 ^ ~x6);
  assign z262 = ~n5079 | ~n5086 | (~x0 & (n5074 | n5077));
  assign n5074 = ~x3 & ((~x4 & ~n5075) | (n4972 & ~n5076));
  assign n5075 = (~x7 | (~x5 ^ ~x6) | (~x1 ^ x2)) & (~x6 | x7 | (x1 ? (~x2 | x5) : (x2 | ~x5)));
  assign n5076 = (x5 | x6 | ~x1 | x2) & (x1 | ~x2 | (~x5 ^ ~x6));
  assign n5077 = x7 & n1188 & (n5078 | (n1364 & n1518));
  assign n5078 = x2 & (x5 ^ ~x6);
  assign n5079 = ~n5082 & ~n5084 & (x2 ? n5080 : n5081);
  assign n5080 = (~x0 | x1 | ~x3 | x5 | ~x7) & (x0 | ((~x1 | (x3 ? (x5 | x7) : (~x5 | ~x7))) & (x1 | x3 | ~x5 | x7)));
  assign n5081 = ((~x1 ^ ~x7) | (x0 ? (x3 | x5) : (~x3 | ~x5))) & (~x0 | ~x1 | x3 | ~x5 | x7) & (x0 | x1 | x5 | ~x7);
  assign n5082 = ~x1 & ((n674 & n547) | (n2061 & ~n5083));
  assign n5083 = (~x4 | ~x7 | ~x2 | x3) & (x4 | x7 | x2 | ~x3);
  assign n5084 = n543 & ((n1044 & n717) | (x2 & ~n5085));
  assign n5085 = (~x5 | ~x7 | ~x3 | x4) & (x5 | x7 | x3 | ~x4);
  assign n5086 = (~x0 | n5089) & (n1198 | (~n5088 & (x0 | n5087)));
  assign n5087 = (x1 | ~x2 | ~x3 | x7) & (~x1 | ((x2 | x7) & (~x4 | ~x7 | ~x2 | ~x3)));
  assign n5088 = x7 & n841 & (~x2 | n828);
  assign n5089 = (~n845 | ~n979) & (x1 | x7 | n5090);
  assign n5090 = (~x5 & x6) | (x5 & ~x6) | (~x2 & (~x3 | (~x4 & ~x6)));
  assign z263 = ~n5104 | ~n5092 | n5100;
  assign n5092 = ~n5094 & ~n5096 & n5098 & (x2 | n5093);
  assign n5093 = x0 ? ((x1 | ~x3 | ~x4 | x6) & (~x1 | x3 | ~x6)) : ((~x1 | x3 | x4 | x6) & (x1 | ~x6 | (~x3 ^ x4)));
  assign n5094 = x3 & ((n845 & n1269) | (n898 & ~n5095));
  assign n5095 = (x1 | ~x2 | ~x4 | ~x5 | x6) & (~x1 | x2 | x4 | x5 | ~x6);
  assign n5096 = ~n643 & (~n5097 | (~n4758 & n3555));
  assign n5097 = (x2 | x3 | ~x0 | x1) & (x0 | ~x2 | (x1 ? (~x3 | ~x4) : x3));
  assign n5098 = (~n829 | ~n3687) & (~n873 | n5099);
  assign n5099 = (~x5 | ~x6 | ~x2 | x4) & (x5 | x6 | x2 | ~x4);
  assign n5100 = ~n640 & (n5102 | ~n5103 | (n841 & n5101));
  assign n5101 = x2 & (~x3 ^ ~x4);
  assign n5102 = n653 & ((n2332 & n804) | (x1 & ~n1122));
  assign n5103 = x0 ? (~n570 | ~n1641) : ~n979;
  assign n5104 = (~x2 | n5105) & (~n1188 | n5106);
  assign n5105 = (~x0 | x1 | x3 | x4 | x6) & (x0 | ((x1 | ~x3 | ~x4 | x6) & (~x1 | ~x6 | (~x3 ^ x4))));
  assign n5106 = (x0 | x2 | ~x4 | x5 | ~x6) & (~x5 | ((~x0 | (x2 ? (~x4 | ~x6) : (x4 | x6))) & (x0 | ~x2 | x4 | x6)));
  assign z264 = ~n5111 | (x6 & (n5109 | (n873 & ~n5108)));
  assign n5108 = (x2 | ~x4 | ~x5 | x7) & (x5 | ~x7 | ~x2 | x4);
  assign n5109 = ~x1 & ((n2705 & n1250) | (x2 & ~n5110));
  assign n5110 = (x0 | ~x3 | x4 | x5 | ~x7) & (~x0 | ~x4 | (x3 ? (~x5 | ~x7) : (x5 | x7)));
  assign n5111 = ~n5120 & ~n5119 & ~n5117 & ~n5112 & n5114;
  assign n5112 = x4 & ((n733 & n1460) | (~x1 & ~n5113));
  assign n5113 = (x0 | x2 | ~x3 | x5 | ~x7) & (x7 | ((x0 | x2 | ~x3 | ~x5) & (~x0 | ~x2 | (~x3 ^ x5))));
  assign n5114 = n5116 & (~x2 | n5115);
  assign n5115 = (x0 | ~x3 | ~x7 | (~x1 ^ x4)) & ((x0 ? (x1 | x4) : (~x1 | ~x4)) | (~x3 ^ x7));
  assign n5116 = (x0 | x1 | ~x2 | x3 | x7) & (x2 | ((x0 | ~x1 | ~x3 | x7) & (~x0 | x3 | (~x1 ^ ~x7))));
  assign n5117 = n1005 & ((n1269 & n2209) | (x0 & ~n5118));
  assign n5118 = (x1 | ~x2 | ~x4 | ~x5 | x7) & (~x1 | x2 | x4 | x5 | ~x7);
  assign n5119 = n572 & ((~x3 & ~x4 & ~x0 & x1) | (~x1 & (x0 ? (x3 & x4) : (x3 ^ x4))));
  assign n5120 = ~x4 & ((~n765 & ~n3676) | (n626 & n5121));
  assign n5121 = x5 & (x2 ? (x3 & x7) : (~x3 & ~x7));
  assign z265 = ~n5132 | n5130 | ~n5123 | n5127;
  assign n5123 = n5126 & (x2 ? (x1 | ~n5125) : n5124);
  assign n5124 = (x3 | ((x0 | ~x1 | ~x4 | x5) & (~x0 | ~x5 | (~x1 ^ ~x4)))) & (x1 | ~x3 | (x0 ? (x4 | x5) : (~x4 ^ x5)));
  assign n5125 = x3 & (x0 ? (x4 ^ x5) : (x4 & x5));
  assign n5126 = ((x0 ? (x1 | x3) : (~x1 | ~x3)) | (~x2 ^ x4)) & (x0 | x3 | (x1 ? (x2 | x4) : (~x2 | ~x4)));
  assign n5127 = ~x2 & ((n830 & n1234) | (~x3 & ~n5128));
  assign n5128 = (n5129 | n3553) & (x0 | ~n1145 | ~n951);
  assign n5129 = x1 ? (~x4 | x6) : (x4 | ~x6);
  assign n5130 = n596 & (x0 ? (n772 & n813) : ~n5131);
  assign n5131 = (x1 | x4 | ~x5 | ~x6 | ~x7) & (~x1 | ((x4 | x5 | ~x6 | x7) & (x6 | ~x7 | ~x4 | ~x5)));
  assign n5132 = x2 ? (~n5136 & (~n1358 | ~n712)) : n5133;
  assign n5133 = (x5 | n5135) & (x1 | ~x5 | n5134);
  assign n5134 = (x4 | x6 | x0 | x3) & (~x4 | ~x6 | ~x0 | ~x3);
  assign n5135 = (~x0 | ~x1 | (x3 ? (x4 | x6) : (~x4 | ~x6))) & (x0 | x1 | x4 | ~x6);
  assign n5136 = ~x0 & ((n696 & n1188) | (x1 & n5137));
  assign n5137 = ~x3 & (x4 ? (x5 & x6) : (~x5 & ~x6));
  assign z266 = ~n5140 | n5143 | ~n5147 | (n1468 & ~n5139);
  assign n5139 = (~x4 | x5 | x6 | ~x0 | x1) & (x0 | ((~x5 | ~x6 | x1 | x4) & (~x1 | (x4 ? (~x5 | x6) : (x5 | ~x6)))));
  assign n5140 = (~x1 | n5141) & (~x0 | x1 | n5142);
  assign n5141 = (~x5 | ~x6 | x0 | ~x3) & (x3 | ((~x5 | ~x6 | ~x0 | x2) & (x0 | x5 | (x2 ^ ~x6))));
  assign n5142 = (~x3 | ~x4 | ~x5 | x6) & (x2 | ((~x3 | x4 | x5 | x6) & (x3 | ~x4 | ~x6)));
  assign n5143 = ~x2 & (n5145 | n5146 | (~n5144 & ~n3587));
  assign n5144 = x1 ? (x3 | x7) : (~x3 | ~x7);
  assign n5145 = ~x7 & ((n653 & n1207) | (n704 & n1234));
  assign n5146 = ~n1040 & ((n841 & n683) | (n543 & n2438));
  assign n5147 = ~n5148 & (n1566 | n5152) & (x1 | n5151);
  assign n5148 = ~x0 & (x4 ? (n1317 & n5149) : ~n5150);
  assign n5149 = ~x5 & (~x2 ^ x6);
  assign n5150 = (x5 | ~x6 | x1 | x3) & (~x1 | ~x5 | x6 | (x2 & ~x3));
  assign n5151 = (x6 | ((x3 | x5 | ~x0 | x2) & (x0 | (~x3 ^ x5)))) & (~x0 | ~x6 | ((~x3 | x5) & (~x2 | x3 | ~x5)));
  assign n5152 = (x0 | x1 | ~x4 | ~x6) & (~x0 | x4 | x6 | (x1 ^ ~x2));
  assign z267 = n5159 | ~n5161 | (x6 ? ~n5157 : ~n5154);
  assign n5154 = ~n5155 & (x2 | (~n5156 & (~n674 | ~n699)));
  assign n5155 = ~n671 & ~n1219;
  assign n5156 = n4089 & ((n626 & n1451) | (x0 & ~n1221));
  assign n5157 = (n1218 | n1215) & (~n3522 | n5158);
  assign n5158 = (x0 | x3 | ~x4 | ~x7) & (x4 | x7 | ~x0 | ~x3);
  assign n5159 = ~x2 & ((n1358 & n1734) | (~x4 & ~n5160));
  assign n5160 = (x6 | ((x3 | x5 | ~x0 | x1) & (x0 | (x1 ? (x3 | ~x5) : (~x3 | x5))))) & (~x0 | ~x6 | (x1 ? x3 : (~x3 | x5)));
  assign n5161 = ~n5164 & (n4226 | ~n5162) & (~n543 | ~n5163);
  assign n5162 = ~x5 & ~x4 & ~x1 & x2;
  assign n5163 = ~x4 & (x5 ^ ~x6);
  assign n5164 = ~x1 & ((x5 & (x0 ? (x4 ^ x6) : (~x4 & ~x6))) | (~x5 & x6 & ~x0 & x4));
  assign z268 = n5171 | (x2 ? ~n5175 : (~n5166 | ~n5176));
  assign n5166 = ~n5167 & (~n689 | n5170);
  assign n5167 = x1 & ((n1070 & n5168) | (~x7 & ~n5169));
  assign n5168 = ~x4 & ~x0 & ~x3;
  assign n5169 = (x4 | x5 | ~x0 | ~x3) & (x0 | x3 | (x4 ? (~x5 ^ x6) : (~x5 ^ ~x6)));
  assign n5170 = (x0 | ~x4 | x5 | x6 | x7) & (~x0 | ~x5 | ~x7 | (~x4 ^ x6));
  assign n5171 = ~x2 & (~n5173 | (x0 & ~n5172));
  assign n5172 = (x5 | x7 | ~x1 | x3) & (x1 | x6 | (x3 ? (x5 | x7) : (~x5 ^ x7)));
  assign n5173 = (~n813 | ~n727) & (n1198 | n5174);
  assign n5174 = (x0 | ~x1 | ~x3 | x7) & (~x0 | ~x7 | (x1 ^ ~x3));
  assign n5175 = (x1 | ((~x0 | (x5 ? (x6 | ~x7) : x7)) & (~x6 | x7 | x0 | ~x5) & (x5 | (~x6 ^ ~x7)))) & (x0 | ((x5 | x6 | ~x7) & (~x1 | (x5 ? (~x6 ^ ~x7) : (~x6 | x7)))));
  assign n5176 = (~x0 | x1 | x5 | ~x6 | x7) & (x0 | ((x1 | (x5 ? (~x6 | x7) : ~x7)) & (~x7 | ((x5 | x6) & (~x1 | ~x5 | ~x6)))));
  assign z269 = ~n5180 | n5182 | (~x2 & (~n5178 | ~n5183));
  assign n5178 = (~n601 | ~n699) & (x7 | ~n2061 | n5179);
  assign n5179 = (x1 | x3 | ~x4 | ~x6) & (x4 | x6 | ~x1 | ~x3);
  assign n5180 = (x2 | x3 | n5181) & (~n2320 | (~x2 & x7));
  assign n5181 = (~x0 | x1 | x4 | ~x6 | x7) & (x0 | ~x1 | ~x7 | (~x4 ^ ~x6));
  assign n5182 = ~x1 & (x0 ? ((x6 & x7) | (x2 & ~x6 & ~x7)) : (x6 ^ x7));
  assign n5183 = (~x0 | ~x1 | x3 | (~x6 ^ ~x7)) & (~x3 | ((x0 | ~x1 | ~x6 | ~x7) & (x6 | x7 | ~x0 | x1)));
  assign z270 = n5185 | n5187 | ~n5188 | (~x2 & ~n5174);
  assign n5185 = n878 & ((n699 & n867) | (x0 & ~n5186));
  assign n5186 = (x1 | x3 | ~x4 | ~x5 | x7) & (~x1 | ~x3 | x4 | x5 | ~x7);
  assign n5187 = n1044 & ((n2296 & n543) | (n841 & n2316));
  assign n5188 = n5189 & (x7 | ~n1044 | n586);
  assign n5189 = (x1 | ~x2 | ~x7) & (x0 | (x1 ? (~x2 | x7) : ~x7));
  assign z271 = ~n5193 | (~x3 & ~n5191) | (n1080 & ~n5192);
  assign n5191 = (~x0 | x1 | x2 | ~x4 | x5) & (x0 | ((x1 | ~x2 | x4 | ~x5) & (~x1 | (x2 ? (~x4 | ~x5) : (x4 | x5)))));
  assign n5192 = (~n577 | ~n699) & (~x0 | n4830);
  assign n5193 = n5197 & (x1 ? n5195 : (x3 | n5194));
  assign n5194 = x0 ? (x2 | x4) : (~x2 | ~x4);
  assign n5195 = (~n696 | ~n594) & (~n653 | n5196);
  assign n5196 = (x2 | x4 | ~x5 | x6) & (~x2 | ~x4 | x5 | ~x6);
  assign n5197 = ~n2435 & ~n4457 & (~n3687 | ~n5198);
  assign n5198 = ~x3 & x2 & ~x0 & ~x1;
  assign z272 = n5208 | ~n5200 | n5205;
  assign n5200 = ~n5201 & (~n742 | ~n2438 | n5204);
  assign n5201 = ~x2 & (x0 ? ~n5202 : ~n5203);
  assign n5202 = (~x1 | ((x3 | ~x5) & (~x3 | x4 | x5 | x6))) & (x3 | (x5 ? x4 : (~x4 & ~x6))) & (x1 | ((x3 | x5) & (~x5 | ~x6 | ~x3 | ~x4)));
  assign n5203 = x3 ? (~x4 & (x1 | (~x5 & ~x6))) : (~x1 | x4 | (x5 & x6));
  assign n5204 = (x1 | x4 | ~x5 | x6) & (~x1 | ~x4 | x5 | ~x6);
  assign n5205 = x2 & (~n5207 | (~x0 & ~n5206));
  assign n5206 = (~x4 | x5 | x6 | ~x1 | x3) & (x1 | x4 | (x3 ? (~x5 | ~x6) : (x5 | x6)));
  assign n5207 = (x1 | (x0 ? x3 : (~x3 | ~x4))) & (x0 | ((~x3 | ~x4 | ~x5) & (~x1 | x3 | x4)));
  assign n5208 = ~x7 & (n3096 | (~x2 & ~n5192));
  assign z273 = n5217 | ~n5220 | (~x5 & (~n5210 | ~n5215));
  assign n5210 = x1 ? (~n5211 & (~n1783 | ~n1395)) : n5213;
  assign n5211 = x6 & (x0 ? (~x2 & ~n1381) : (x2 & n5212));
  assign n5212 = x3 & (~x4 ^ ~x7);
  assign n5213 = (~n548 | ~n549) & (~n653 | n5214);
  assign n5214 = (~x2 | x4 | ~x6 | x7) & (x2 | ~x4 | x6 | ~x7);
  assign n5215 = x3 ? n5216 : (~n626 | n1977);
  assign n5216 = (x0 | x1 | x2 | ~x4 | ~x6) & (x6 | ((x2 | x4 | ~x0 | ~x1) & (x0 | (x1 ? (~x2 | ~x4) : (x2 | x4)))));
  assign n5217 = x5 & ((~x2 & ~n5218) | (n3818 & ~n5219));
  assign n5218 = x6 ? (n1218 | ~n873) : (~n841 | n3972);
  assign n5219 = (~x6 | ~x7 | ~x0 | x3) & (x6 | x7 | x0 | ~x3);
  assign n5220 = ~n5227 & ~n5225 & n5221 & n5222;
  assign n5221 = (x0 | x1 | x2 | ~x4 | ~x5) & ((~x2 ^ ~x5) | (x0 ? (x1 | ~x4) : (~x1 | x4)));
  assign n5222 = (~n5223 | n5194) & (n5224 | (~n2857 & ~n2094));
  assign n5223 = x5 & ~x1 & ~x3;
  assign n5224 = x1 ? (x2 | ~x5) : (~x2 | x5);
  assign n5225 = ~n1408 & (n5226 | (x2 & n543 & n1451));
  assign n5226 = x5 & x3 & ~x2 & x0 & ~x1;
  assign n5227 = ~n791 & ((n570 & n3021) | (n632 & n3575));
  assign z274 = n5229 | ~n5234 | ~n5237 | (~n1548 & ~n5233);
  assign n5229 = ~x2 & (n5230 | n5231);
  assign n5230 = ~n1008 & ((n841 & n598) | (n543 & n2352));
  assign n5231 = x6 & ((n1234 & n2209) | (~x0 & ~n5232));
  assign n5232 = (x1 | ~x3 | ~x4 | ~x5 | ~x7) & (~x1 | x4 | (x3 ? (x5 | ~x7) : (~x5 | x7)));
  assign n5233 = x0 ? ((~x1 | x2 | x5 | x6) & (x1 | (x2 ? ~x5 : (x5 | ~x6)))) : ((~x1 | x2 | ~x5 | x6) & (x1 | ~x2 | x5 | ~x6));
  assign n5234 = (n1097 | n5235) & (n604 | n5236);
  assign n5235 = (~x0 | ~x1 | x2 | x3 | x4) & (x0 | ((x1 | x2 | ~x3 | x4) & (x3 | ~x4 | ~x1 | ~x2)));
  assign n5236 = (x0 | ~x1 | x2 | ~x5) & (x1 | (x0 ? (~x2 ^ ~x5) : (~x2 | x5)));
  assign n5237 = ~n5238 & ~n5242 & ~n5245 & (~n742 | n5241);
  assign n5238 = ~x2 & ((~n823 & ~n5239) | (~x0 & ~n5240));
  assign n5239 = (x3 | x4 | x5 | ~x6) & (~x3 | ~x4 | ~x5 | x6);
  assign n5240 = (~x3 | ((~x5 | ~x6 | ~x1 | x4) & (x5 | x6 | x1 | ~x4))) & (x1 | x3 | ~x5 | (x4 & ~x6));
  assign n5241 = x1 ? ((~x5 | ~x6 | x3 | x4) & (~x3 | x5 | x6)) : (~x4 | x6 | (~x3 ^ ~x5));
  assign n5242 = ~n765 & ((n543 & n5244) | (x4 & ~n5243));
  assign n5243 = (~x0 | ((x1 | ~x2 | ~x3 | x6) & (~x1 | x2 | x3 | ~x6))) & (x0 | x1 | x2 | x3 | x6);
  assign n5244 = x2 & ~x4 & (x3 ^ ~x6);
  assign n5245 = x2 & ((n866 & n931) | (n1145 & ~n5246));
  assign n5246 = (x0 | x3 | x5 | ~x6 | x7) & ((~x5 ^ x7) | (x0 ? (x3 | ~x6) : (~x3 | x6)));
  assign z275 = n5266 | n5263 | ~n5253 | n5248 | n5250;
  assign n5248 = ~n640 & ((n746 & n1311) | (~x5 & ~n5249));
  assign n5249 = (x0 | ~x1 | ~x2 | x3 | x4) & (x1 | ~x3 | (x0 ? (~x2 ^ ~x4) : (~x2 | x4)));
  assign n5250 = ~x0 & (x1 ? ~n5252 : ~n5251);
  assign n5251 = (x2 | ~x3 | ~x4 | x5 | x6) & (~x2 | x3 | x4 | ~x5 | ~x6);
  assign n5252 = (x2 | x3 | x4 | x5 | x6) & (~x3 | ~x6 | (x2 ? (~x4 | ~x5) : (~x4 ^ x5)));
  assign n5253 = n5262 & ~n5261 & ~n5259 & ~n5254 & ~n5256;
  assign n5254 = ~x6 & ~n5255;
  assign n5255 = (x0 | ~x2 | ~x4 | (~x1 ^ x3)) & (x2 | ((x0 | x1 | ~x3 | x4) & (~x0 | (x1 ? (x3 | x4) : (~x3 | ~x4)))));
  assign n5256 = ~x1 & ((n1044 & n5257) | (x5 & ~n5258));
  assign n5257 = x4 & ~x5 & (x6 ^ ~x7);
  assign n5258 = (x2 | x3 | ~x4 | x6 | x7) & (~x2 | ~x3 | x4 | ~x6 | ~x7);
  assign n5259 = n5260 & (n2537 | (n681 & n1044));
  assign n5260 = x6 & x0 & ~x1;
  assign n5261 = ~n1119 & ((n1156 & n813) | (n530 & n1518));
  assign n5262 = (~n576 | ~n2402) & (~x6 | n1685 | ~n4808);
  assign n5263 = ~n643 & (x0 ? ~n5265 : ~n5264);
  assign n5264 = x1 ? ((~x3 | ((x4 | x5) & (~x2 | (x4 & x5)))) & (x2 | x3 | (~x4 & ~x5))) : ((x2 | ~x3 | ~x4 | ~x5) & (~x2 | x3 | x4 | x5));
  assign n5265 = x1 ? (x2 | (x3 ? (x4 | x5) : ~x4)) : (~x2 | x3 | (x4 & x5));
  assign n5266 = ~x1 & (n5270 | (x5 & (n5267 | n5268)));
  assign n5267 = ~x0 & ((n885 & n1786) | (n1044 & n1668));
  assign n5268 = x0 & ((n885 & n3790) | (n1084 & ~n5269));
  assign n5269 = x3 ? (x6 | x7) : (~x6 | ~x7);
  assign n5270 = n3434 & n817;
  assign z276 = n5278 | ~n5280 | (x1 ? ~n5272 : ~n5274);
  assign n5272 = x0 ? (~n1044 | ~n931) : (~n5273 & (~n1044 | ~n1950));
  assign n5273 = ~n643 & ((~x4 & ~x5 & x2 & x3) | (~x2 & x4 & (x3 ^ ~x5)));
  assign n5274 = ~n5277 & (n1218 | n5275) & (x6 | n5276);
  assign n5275 = (x0 | x2 | ~x3 | x5 | x6) & (~x2 | ((~x0 | ~x6 | (~x3 ^ ~x5)) & (x0 | x3 | ~x5 | x6)));
  assign n5276 = (~x3 | ~n670 | x0 | ~x2) & (x2 | x3 | ~n867);
  assign n5277 = ~n835 & n743 & x6 & n2332;
  assign n5278 = ~n671 & ~n5279;
  assign n5279 = (~x0 | ((x1 | ~x2 | ~x3 | x5) & (~x1 | x2 | x3 | ~x5))) & (x1 | x2 | ((x3 | x5) & (x0 | ~x3 | ~x5)));
  assign n5280 = n5289 & ~n5287 & ~n5285 & ~n5281 & ~n5284;
  assign n5281 = ~x0 & (x2 ? ~n5282 : ~n5283);
  assign n5282 = x1 ? (~x5 | ((~x4 | ~x7) & (~x3 | x4 | x7))) : (x5 | ((x4 | x7) & (x3 | ~x4 | ~x7)));
  assign n5283 = (x1 | ~x3 | x4 | x5 | ~x7) & (x7 | ((x3 | ~x4 | ~x5) & (~x1 | (x3 ? (x4 | x5) : ~x5))));
  assign n5284 = n1188 & (x0 ? (~x2 & ~n1218) : (x2 & n4972));
  assign n5285 = ~n1205 & ~n5286;
  assign n5286 = x0 ? ((x1 | ~x2 | ~x4 | ~x5) & (~x1 | x2 | x4 | x5)) : (~x2 | (x1 ? (~x4 | x5) : (x4 | ~x5)));
  assign n5287 = ~n714 & ~n5288;
  assign n5288 = (~x2 | x3 | x7 | ~x0 | x1) & (x0 | ~x1 | x2 | ~x3 | ~x7);
  assign n5289 = (~n2765 | ~n746) & (~n560 | ~n5290);
  assign n5290 = ~x7 & x5 & ~x3 & x4;
  assign z277 = ~n5303 | ~n5299 | n5292 | n5296;
  assign n5292 = ~x0 & (n5293 | (n619 & ~n5295));
  assign n5293 = x1 & ((n1070 & n1556) | (~x7 & ~n5294));
  assign n5294 = x2 ? ((~x3 | x4 | ~x5 | ~x6) & (x3 | (x4 ? (~x5 | x6) : (x5 | ~x6)))) : ((x3 | ~x5 | ~x6) & (x5 | x6 | ~x3 | ~x4));
  assign n5295 = ((x3 ? (~x4 | x5) : (x4 | ~x5)) | (~x2 ^ x6)) & (~x2 | x3 | ~x4 | ~x5 | ~x6) & (x5 | x6 | x2 | x4);
  assign n5296 = x0 & ((n576 & n1626) | (~x1 & ~n5297));
  assign n5297 = (n1353 | n5298) & (~x7 | n615 | ~n691);
  assign n5298 = (~x2 | ~x7 | (~x3 ^ ~x5)) & (x5 | x7 | x2 | x3);
  assign n5299 = ~n5301 & (x4 | n1356) & (n1198 | n5300);
  assign n5300 = x1 ? ((x2 | x3 | ~x4) & (~x3 | x4 | x0 | ~x2)) : ((x3 | x4 | ~x0 | ~x2) & (x0 | ~x3 | (~x2 ^ ~x4)));
  assign n5301 = x2 & ((~n2259 & n5302) | (n696 & n699));
  assign n5302 = ~x1 & (~x0 ^ x3);
  assign n5303 = ~n5305 & (~x4 | n5304);
  assign n5304 = (x0 | ~x1 | ~x2 | (~x3 ^ ~x5)) & (x1 | (x0 ? (x2 ? (x3 | ~x5) : (~x3 | x5)) : (x2 | (~x3 ^ ~x5))));
  assign n5305 = ~x2 & (x5 ? ~n5306 : (n841 & n598));
  assign n5306 = (~x0 | x1 | x3 | ~x6) & (x0 | ~x1 | (x3 ? (~x4 | ~x6) : (x4 | x6)));
  assign z278 = ~n5324 | ~n5316 | n5313 | n5308 | n5311;
  assign n5308 = ~x3 & ((~x1 & ~n5309) | (n543 & ~n5310));
  assign n5309 = (x0 | x4 | (x2 ? (~x5 ^ ~x6) : (x5 | ~x6))) & (~x4 | ((x0 | ~x2 | x5 | ~x6) & (~x0 | ~x5 | (x2 & x6))));
  assign n5310 = x4 ? (x2 ? (~x5 ^ ~x6) : (x5 | ~x6)) : (~x5 | x6);
  assign n5311 = x3 & ((~x0 & ~n1278) | (n841 & ~n5312));
  assign n5312 = (x2 | x4 | x5 | ~x6) & (~x2 | (x4 ? (x5 | ~x6) : (~x5 ^ ~x6)));
  assign n5313 = ~n671 & ((n804 & ~n5315) | (x2 & ~n5314));
  assign n5314 = (x0 | x1 | x3 | ~x5 | x6) & ((~x3 ^ ~x5) | (x0 ? (x1 | x6) : (~x1 | ~x6)));
  assign n5315 = x0 ? (x3 ? (~x5 | ~x6) : (x5 | x6)) : (x3 ? (x5 | x6) : (~x5 | ~x6));
  assign n5316 = n5319 & ~n5321 & ~n5323 & (n5317 | n5318);
  assign n5317 = (x3 | x5) & (~x2 | ~x3 | ~x5);
  assign n5318 = (x0 | ~x1 | x4 | x6 | x7) & (~x0 | x1 | ~x4 | ~x6 | ~x7);
  assign n5319 = (n2128 | n2953) & (~n3818 | n5320);
  assign n5320 = x0 ? (x3 | ~x6) : (~x3 | x6);
  assign n5321 = ~n682 & ~n5322;
  assign n5322 = (x3 | x4 | ~x0 | x2) & (x0 | ~x3 | (~x2 ^ ~x4));
  assign n5323 = n1518 & (x0 ? (x1 ? (~x3 & x6) : (x3 & ~x6)) : (x1 ? (x3 & x6) : (~x3 & ~x6)));
  assign n5324 = ~n5327 & (x4 | (~n5325 & (~n1283 | ~n1403)));
  assign n5325 = ~x7 & ((n3269 & n837) | (~x1 & n5326));
  assign n5326 = (x2 ? (~x5 & x6) : (x5 & ~x6)) & (~x0 ^ x3);
  assign n5327 = n566 & ((n576 & n658) | (x7 & ~n5328));
  assign n5328 = (x1 | x2 | ~x3 | x5 | ~x6) & (x3 | ~x5 | (x1 ? (x2 ^ ~x6) : (~x2 | ~x6)));
  assign z279 = ~n5344 | ~n5339 | ~n5337 | n5330 | n5334;
  assign n5330 = x1 & (n4374 | n5331);
  assign n5331 = ~x0 & (x3 ? ~n5332 : ~n5333);
  assign n5332 = x2 ? ((~x6 | ~x7 | ~x4 | ~x5) & (x6 | x7 | x4 | x5)) : (x4 ? (x5 ? (~x6 | x7) : (x6 | ~x7)) : (x7 | (~x5 ^ x6)));
  assign n5333 = (x2 | x4 | x5 | x6 | ~x7) & (~x6 | ((x2 | ~x4 | x5 | x7) & (~x2 | (x4 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n5334 = ~x1 & (x2 ? ~n5335 : ~n5336);
  assign n5335 = x0 ? ((~x5 | ~x7 | ~x3 | ~x4) & (x3 | (x4 ? (x5 | ~x7) : (~x5 | x7)))) : ((x3 | ~x4 | ~x5 | ~x7) & (~x3 | x4 | x5 | x7));
  assign n5336 = (x0 | ~x3 | x4 | ~x5 | x7) & (x5 | ((x0 | ~x3 | ~x4 | ~x7) & (~x0 | (x3 ? (x4 | x7) : (~x4 | ~x7)))));
  assign n5337 = (n643 | n5338) & (~x3 | n1040 | ~n2940);
  assign n5338 = x3 ? (~n570 | n1679) : (n1164 | n2267);
  assign n5339 = ~n5340 & (n1353 | n5342) & (x3 | n5343);
  assign n5340 = ~n2803 & ~n5341;
  assign n5341 = x1 ? (x2 | (x0 ? (x3 | ~x5) : (~x3 ^ ~x5))) : ((~x3 | ~x5 | x0 | ~x2) & ((~x2 ^ x5) | (x0 ^ x3)));
  assign n5342 = x0 ? ((x1 | ~x2 | ~x3 | x5) & (~x1 | x2 | x3 | ~x5)) : (x1 | ~x2 | (~x3 ^ ~x5));
  assign n5343 = (~x2 | ~n926 | x0 | ~x1) & (~x0 | x1 | x2 | ~n2720);
  assign n5344 = x1 ? n5345 : (~n5347 & (x2 | n5348));
  assign n5345 = x0 ? (~n1044 | ~n2209) : n5346;
  assign n5346 = (~x2 | ~x3 | (x4 ? (x5 | x7) : (~x5 | ~x7))) & (x3 | ((x5 | ~x7 | ~x2 | x4) & (x2 | ~x5 | (~x4 ^ ~x7))));
  assign n5347 = ~n2466 & ~n1113;
  assign n5348 = (n2129 | n5349) & (x7 | ~n828 | n4880);
  assign n5349 = (x4 | ~x5 | x6 | ~x7) & (~x4 | ~x6 | (~x5 ^ ~x7));
  assign z280 = n5351 | ~n5356 | ~n5364 | (~x0 & ~n5354);
  assign n5351 = ~n640 & ((~x1 & ~n5352) | (n2074 & ~n5353));
  assign n5352 = (x0 | ~x2 | ~x3 | x4 | ~x5) & (~x4 | ((x0 | x2 | ~x3 | ~x5) & (~x0 | (x2 ? (x3 | ~x5) : (~x3 | x5)))));
  assign n5353 = (x3 | x4 | ~x0 | x2) & (x0 | ~x2 | (~x3 ^ ~x4));
  assign n5354 = ~n5355 & (~n1017 | (~n2409 & (x3 | ~n881)));
  assign n5355 = ~x1 & (x2 ? n2202 : (n1392 & n813));
  assign n5356 = ~n5357 & ~n5360 & ~n5362 & (n1389 | n5361);
  assign n5357 = x3 & ((~x0 & ~n5358) | (n841 & ~n5359));
  assign n5358 = (~x1 | x4 | ~x5 | (~x2 ^ ~x6)) & (~x4 | x5 | (x1 ? (~x2 | ~x6) : (x2 ^ ~x6)));
  assign n5359 = (x2 | x4 | x5 | ~x6) & (~x5 | (x2 ? (~x4 ^ ~x6) : (~x4 | x6)));
  assign n5360 = n793 & ((n4894 & n658) | (~x1 & ~n2055));
  assign n5361 = (x6 | x7 | ~x2 | x5) & (~x6 | ~x7 | x2 | ~x5);
  assign n5362 = ~n2063 & (n5363 | (x3 & n1181 & ~n1164));
  assign n5363 = ~x4 & ~x3 & x2 & x0 & ~x1;
  assign n5364 = ~n5367 & (n643 | (~x2 & n5365) | (x2 & n5366));
  assign n5365 = x0 ? ((x4 | x5 | ~x1 | ~x3) & (x3 | ((~x4 | ~x5) & (x1 | (~x4 & ~x5))))) : (x1 ? (x3 ? ~x4 : (x4 | x5)) : (~x3 | x4));
  assign n5366 = (x0 | ~x1 | ~x3 | x4 | x5) & (x1 | (x0 ? (x3 ? (~x4 | x5) : x4) : (~x4 | (~x3 ^ ~x5))));
  assign n5367 = ~x3 & ((~x5 & ~n5368) | (n1380 & ~n5369));
  assign n5368 = (~x0 | x2 | x6 | (~x1 ^ ~x4)) & (~x6 | (x0 ? (x1 ? (x2 | x4) : (~x2 | ~x4)) : (x1 ? (~x2 ^ x4) : (x2 | x4))));
  assign n5369 = (~x1 | ~x2 | ~x4 | x6) & (x1 | (x2 ? (~x4 ^ ~x6) : (~x4 | x6)));
  assign z281 = n5380 | ~n5382 | (x1 ? ~n5371 : ~n5375);
  assign n5371 = ~n5374 & (x0 | (x2 & n5372) | (~x2 & n5373));
  assign n5372 = (x3 | ~x4 | x5 | ~x6 | ~x7) & (x6 | (x3 ? (x4 ? (x5 | ~x7) : (~x5 | x7)) : (~x4 | (~x5 ^ ~x7))));
  assign n5373 = (x3 | x4 | ~x5 | x6 | ~x7) & (~x6 | ((x4 | x5 | ~x7) & (~x3 | ~x4 | (~x5 ^ ~x7))));
  assign n5374 = n600 & n845;
  assign n5375 = x3 ? n5378 : n5376;
  assign n5376 = x6 ? n5377 : (~n742 | (~n674 & ~n2705));
  assign n5377 = x2 ? (x4 | (x0 ? (~x5 ^ ~x7) : (x5 | ~x7))) : (~x4 | ((x5 | ~x7) & (~x0 | ~x5 | x7)));
  assign n5378 = (~n658 | ~n3996) & (x4 | n5379);
  assign n5379 = (x0 | x2 | x5 | ~x6 | x7) & ((x0 ? (~x2 | x5) : (x2 | ~x5)) | (~x6 ^ ~x7));
  assign n5380 = ~n643 & ((n1716 & n1269) | (x5 & ~n5381));
  assign n5381 = (x0 | x1 | ~x2 | ~x3 | ~x4) & (x2 | (x1 ? (x3 | ~x4) : (x4 | (~x0 & x3))));
  assign n5382 = ~n5383 & n5385 & ~n5387 & (~n1181 | n5390);
  assign n5383 = ~n671 & ~n5384;
  assign n5384 = (x0 | ~x1 | ~x3 | ~x5) & (x1 | x2 | x5 | (~x0 & x3));
  assign n5385 = (n1337 | (~n587 & ~n1101)) & (n2129 | n5386);
  assign n5386 = (~x1 | x2 | x4 | x5 | x7) & (x1 | ~x4 | ((~x5 | ~x7) & (~x2 | x5 | x7)));
  assign n5387 = x2 & (x5 ? ~n5389 : (~n1205 & n5388));
  assign n5388 = ~x4 & ~x0 & x1;
  assign n5389 = (x0 | ~x1 | x3 | x4 | x7) & (~x0 | x1 | (x3 ? (x4 | ~x7) : (~x4 | x7)));
  assign n5390 = (x1 | ~x3 | ~x4 | ~x5 | x7) & (x5 | ((x1 | ~x3 | ~x4 | ~x7) & (~x1 | (x3 ? (x4 | x7) : (~x4 | ~x7)))));
  assign z282 = ~n5396 | ~n5402 | ~n5406 | (~x1 & ~n5392);
  assign n5392 = n5394 & (x5 | (~n5393 & (~n2435 | ~n1585)));
  assign n5393 = n1051 & ((n1181 & n4089) | (x0 & ~n3770));
  assign n5394 = (n1977 | ~n4365) & (n1408 | n5395);
  assign n5395 = (~x3 | x5 | x7 | ~x0 | x2) & (x0 | ~x2 | x3 | ~x5 | ~x7);
  assign n5396 = ~n5398 & n5400 & (n1097 | n5397);
  assign n5397 = x2 ? ((x1 | ~x3 | ~x4) & (x0 | (x1 ? (~x3 | x4) : ~x4))) : ((~x1 | x3 | ~x4) & (~x0 | x1 | x4));
  assign n5398 = ~x1 & ((~n1408 & ~n5399) | (n547 & n577));
  assign n5399 = (x0 | x2 | ~x3 | ~x5) & (x3 | x5 | ~x0 | ~x2);
  assign n5400 = x1 ? (~n1044 | ~n728) : n5401;
  assign n5401 = (x2 | x3 | ~x4 | ~x5 | x6) & (~x2 | ~x3 | x4 | x5 | ~x6);
  assign n5402 = ~n5403 & (n671 | (~n5405 & (~n3436 | n4869)));
  assign n5403 = ~n2227 & ~n5404;
  assign n5404 = (~x0 | x1 | ~x4 | ~x5 | x6) & (x0 | ((~x1 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (x5 | ~x6 | x1 | x4)));
  assign n5405 = n971 & ((n543 & n934) | (x0 & ~n753));
  assign n5406 = ~n5407 & (~x1 | (~n2581 & ~n5410));
  assign n5407 = ~n1218 & ((n543 & ~n5409) | (~x1 & ~n5408));
  assign n5408 = (~x0 | ~x2 | ~x3 | ~x5 | x6) & (x5 | ~x6 | x2 | x3);
  assign n5409 = (~x5 | ~x6 | ~x2 | x3) & (x5 | x6 | x2 | ~x3);
  assign n5410 = ~x0 & ((n1070 & n2003) | (~n1134 & ~n5411));
  assign n5411 = (x6 | x7 | ~x2 | x3) & (~x6 | ~x7 | x2 | ~x3);
  assign z283 = ~n5429 | n5425 | ~n5419 | n5413 | n5416;
  assign n5413 = ~n1008 & (x2 ? ~n5414 : ~n5415);
  assign n5414 = x3 ? (~x6 | ((x1 | ~x4) & (x0 | (x1 & ~x4)))) : (x4 | x6 | (~x0 ^ x1));
  assign n5415 = (~x0 | ~x1 | x3 | x4 | ~x6) & (x0 | ((~x3 | ~x4 | x6) & (x4 | ~x6 | x1 | x3)));
  assign n5416 = ~x2 & (n5417 | n5418 | (n699 & n809));
  assign n5417 = ~x1 & ((n825 & n809) | (x0 & ~n4754));
  assign n5418 = ~n1008 & ((n1392 & n922) | (~x0 & ~n1820));
  assign n5419 = ~n5420 & n5423 & (~n1465 | n5422);
  assign n5420 = ~x2 & (x0 ? (n813 & n1317) : ~n5421);
  assign n5421 = (~x1 | x3 | x5 | x6 | x7) & (~x6 | ~x7 | ~x3 | ~x5);
  assign n5422 = (x2 | x5 | ~x0 | x1) & (x0 | ~x1 | (~x2 ^ ~x5));
  assign n5423 = (~n1365 | ~n3435) & (~x2 | n823 | n5424);
  assign n5424 = (x3 | x5 | ~x6 | x7) & (~x3 | ~x5 | x6 | ~x7);
  assign n5425 = ~x2 & (n5426 | (~x1 & (n5427 | n5428)));
  assign n5426 = x1 & ((n951 & n2204) | (n978 & n1074));
  assign n5427 = x0 & ((~n693 & ~n1097) | (n774 & n813));
  assign n5428 = n1310 & (n1525 | (x3 & ~n3319));
  assign n5429 = ~x2 | (n5430 & ~n5432 & (~n626 | n5434));
  assign n5430 = x0 ? (~n689 | ~n717) : n5431;
  assign n5431 = (~x3 | x4 | x5 | x7) & (x1 | x3 | (x4 ? (x5 | x7) : (~x5 | ~x7)));
  assign n5432 = ~n2803 & (n5433 | (n3151 & n841));
  assign n5433 = ~x5 & x3 & ~x0 & x1;
  assign n5434 = (x3 | x4 | x5 | ~x6 | x7) & (x6 | (x3 ? (x4 ? (x5 | x7) : (~x5 | ~x7)) : (~x5 | (~x4 ^ ~x7))));
  assign z284 = n5436 | ~n5438 | n5444 | (~x6 & ~n5450);
  assign n5436 = ~n640 & ((n731 & n1269) | (~x3 & ~n5437));
  assign n5437 = (x1 & ((x0 & (x2 | (~x4 & ~x5))) | (x2 & ~x4 & ~x5) | (x5 & (x4 | (~x0 & ~x2))))) | (x0 & x2 & ~x4) | (~x1 & ((~x2 & x4) | (~x0 & (x4 | (~x2 & ~x5)))));
  assign n5438 = x3 ? (~n5441 & ~n5443) : (~n5439 & n5440);
  assign n5439 = ~n1998 & ((n1723 & n772) | (x1 & ~n2819));
  assign n5440 = (x0 | ~x1 | x2 | ~n1364) & (x1 | n1559);
  assign n5441 = n5442 & (x0 ? n2359 : n1479);
  assign n5442 = ~x1 & (~x2 | ~x5);
  assign n5443 = n543 & ((n706 & n859) | (~x2 & ~n1040));
  assign n5444 = x6 & (n5445 | ~n5447);
  assign n5445 = ~x0 & ((n674 & n676) | (~x4 & ~n5446));
  assign n5446 = (~x1 | ((~x3 | ~x5 | x7) & (~x2 | x3 | x5 | ~x7))) & (x2 | ~x3 | ~x5 | x7) & (x1 | x5 | ((~x3 | x7) & (x2 | x3 | ~x7)));
  assign n5447 = (x2 | ((~x4 | n5449) & (~x1 | x4 | ~n5448))) & (x1 | ~x4 | ~n5448) & (~x2 | x4 | n5449);
  assign n5448 = ~x7 & ~x5 & x0 & x3;
  assign n5449 = (x0 | ~x1 | ~x3 | x5 | x7) & (~x0 | x1 | ~x5 | (~x3 ^ x7));
  assign n5450 = ~n5453 & (x0 | (~n5451 & (~x7 | n5452)));
  assign n5451 = ~n1090 & ((n885 & n4089) | (~x2 & ~n3972));
  assign n5452 = (~x1 | ~x3 | ~x4 | x5) & (x1 | x4 | ((~x3 | ~x5) & (x2 | x3 | x5)));
  assign n5453 = n1365 & (n4972 | (n1429 & n1084));
  assign z285 = x4 ? (~n5455 | ~n5464) : (~n5459 | ~n5467);
  assign n5455 = ~n5456 & (~n1080 | n5458);
  assign n5456 = x2 & ((~n5269 & ~n3394) | (~x0 & ~n5457));
  assign n5457 = (~x1 | ~x3 | x5 | ~x6 | ~x7) & (x1 | ~x5 | ((~x6 | x7) & (x3 | x6 | ~x7)));
  assign n5458 = (x0 | ~x1 | x3 | ~x5 | x6) & (x1 | ((x5 | x6 | x0 | x3) & (~x0 | ~x6 | (~x3 ^ x5))));
  assign n5459 = x2 ? n5462 : (~n5460 & (x5 | n5461));
  assign n5460 = ~n1090 & ((n569 & n622) | (~x0 & ~n871));
  assign n5461 = (x0 | x1 | x3 | ~x6 | x7) & (~x0 | ~x3 | x6 | (~x1 ^ ~x7));
  assign n5462 = (~x3 | x7 | (x6 ? n3394 : ~n5463)) & (~x7 | (x6 ? ~n5463 : n3394));
  assign n5463 = x5 & ~x0 & ~x1;
  assign n5464 = n5466 & (x1 | n5465);
  assign n5465 = (~x0 | x7 | (x2 ? x3 : (~x3 | ~x5))) & (~x7 | ((x2 | x3 | x5) & (x0 | (x2 & x5))));
  assign n5466 = (~n746 | ~n2575) & (n765 | n3771);
  assign n5467 = n5469 & (~n1986 | n3625) & (x2 | n5468);
  assign n5468 = (~x1 | x5 | (x0 ? (x3 | ~x7) : (~x3 ^ ~x7))) & (~x0 | x1 | (x3 ? ~x7 : (~x5 | x7)));
  assign n5469 = x1 | ~x2 | (x0 ? ~n757 : ~n1453);
  assign z286 = n5474 | ~n5482 | (x4 ? ~n5471 : ~n5477);
  assign n5471 = ~n5472 & (x3 | ~n1723 | ~n742 | n1543);
  assign n5472 = ~x6 & ((n543 & n5121) | (~x1 & ~n5473));
  assign n5473 = (x0 | x2 | x3 | ~x5 | ~x7) & (x7 | ((x3 | x5 | x0 | x2) & (~x0 | ~x3 | (~x2 ^ ~x5))));
  assign n5474 = ~x2 & ((~n2290 & ~n5475) | (x3 & ~n5476));
  assign n5475 = (x0 & x3) | (~x6 & (~x4 | (~x0 & ~x3)));
  assign n5476 = (x4 | x6 | (x0 ? (~x1 | x5) : (x1 | ~x5))) & (~x0 | x1 | ~x5 | (~x4 & ~x6));
  assign n5477 = ~n5478 & ~n5481 & (x3 | ~n1181 | ~n951);
  assign n5478 = ~x7 & ((n3269 & n816) | (n5479 & ~n5480));
  assign n5479 = x0 & x6;
  assign n5480 = (~x1 | x2 | ~x3 | x5) & (x1 | ~x2 | x3 | ~x5);
  assign n5481 = ~n765 & (x0 ? (~x1 & n878) : (x1 & n1146));
  assign n5482 = ~n5485 & (~x2 | (n5484 & (~x5 | n5483)));
  assign n5483 = (x1 | ~x3 | x4 | x6) & (x0 | ~x1 | x3 | ~x4 | ~x6);
  assign n5484 = (x1 | (x3 ? (x5 | ~x6) : (~x5 | x6))) & (x0 | ~x1 | ((x5 | x6) & (~x3 | ~x5 | ~x6)));
  assign n5485 = ~n1008 & ((~n913 & n3436) | (~x3 & ~n5486));
  assign n5486 = (x0 | x1 | ~x2 | x4 | ~x6) & (~x0 | ((x1 | ~x2 | ~x4 | ~x6) & (~x1 | x2 | x4 | x6)));
  assign z287 = n5495 | ~n5498 | (x1 ? ~n5488 : ~n5491);
  assign n5488 = ~n3926 & (x0 | (~x3 & n5490) | (x3 & n5489));
  assign n5489 = (x2 | x4 | ~x5 | ~x6 | x7) & (~x2 | ~x4 | x5 | x6 | ~x7);
  assign n5490 = x2 ? ((~x4 | x5 | ~x6 | x7) & (x4 | ~x5 | x6 | ~x7)) : ((~x4 | x5 | x6 | ~x7) & (x4 | (x5 ? (~x6 | x7) : (~x6 ^ ~x7))));
  assign n5491 = ~n5493 & (~x2 | (~n5492 & (~n2438 | n1082)));
  assign n5492 = ~x3 & ~n1198 & (x0 ? n4089 : n1379);
  assign n5493 = n1080 & ~n5494;
  assign n5494 = x0 ? ((x5 | x6 | ~x3 | ~x4) & (x3 | ~x6 | (~x4 ^ x5))) : (x4 | (x3 ? (~x5 ^ ~x6) : (~x5 | x6)));
  assign n5495 = ~x3 & ((n4464 & ~n5496) | (x2 & ~n5497));
  assign n5496 = x0 ? (~x4 | ~x6) : (x4 | x6);
  assign n5497 = x6 ? (x7 | (x0 ? x1 : x4)) : (~x7 | ((x1 | ~x4) & (x0 | (x1 & ~x4))));
  assign n5498 = n5501 & (n640 | n5499) & (~n1188 | n5500);
  assign n5499 = (~x3 | ~x4 | x0 | ~x2) & (x2 | ((x0 | x3 | ~x4) & (x4 | (~x0 ^ (x1 & x3)))));
  assign n5500 = (~x0 | ~x2 | ~x4 | x6 | x7) & (x0 | x2 | x4 | ~x6 | ~x7);
  assign n5501 = (~n2352 | ~n837) & (~x3 | n710 | n1977);
  assign z288 = ~n5503 | n5507 | n5513 | (~x1 & ~n5511);
  assign n5503 = (~x2 | n5506) & (~n543 | n5504) & (x2 | n5505);
  assign n5504 = (x2 | x3 | x4 | ~x5 | ~x7) & (x7 | (x2 ? (x3 ? (~x4 | ~x5) : (~x4 ^ x5)) : ((x4 | x5) & (x3 | ~x4 | ~x5))));
  assign n5505 = x3 ? ((x0 | ~x4 | ~x7) & (x1 | ((~x4 | ~x7) & (~x0 | x4 | x7)))) : (x0 ? (~x1 | (~x4 ^ ~x7)) : (x1 | (~x4 ^ x7)));
  assign n5506 = (x0 | ~x1 | ~x3 | x4 | ~x7) & (x1 | (x0 ? (x3 ? (x4 | ~x7) : (~x4 | x7)) : (x7 | (~x3 ^ ~x4))));
  assign n5507 = x5 & (n5508 | (~x4 & n825 & ~n5510));
  assign n5508 = ~x3 & (x2 ? ~n5509 : (n841 & n2467));
  assign n5509 = (x0 | ~x1 | ~x4 | (~x6 ^ ~x7)) & (~x0 | x1 | x4 | ~x6 | x7);
  assign n5510 = (x1 | ~x2 | x6 | ~x7) & (~x1 | x2 | (~x6 ^ ~x7));
  assign n5511 = x0 ? n5512 : (~n3032 & (n765 | n2099));
  assign n5512 = x2 ? ((x5 | ~x7 | x3 | x4) & (~x3 | ~x4 | (~x5 ^ x7))) : (x3 | (x4 ? (x5 | ~x7) : (~x5 ^ ~x7)));
  assign n5513 = ~x5 & ((~x6 & ~n5514) | (n1686 & ~n5516));
  assign n5514 = (x2 | n5515) & (~x2 | ~x7 | ~n543 | n1744);
  assign n5515 = (x0 | ~x1 | x3 | ~x4 | ~x7) & (~x0 | ~x3 | (x1 ? (x4 | ~x7) : (~x4 | x7)));
  assign n5516 = (~x1 | x2 | x3 | x4 | ~x7) & (~x2 | ((~x4 | ~x7 | x1 | x3) & (~x1 | x7 | (~x3 ^ ~x4))));
  assign z289 = n5518 | ~n5523 | ~n5529 | (x5 & ~n5522);
  assign n5518 = x6 & (n5519 | (n743 & ~n5521));
  assign n5519 = ~x0 & (x7 ? (n2074 & ~n2075) : ~n5520);
  assign n5520 = (x1 | ~x2 | (x3 ? (x4 | ~x5) : (~x4 | x5))) & (x3 | x5 | ~x1 | x2);
  assign n5521 = (~x1 | ~x3 | x4 | x5 | x7) & (x1 | ~x7 | (x3 ? (~x4 ^ ~x5) : (~x4 | x5)));
  assign n5522 = x2 ? ((x3 | ~x4 | ~x0 | x1) & (x0 | ~x1 | ~x3 | x4)) : ((x4 | (x0 ? (~x1 ^ x3) : (x1 | x3))) & (x0 | ~x1 | ~x3 | ~x4));
  assign n5523 = n5527 & (x3 | (~n5524 & (~n559 | ~n837)));
  assign n5524 = n3074 & (n5526 | (x1 & (~x5 | n5525)));
  assign n5525 = x5 & x2 & x4;
  assign n5526 = ~x5 & x4 & ~x1 & x2;
  assign n5527 = (n627 | n5528) & (~n1287 | ~n841);
  assign n5528 = (x0 | x1 | ~x5 | (~x2 ^ x4)) & (x5 | (x0 ? (x1 ? (x2 | x4) : (~x2 | ~x4)) : (x1 ? (~x2 | ~x4) : (x2 | x4))));
  assign n5529 = ~n5531 & (x6 | (~n5530 & (x1 | n5533)));
  assign n5530 = n733 & n757 & n774;
  assign n5531 = x3 & ((n728 & n733) | (x6 & ~n5532));
  assign n5532 = (x4 | x5 | x0 | x2) & (x1 | (x0 ? (~x2 | (~x4 ^ x5)) : (x5 ? ~x4 : (x2 & x4))));
  assign n5533 = (~x2 | n5534) & (x7 | n4129 | ~x0 | x2);
  assign n5534 = (~x0 | x3 | x4 | ~x5 | x7) & (x0 | ~x3 | ~x7 | (~x4 ^ ~x5));
  assign z290 = n5544 | (x3 ? (n5536 | ~n5538) : ~n5548);
  assign n5536 = ~x1 & ~n5537;
  assign n5537 = x0 ? (x4 | ~x5 | (x2 ^ ~x6)) : (~x4 | x5 | (~x2 ^ ~x6));
  assign n5538 = ~n5541 & ~n5542 & n5543 & (x1 | n5539);
  assign n5539 = (x0 | ~x4 | ~x5 | n3929) & (x5 | n5540 | ~x0 | x4);
  assign n5540 = x2 ? (~x6 | ~x7) : (x6 | x7);
  assign n5541 = ~x0 & ((n1145 & ~n3929) | (n632 & n1668));
  assign n5542 = ~n1580 & ~n5540;
  assign n5543 = (~n926 | ~n746) & (~n733 | ~n1725);
  assign n5544 = ~n643 & (n5546 | n5547 | (~x2 & ~n5545));
  assign n5545 = (x1 | ~x3 | ~x4 | ~x5) & (x5 | (x0 ? (x1 | (~x3 ^ x4)) : (~x1 | (x3 & ~x4))));
  assign n5546 = ~n1566 & ((x0 & ~n913) | (~n3802 & n1167));
  assign n5547 = n742 & ((n1121 & n927) | (~x1 & ~n856));
  assign n5548 = n5550 & n5554 & (~n1310 | n5549);
  assign n5549 = (~x4 | x6 | x7 | ~x1 | x2) & (x1 | x4 | ~x7 | (~x2 ^ ~x6));
  assign n5550 = (~x6 & (x5 | n5553)) | (~n5551 & ~n5552 & (n5553 | (~x5 & x6)));
  assign n5551 = ~x1 & ((x4 & x5 & ~x0 & x2) | (x0 & ~x4 & ~x5));
  assign n5552 = x5 & x4 & ~x2 & ~x0 & x1;
  assign n5553 = (x0 | ~x1 | x2 | x4 | x7) & (~x0 | x1 | ~x2 | ~x4 | ~x7);
  assign n5554 = (x6 | n5012) & (n714 | n5555);
  assign n5555 = x0 ? ((x1 | x6 | x7) & (~x1 | x2 | ~x6 | ~x7)) : (~x6 | ~x7 | (~x1 ^ ~x2));
  assign z291 = ~n5572 | ~n5563 | n5557 | n5560;
  assign n5557 = ~x1 & (~n5559 | (x3 & (n3175 | n5558)));
  assign n5558 = ~x2 & ((n1070 & n1167) | (x0 & ~n2055));
  assign n5559 = (n4226 | n4213) & (~n1783 | ~n993);
  assign n5560 = ~n1008 & ((n841 & ~n5562) | (~x0 & ~n5561));
  assign n5561 = x1 ? ((x2 | ~x3 | ~x4 | ~x6) & (~x2 | x3 | x4 | x6)) : ((x4 | x6 | x2 | x3) & (~x2 | ~x3 | (~x4 ^ x6)));
  assign n5562 = (x4 | x6 | x2 | x3) & (~x2 | ~x4 | (~x3 ^ ~x6));
  assign n5563 = ~n5564 & n5567 & ~n5569 & (n2063 | n5571);
  assign n5564 = ~n643 & ((n720 & ~n5565) | (~x2 & ~n5566));
  assign n5565 = x1 ? (~x3 | ~x5) : (x3 | x5);
  assign n5566 = (x0 | ((~x1 | x3 | x5) & (x1 | ~x3 | x4 | ~x5))) & (~x4 | ((~x1 | x3 | x5) & (~x0 | x1 | ~x3 | ~x5)));
  assign n5567 = (n1008 | n5568) & (x1 | n1014 | n3486);
  assign n5568 = x0 ? (x3 | x4 | (x1 ^ ~x2)) : (~x3 | ~x4 | (~x1 ^ ~x2));
  assign n5569 = x1 & ((~n4213 & ~n5570) | (n547 & n867));
  assign n5570 = x0 & x2;
  assign n5571 = (x0 | x1 | x2 | ~x3 | ~x4) & (~x0 | x3 | x4 | (x1 ^ ~x2));
  assign n5572 = (n1014 | n5573) & (~x1 | (~n609 & ~n5574));
  assign n5573 = (x1 | ((x2 | x3 | ~x6) & (~x0 | ~x2 | ~x3 | x6))) & (x0 | ~x1 | (x2 ? (x3 | ~x6) : (~x3 | x6)));
  assign n5574 = ~x0 & (~n4164 | (n1857 & ~n1150));
  assign z292 = ~n5585 | ~n5591 | (x1 ? ~n5576 : ~n5579);
  assign n5576 = ~n5374 & (x0 | (~x2 & n5577) | (x2 & n5578));
  assign n5577 = (~x3 | ~x4 | (x5 ? (x6 | ~x7) : (~x6 | x7))) & (x4 | ((~x6 | ~x7 | ~x3 | x5) & (x3 | (x5 ? ~x7 : (~x6 | x7)))));
  assign n5578 = (x4 | ~x5 | x6 | x7) & (x3 | ~x7 | (x4 ? (~x5 | x6) : (x5 | ~x6)));
  assign n5579 = ~n5582 & (x4 ? n5583 : n5580);
  assign n5580 = x6 ? n5581 : (~n3237 & (~n743 | ~n2575));
  assign n5581 = (x0 | x5 | (x2 ? (~x3 | x7) : (x3 | ~x7))) & (~x5 | ((~x0 | (x2 ? (~x3 | ~x7) : (x3 | x7))) & (x0 | x2 | ~x3 | x7)));
  assign n5582 = ~n981 & (x0 ? (x2 & ~n671) : (~x2 & ~n1218));
  assign n5583 = x0 ? (~n1044 | ~n658) : n5584;
  assign n5584 = (x2 | x3 | x5 | x6 | ~x7) & (~x2 | ~x3 | (x5 ? (x6 | x7) : (~x6 | ~x7)));
  assign n5585 = x5 ? (~n5590 & (~x2 | n5589)) : n5586;
  assign n5586 = x1 ? n5587 : n5588;
  assign n5587 = (x0 | ~x2 | x3 | x4 | x6) & (x2 | (x3 ? (x4 | x6) : (~x4 | ~x6)));
  assign n5588 = (x0 | ~x2 | ~x4 | x6) & (~x6 | ((~x3 | ~x4 | ~x0 | ~x2) & (x0 | x4 | (x2 ^ ~x3))));
  assign n5589 = (x4 | x6 | ~x0 | x1) & (x0 | ((x1 | ~x3 | ~x4 | ~x6) & (~x1 | ((x4 | ~x6) & (~x3 | ~x4 | x6)))));
  assign n5590 = x4 & n804 & (x0 ? x6 : (~x3 & ~x6));
  assign n5591 = ~n5592 & (n640 | (~x0 & n5595) | (x0 & n5596));
  assign n5592 = ~n643 & (x2 ? ~n5593 : ~n5594);
  assign n5593 = (x0 | ~x1 | ~x4 | x5) & (x1 | (x0 ? (x3 ? (~x4 | ~x5) : (x4 | x5)) : (x4 | ~x5)));
  assign n5594 = (~x1 | x3 | ~x4 | ~x5) & (~x0 | x1 | x5 | (~x3 ^ x4));
  assign n5595 = (x1 | ~x2 | x3 | ~x4 | ~x5) & (~x3 | ((~x1 | x4 | (x2 ^ ~x5)) & (x1 | x2 | ~x4 | ~x5)));
  assign n5596 = (~x1 | x2 | x3 | x4 | ~x5) & (x1 | x5 | (x2 ? (x3 | ~x4) : (~x3 ^ ~x4)));
  assign z293 = ~n5610 | n5606 | n5604 | n5598 | n5601;
  assign n5598 = ~x1 & (n5599 | (n830 & n1783));
  assign n5599 = x4 & ((n978 & n2435) | (n1769 & ~n5600));
  assign n5600 = (x0 | ~x2 | x3 | ~x5) & (~x0 | x5 | (~x2 ^ ~x3));
  assign n5601 = ~n1198 & (n5602 | (~x3 & ~n5603));
  assign n5602 = x3 & ((~x0 & x1 & ~x2 & x7) | (~x1 & (x0 ? (x2 & ~x7) : (x2 ^ ~x7))));
  assign n5603 = (~x0 | ~x1 | x2 | x4 | x7) & (x0 | ((x1 | x2 | ~x4 | x7) & (x4 | ~x7 | ~x1 | ~x2)));
  assign n5604 = ~x7 & ((n1268 & n1269) | (x1 & ~n5605));
  assign n5605 = (x0 | ~x2 | ~x3 | ~x4 | ~x5) & (~x0 | x2 | x5 | (~x3 ^ x4));
  assign n5606 = ~n1097 & (n5608 | (~n5607 & (~x3 | n774)));
  assign n5607 = (x0 | (x1 ? (~x2 | x7) : (x2 | ~x7))) & (~x2 | ~x7 | ~x0 | x1);
  assign n5608 = n1084 & ((n543 & n683) | (x0 & n5609));
  assign n5609 = ~x1 & (~x3 ^ ~x7);
  assign n5610 = n5612 & ~n5613 & n5614 & (n3309 | n5611);
  assign n5611 = (~x0 | x1 | ~x3 | ~x4 | ~x5) & (x0 | x3 | (x1 ? (~x4 | x5) : (x4 | ~x5)));
  assign n5612 = (n1246 | n1387) & (~n526 | ~n1029 | ~n816);
  assign n5613 = n543 & n778 & (n923 | n1598);
  assign n5614 = (n3924 | ~n1283) & (~n841 | n5615);
  assign n5615 = (~x2 | x3 | ~x5 | x7) & (x2 | ~x3 | x5 | ~x7);
  assign z294 = n5632 | n5628 | ~n5617 | ~n5621;
  assign n5617 = n5619 & (~n5260 | n5618);
  assign n5618 = (x2 | x3 | ~x4 | ~x5 | x7) & (~x2 | x5 | (x3 ? (~x4 | x7) : (x4 | ~x7)));
  assign n5619 = (n1171 | n1682) & (~n632 | n5620);
  assign n5620 = (~x0 | ~x3 | x4 | x5 | x6) & (x0 | ~x6 | (x3 ? (~x4 | ~x5) : (x4 | x5)));
  assign n5621 = ~n5622 & ~n5625 & (~x4 | n5624);
  assign n5622 = ~n643 & ((x3 & ~n5623) | (x1 & ~x3 & ~n5194));
  assign n5623 = (x0 | ~x1 | ~x2 | x4 | x5) & (x1 | (x0 ? (x2 ? (~x4 | ~x5) : x4) : (x2 | ~x4)));
  assign n5624 = (x0 | x1 | x2 | x3 | ~x6) & (x6 | ((x2 | x3 | ~x0 | ~x1) & (x0 | ~x2 | (~x1 ^ ~x3))));
  assign n5625 = ~x1 & ((n1051 & ~n5626) | (n825 & n5627));
  assign n5626 = (x0 | ~x2 | x4 | ~x5) & (~x0 | (x2 ? (x4 | x5) : (~x4 | ~x5)));
  assign n5627 = x6 & (x2 ? (x4 & x5) : (~x4 & ~x5));
  assign n5628 = ~n640 & (~n5631 | (~x1 & (~n5629 | ~n5630)));
  assign n5629 = (x0 | ~x2 | ~x3 | ~x4 | x5) & (x3 | ((x0 | x2 | x4 | ~x5) & (~x0 | (x2 ? (x4 | ~x5) : (~x4 | x5)))));
  assign n5630 = (x0 | ~x2 | ~x3 | x4) & (~x0 | x3 | (~x2 ^ ~x4));
  assign n5631 = (~n543 | ~n949) & (~n733 | ~n1641);
  assign n5632 = ~x0 & ((~n3855 & n4569) | (~x4 & ~n5633));
  assign n5633 = (x5 | ~x7 | ~n689 | n815) & (~x5 | n5634);
  assign n5634 = (x1 | x2 | ~x3 | ~x6 | x7) & (~x1 | ((x2 | x3 | ~x6 | x7) & (x6 | ~x7 | ~x2 | ~x3)));
  assign z295 = ~n5645 | n5642 | n5636 | n5639;
  assign n5636 = ~x0 & ((~n976 & ~n2693) | (~x1 & ~n5637));
  assign n5637 = x7 ? (~x2 | (~n1748 & ~n5137)) : n5638;
  assign n5638 = (x2 | ~x3 | x4 | ~x5 | x6) & (x3 | ((~x2 | (x4 ? (~x5 | x6) : (x5 | ~x6))) & (x5 | ~x6 | x2 | ~x4)));
  assign n5639 = ~x5 & (x3 ? ~n5640 : ~n5641);
  assign n5640 = x2 ? ((~x0 | x1 | ~x4 | x7) & (x0 | ~x1 | x4 | ~x7)) : ((x0 | ~x1 | ~x4 | ~x7) & (x4 | (x0 ? (x1 ^ ~x7) : (x1 | x7))));
  assign n5641 = (~x0 | ~x1 | x2 | x4 | ~x7) & (x1 | ~x2 | (x0 ? (~x4 ^ ~x7) : (~x4 | x7)));
  assign n5642 = x0 & ((n576 & n1725) | (~x1 & ~n5643));
  assign n5643 = (x4 | n5644) & (~x2 | ~x4 | ~x7 | n975);
  assign n5644 = (~x2 | x3 | x5 | ~x6 | ~x7) & (x2 | x6 | (x3 ? (~x5 | ~x7) : (x5 | x7)));
  assign n5645 = ~n5646 & ~n5649 & ~n5650 & (x0 | n5648);
  assign n5646 = x5 & ((n733 & n3090) | (~x1 & ~n5647));
  assign n5647 = (x0 | x2 | x3 | ~x4 | x7) & (~x2 | (~x3 ^ ~x4) | (~x0 ^ ~x7));
  assign n5648 = (x1 | x2 | x3 | x4 | ~x7) & (~x1 | (x2 ? (~x4 | (~x3 ^ x7)) : (x4 | (~x3 ^ ~x7))));
  assign n5649 = ~n1532 & ((n841 & n1903) | (~x0 & ~n5144));
  assign n5650 = n793 & (n619 | n5651);
  assign n5651 = ~x7 & x1 & x4;
  assign z296 = ~n5664 | n5661 | n5653 | n5656;
  assign n5653 = ~x2 & (n5654 | (n610 & n1734));
  assign n5654 = ~x1 & ((n5168 & n951) | (x0 & ~n5655));
  assign n5655 = (x3 | x4 | x5 | x6 | ~x7) & (~x5 | ((x3 | (x4 ? (x6 | ~x7) : (~x6 | x7))) & (~x3 | ~x4 | x6 | x7)));
  assign n5656 = x2 & (n5657 | (~x3 & ~n5659));
  assign n5657 = x3 & ((~x1 & ~n2055) | (~x0 & x1 & ~n5658));
  assign n5658 = (~x4 | x5 | ~x6 | x7) & (x4 | ~x5 | x6 | ~x7);
  assign n5659 = (x4 | ~n1070 | ~x0 | x1) & (x0 | ~x1 | n5660);
  assign n5660 = (x4 | x5 | ~x6 | x7) & (~x4 | (x5 ? (~x6 | x7) : (x6 | ~x7)));
  assign n5661 = ~x3 & (~n5663 | (~x0 & ~n5662));
  assign n5662 = (x1 | ~x2 | ~x4 | ~x5 | ~x6) & (x5 | (x1 ? (x6 | (x2 ^ ~x4)) : (~x6 | (x2 & x4))));
  assign n5663 = (n1198 | n3956) & (~n559 | ~n560);
  assign n5664 = n5666 & (~n825 | n5665);
  assign n5665 = (x1 | x2 | x4 | ~x5 | ~x6) & (~x1 | ((~x2 | (x4 ? (x5 | x6) : (~x5 | ~x6))) & (x2 | x4 | ~x5 | x6)));
  assign n5666 = (~x3 | n5669) & (x3 | n5667) & (n2063 | n5668);
  assign n5667 = (~x0 | ~x1 | x2 | ~x4 | x5) & (x1 | ~x5 | ((~x2 | x4) & (x0 | x2 | ~x4)));
  assign n5668 = (~x1 | x2 | x3 | x4) & (~x0 | x1 | (x2 ? (x3 | ~x4) : (~x3 | x4)));
  assign n5669 = (x1 | x2 | ~x4 | x5) & ((~x4 ^ ~x5) | ((x1 | ~x2) & (x0 | ~x1 | x2)));
  assign z297 = ~n5680 | n5671 | ~n5676;
  assign n5671 = ~n1097 & (~n5673 | (x0 & ~n5672));
  assign n5672 = (x3 | ~x4 | ~x1 | x2) & (x1 | ((~x2 | (x3 ? x4 : (~x4 | ~x7))) & (~x3 | (x4 ? x2 : ~x7))));
  assign n5673 = ~n5674 & ~n5675 & (~n1269 | ~n2648);
  assign n5674 = x7 & ((~x3 & ~x4 & x0 & ~x2) | (~x0 & ((x3 & ~x4) | (x2 & ~x3 & x4))));
  assign n5675 = ~x0 & x3 & ~x7 & (~x2 | ~x4);
  assign n5676 = ~n5677 & (~n1986 | (~n5679 & (~n570 | ~n2089)));
  assign n5677 = x1 & (x0 ? (n704 & n1044) : ~n5678);
  assign n5678 = (~x4 | (x3 ? (~x5 | x6) : (x5 | ~x6))) & (x3 | ((x2 | x5 | ~x6) & (~x2 | x4 | ~x5 | x6)));
  assign n5679 = ~x2 & (~n2077 | (n689 & n577));
  assign n5680 = ~n5681 & (~x7 | (~n5684 & ~n5686));
  assign n5681 = ~x1 & (x0 ? ~n5682 : ~n5683);
  assign n5682 = (x5 | ((~x2 | x3 | ~x4 | ~x6) & (x2 | ((x4 | ~x6) & (x3 | ~x4 | x6))))) & (~x2 | ~x5 | x6 | (~x3 ^ ~x4));
  assign n5683 = (~x3 | ~x4 | ~x5 | x6) & (x3 | ((x2 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (x5 | ~x6 | ~x2 | x4)));
  assign n5684 = ~x0 & ((x1 & ~x2 & ~n928) | (x2 & ~n5685));
  assign n5685 = (~x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (~x1 | x3 | x4 | x5 | ~x6);
  assign n5686 = x0 & ((n576 & n1358) | (~x1 & ~n5687));
  assign n5687 = (~x5 | x6 | x2 | ~x4) & (~x2 | ((~x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (x5 | ~x6 | x3 | x4)));
  assign z298 = n5689 | ~n5692 | n5697 | (~n1116 & ~n5696);
  assign n5689 = ~n1008 & ((~n784 & ~n5690) | (~x3 & ~n5691));
  assign n5690 = x0 ? (x1 | x4) : (~x3 ^ ~x4);
  assign n5691 = (x2 | ~x4 | ~x6 | (x0 & ~x1)) & (x6 | ((~x2 | ~x4 | x0 | ~x1) & (~x0 | (x1 ? (x2 | x4) : (~x2 | ~x4)))));
  assign n5692 = ~n5694 & n5695 & (n5693 | (n1701 & n1097));
  assign n5693 = (~x0 | x1 | ~x2 | ~x3 | ~x4) & (x0 | ((x2 | ~x3 | x4) & (x1 | ~x2 | x3 | ~x4)));
  assign n5694 = ~n5361 & (x0 ? (~x1 & ~x4) : ((~x3 & ~x4) | (~x1 & x3 & x4)));
  assign n5695 = (~n601 | ~n880) & (~n1549 | n5179);
  assign n5696 = (x1 & (x3 ? x0 : x2)) | (x0 & ~x3 & (x2 | (~x1 & x4))) | (x2 & x4) | (~x2 & ~x4 & (~x0 | x3));
  assign n5697 = x4 & ((n746 & n2409) | (~x3 & ~n5698));
  assign n5698 = (n823 | n3855) & (x7 | ~n743 | n5699);
  assign n5699 = x1 ? (x5 | x6) : (~x5 | ~x6);
  assign z299 = n5701 | ~n5707 | ~n5717 | (n841 & ~n5712);
  assign n5701 = ~x0 & (n5702 | (x7 & (n5705 | ~n5706)));
  assign n5702 = ~x7 & (x2 ? ~n5703 : ~n5704);
  assign n5703 = (x3 | ((x4 | ~x5 | x6) & (x5 | ~x6 | ~x1 | ~x4))) & (x1 | ~x3 | (x4 ? (~x5 | x6) : (~x5 ^ ~x6)));
  assign n5704 = (x1 | ~x3 | x4 | (~x5 ^ ~x6)) & (x3 | ((x4 | ~x5 | x6) & (~x1 | ((~x4 | x5 | ~x6) & (~x5 | x6)))));
  assign n5705 = ~x1 & (n606 | (n1723 & (n949 | n5101)));
  assign n5706 = (~n559 | ~n2135) & (n1097 | n2965);
  assign n5707 = ~n5710 & (x3 | (~n5708 & (x0 | n5709)));
  assign n5708 = ~n1954 & (x0 ? (n2317 | (x4 & n526)) : (~x4 & n526));
  assign n5709 = (~x5 | ~x7 | ~x1 | ~x4) & (x1 | ((~x4 | x5 | x7) & (~x5 | ~x7 | x2 | x4)));
  assign n5710 = ~n2803 & ~n5711;
  assign n5711 = (x0 | ~x1 | ~x3 | x5) & (~x0 | x3 | ~x5 | (x1 ^ ~x2));
  assign n5712 = ~n5713 & n5715 & (x7 | ~n681 | n5714);
  assign n5713 = ~n640 & (n2775 | (n1477 & n885));
  assign n5714 = (~x2 | x3 | x6) & (~x3 | ~x6);
  assign n5715 = (n3319 | n5716) & (~n530 | ~n2385);
  assign n5716 = (~x3 | ~x5) & (x2 | x3 | x5);
  assign n5717 = ~n5718 & ~n5720;
  assign n5718 = x3 & ((n837 & n2209) | (~x0 & ~n5719));
  assign n5719 = (x5 | x7 | ~x1 | x4) & (~x4 | ((x2 | ~x5 | x7) & (~x1 | (~x5 ^ x7))));
  assign n5720 = ~n643 & (x3 ? (n2332 & n543) : ~n5721);
  assign n5721 = (x0 | x1 | ~x2 | ~x4 | ~x5) & (x5 | (x0 ? (~x4 | (x1 ^ ~x2)) : (x4 | (x1 & x2))));
  assign z300 = n5723 | n5730 | ~n5732 | (x1 & ~n5727);
  assign n5723 = ~x0 & (n5724 | (n1723 & ~n5726));
  assign n5724 = x5 & ((n3236 & ~n2541) | (~x6 & ~n5725));
  assign n5725 = x1 ? (x2 | (x3 ? (x4 | x7) : ~x7)) : (~x2 | ((~x3 | x4 | ~x7) & (~x4 | x7)));
  assign n5726 = (~x1 | x2 | x3 | x4 | x7) & (x1 | (~x2 & ~x3) | (~x4 ^ ~x7));
  assign n5727 = (x2 | n5729) & (x0 | ~x2 | ~x5 | n5728);
  assign n5728 = (~x4 | x6) & (x3 | x4 | ~x6);
  assign n5729 = x0 ? (x5 | ((x4 | x6) & (x3 | ~x4 | ~x6))) : (~x3 | ~x5 | (~x4 ^ x6));
  assign n5730 = ~x1 & ((n859 & ~n4024) | (~x2 & ~n5731));
  assign n5731 = x0 ? (~x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))) : (x5 | ((~x4 | x6) & (x3 | x4 | ~x6)));
  assign n5732 = ~n5733 & ~n5739 & (n643 | (~n5736 & n5737));
  assign n5733 = n841 & (x6 ? (n691 & ~n5735) : ~n5734);
  assign n5734 = (x2 | x3 | ~x4 | ~x5 | x7) & (x5 | ((~x2 | ((x4 | ~x7) & (x3 | ~x4 | x7))) & (~x3 | ((x4 | ~x7) & (x2 | ~x4 | x7)))));
  assign n5735 = x3 ? (x4 | ~x7) : x7;
  assign n5736 = x4 & n743 & (x1 ? (~x3 & x5) : (x3 ^ ~x5));
  assign n5737 = ~n3915 & ~n5738 & (~n1311 | ~n1269);
  assign n5738 = ~x0 & ((x1 & x4 & ~x5) | (~x4 & x5 & ~x1 & ~x2));
  assign n5739 = ~n640 & (~n5741 | (n1084 & ~n5740));
  assign n5740 = (x0 | ~x1 | ~x3 | x5) & (~x0 | x3 | (~x1 ^ ~x5));
  assign n5741 = (x0 | ((~x4 | ~x5 | x1 | x2) & (x4 | x5 | ~x1 | ~x2))) & (~x0 | x1 | ~x2 | x4 | ~x5);
  assign z301 = n5743 | ~n5747 | ~n5751 | (~x0 & ~n5746);
  assign n5743 = ~x1 & (n5744 | (n1241 & n1783));
  assign n5744 = ~x2 & ((n942 & n5168) | (n1479 & ~n5745));
  assign n5745 = (~x0 | (x3 ? (x5 | ~x7) : (~x5 | x7))) & (x0 | x3 | ~x5 | ~x7);
  assign n5746 = (~x1 | x2 | ~x3 | x5 | ~x7) & (~x2 | ((x5 | x7 | x1 | x3) & (~x1 | ((~x5 | x7) & (x3 | x5 | ~x7)))));
  assign n5747 = ~n5748 & ~n5750 & (n3924 | n1350);
  assign n5748 = ~n5749 & x4 & n632;
  assign n5749 = (x0 | (x3 ? (~x5 | x7) : (x5 | ~x7))) & (~x5 | ~x7 | ~x0 | x3);
  assign n5750 = x0 & ((n632 & n4531) | (n570 & n2575));
  assign n5751 = ~n5752 & ~n5754 & (n1097 | (~n5756 & n5757));
  assign n5752 = ~n1198 & ((n733 & n2647) | (~x1 & ~n5753));
  assign n5753 = (~x7 & (~x0 | (x2 & x3 & x4))) | (~x2 & ~x3) | (x0 & x7);
  assign n5754 = ~x1 & ((n3434 & n867) | (~x2 & ~n5755));
  assign n5755 = (x5 | x7 | x0 | ~x4) & (~x0 | ~x5 | (x3 ? (~x4 | ~x7) : (x4 | x7)));
  assign n5756 = ~x0 & ((~x1 & x2 & x3 & ~x7) | (x1 & (x2 ? (x3 & x7) : (~x3 & ~x7))));
  assign n5757 = (~n841 | ~n5758) & (x4 | ~n902 | n3134);
  assign n5758 = x7 & ~x2 & ~x3;
  assign z302 = n5760 | n5763 | ~n5768 | (~n640 & ~n5766);
  assign n5760 = ~x2 & (n5761 | (n610 & n661));
  assign n5761 = ~x0 & ((n530 & n944) | (~x4 & ~n5762));
  assign n5762 = (x1 | x3 | x5 | x6 | ~x7) & (~x1 | ~x5 | (x3 ? (x6 | ~x7) : (~x6 | x7)));
  assign n5763 = ~x2 & ((x0 & ~n5764) | (n3074 & ~n5765));
  assign n5764 = x1 ? (x3 | x6) : (~x6 | (~x3 ^ (x4 & x5)));
  assign n5765 = x1 ? (~x3 | ~x4) : (x3 | (~x4 & ~x5));
  assign n5766 = ~n1613 & ~n5767 & (x5 | n1998 | ~n4569);
  assign n5767 = ~x0 & (x1 ? (x2 & x3) : (x2 ? (~x3 & ~x4) : x3));
  assign n5768 = ~n5771 & (n5769 | n5770) & (~x2 | n5773);
  assign n5769 = (x4 | x5 | ~x1 | x2) & (~x4 | ~x5 | x1 | ~x2);
  assign n5770 = x0 ? (~x3 | x6) : (x3 | ~x6);
  assign n5771 = ~n643 & (~n5772 | (n902 & ~n1939));
  assign n5772 = (x0 | ~x1 | x2 | x3 | ~x4) & (~x0 | x1 | ~x2 | (x3 & x4));
  assign n5773 = (x0 | (x1 ? (x3 | x6) : (~x3 | ~x6))) & (~x0 | x1 | ~x3 | ~n926);
  assign z303 = ~n5779 | ~n5783 | (~x2 & (~n5775 | ~n5778));
  assign n5775 = (~x0 | ~n5776) & (x4 | n5777);
  assign n5776 = ~x1 & x4 & (x3 ? (x5 ^ ~x7) : (~x5 & x7));
  assign n5777 = (~x0 | ~x1 | ~x3 | x5 | x7) & (x0 | ((x1 | x3 | ~x5 | x7) & (x5 | ~x7 | ~x1 | ~x3)));
  assign n5778 = (x0 | x3 | x7 | (~x1 ^ x4)) & ((x0 ? (x1 | x4) : (~x1 | ~x4)) | (~x3 ^ x7));
  assign n5779 = ~n5780 & ~n5781 & ~n5782 & (~n1269 | ~n5290);
  assign n5780 = ~x3 & ((~x0 & x1 & x2 & ~x7) | (x0 & (x1 ? (~x2 & ~x7) : (x2 & x7))));
  assign n5781 = ~x0 & x3 & (x1 ? (x2 & x7) : (x2 ^ x7));
  assign n5782 = n1241 & n2144;
  assign n5783 = (x0 | n5784) & (~n570 | (~n900 & (~x0 | ~n5212)));
  assign n5784 = (n538 | n5785) & (n5786 | ~n5787);
  assign n5785 = (x1 | x3 | ~x4 | ~x7) & (x4 | x7 | ~x1 | ~x3);
  assign n5786 = x1 ? (~x5 | ~x7) : (x5 | x7);
  assign n5787 = x6 & ~x4 & ~x2 & ~x3;
  assign z304 = x7 ? (~n553 | ~n5789) : ~n5791;
  assign n5789 = (~n746 | ~n2145) & (x3 | (~n5790 & (~n696 | ~n746)));
  assign n5790 = ~n2341 & ((~x4 & x5 & x1 & ~x2) | (~x1 & x4 & (x2 ^ x5)));
  assign n5791 = n5794 & (x0 | n5792) & (x6 | n5793);
  assign n5792 = (~x1 | ((~x3 | ~x4) & (~x2 | x3 | x4 | x5))) & (~x3 | (x2 ? (x4 | ~x5) : (~x4 | x5))) & (x1 | ((~x3 | x4) & (~x2 | x3 | ~x4 | ~x5)));
  assign n5793 = (~n622 | n1284) & (~x4 | n968 | ~n1922);
  assign n5794 = (~x6 | n968 | ~n3047) & (~x0 | n5795);
  assign n5795 = (~x1 | x2 | x3 | x4 | x5) & (x1 | ((~x3 | ~x4 | ~x5) & (~x2 | (~x3 ^ ~x4))));
  assign z305 = ~n5807 | ~n5806 | n5804 | n5797 | n5801;
  assign n5797 = ~x6 & (n5798 | (~x5 & n885 & ~n5800));
  assign n5798 = ~x2 & ((n2296 & n1244) | (x5 & ~n5799));
  assign n5799 = x0 ? (x7 | (x1 ? (x3 | ~x4) : (~x3 | x4))) : (~x3 | ~x7 | (~x1 ^ x4));
  assign n5800 = (x4 | x7 | ~x0 | x1) & (x0 | ~x7 | (x1 ^ ~x4));
  assign n5801 = x6 & (n5803 | (n5802 & n816));
  assign n5802 = x7 & x5 & ~x3 & x4;
  assign n5803 = x2 & ((n635 & n1244) | (~n1920 & ~n3961));
  assign n5804 = ~n968 & ~n5805;
  assign n5805 = (x0 | ~x1 | (x3 ? (x4 | ~x6) : (~x4 | x6))) & (x1 | (~x4 ^ ~x6) | (x0 ^ ~x3));
  assign n5806 = (~x0 | x1 | x2 | x4 | x5) & (x0 | ((x1 | ~x2 | ~x4 | ~x5) & (~x1 | (x2 ? (x4 | ~x5) : (~x4 | x5)))));
  assign n5807 = n5810 & (x1 | n5808) & (~n1875 | n5809);
  assign n5808 = (x0 | ~x2 | x3 | x4 | x5) & (~x0 | x2 | ~x3 | ~x4 | ~x5) & ((~x3 ^ x5) | (x0 ? (~x2 | ~x4) : (x2 | x4)));
  assign n5809 = (x1 | ~x2 | ~x3 | ~x4 | x6) & (~x1 | x2 | x3 | x4 | ~x6);
  assign n5810 = (~n1268 | ~n837) & (~n816 | ~n1228);
  assign z306 = ~n5820 | (x0 ? (n5816 | n5818) : ~n5812);
  assign n5812 = ~n5815 & (~n1084 | n5813) & (n627 | n5814);
  assign n5813 = x1 ? ((x3 | x5 | ~x6 | x7) & (x6 | ~x7 | ~x3 | ~x5)) : ((~x3 | x5 | ~x6 | x7) & (x3 | x6 | (~x5 ^ x7)));
  assign n5814 = x5 ? ((~x2 | x4 | x7) & (x1 | x2 | ~x4 | ~x7)) : ((x1 | ~x2 | ~x4 | ~x7) & (~x1 | (x2 ? (x4 | ~x7) : (~x4 | x7))));
  assign n5815 = x2 & ((n813 & n3192) | (n530 & n1288));
  assign n5816 = ~n765 & ~n5817;
  assign n5817 = (~x1 | x2 | x3 | ~x4 | x6) & (x1 | ~x3 | (x2 ? (~x4 | ~x6) : (x4 | x6)));
  assign n5818 = ~x1 & ((n3431 & ~n4754) | (x6 & ~n5819));
  assign n5819 = (~x2 | x3 | x4 | x5 | ~x7) & (x2 | x7 | (x3 ? (~x4 | ~x5) : (x4 | x5)));
  assign n5820 = (x2 & n5825) | (~x2 & ~n5821 & ~n5823 & n5824);
  assign n5821 = ~x3 & ~n5822;
  assign n5822 = x0 ? ((x4 | ~x5 | ~x6) & (x1 | ~x4 | x5 | x6)) : (~x4 | x5 | (x1 ^ ~x6));
  assign n5823 = ~n1408 & ((n1301 & n841) | (~x0 & ~n5565));
  assign n5824 = (x0 | ~x3 | (n2819 & (x1 | n2259))) & (x3 | n2819 | (~x0 & ~x1));
  assign n5825 = (x0 | ((~n4894 | n975) & (~x1 | n5826))) & (x1 | (x0 ? n5826 : n975));
  assign n5826 = (x3 | x4 | ~x5 | x6) & (x5 | (x3 ? (~x4 ^ x6) : (~x4 | ~x6)));
  assign z307 = ~n5841 | (x2 ? (n5834 | ~n5837) : ~n5828);
  assign n5828 = x3 ? n5831 : (x1 ? n5829 : n5830);
  assign n5829 = x7 ? (x0 ? (~x4 | x6) : (x5 | ~x6)) : (x0 ? (~x6 | (x4 ^ ~x5)) : (x6 | (~x4 & ~x5)));
  assign n5830 = ((x0 ? (x4 | x5) : (~x4 | ~x5)) | (~x6 ^ ~x7)) & (~x0 | ~x4 | x5 | ~x6 | x7) & (x0 | x4 | ((x6 | ~x7) & (x5 | ~x6 | x7)));
  assign n5831 = (n643 | n5832) & (x1 | n5833);
  assign n5832 = x0 ? (x1 | x4) : (x1 ? (~x4 ^ x5) : (~x4 | ~x5));
  assign n5833 = (x0 | x4 | x5 | x6 | x7) & (~x6 | ((~x0 | ~x4 | ~x5 | ~x7) & (x0 | x5 | (x4 ^ ~x7))));
  assign n5834 = ~x1 & ((~x5 & ~n5836) | (~x0 & n5835));
  assign n5835 = ~x3 & x5 & (x4 ? (~x6 & ~x7) : (x6 & x7));
  assign n5836 = (x0 | x3 | x4 | x6 | ~x7) & (~x0 | ((x3 | ~x4 | ~x6 | x7) & (~x3 | x4 | x6 | ~x7)));
  assign n5837 = ~n5840 & (x6 ? (x7 ? n5839 : n5838) : (x7 ? n5838 : n5839));
  assign n5838 = (x1 | ~x4 | (x0 ? (x3 | ~x5) : (~x3 | x5))) & (x0 | ~x3 | x4 | (~x1 & ~x5));
  assign n5839 = (x0 | ~x1 | ~x5 | (~x3 ^ ~x4)) & (x1 | ((x0 | x3 | ~x4 | x5) & (~x0 | (x3 ? ~x4 : (x4 | x5)))));
  assign n5840 = ~n2803 & n543 & ~x3 & ~x5;
  assign n5841 = ~n5844 & (~n543 | n5842) & (n627 | n5843);
  assign n5842 = (x2 | ~x3 | x4 | x5 | ~x6) & (x3 | ((x4 | x5 | x6) & (~x5 | ~x6 | ~x2 | ~x4)));
  assign n5843 = x0 ? ((~x1 | x2 | x4 | x5) & (x1 | ~x5 | (~x2 ^ x4))) : (~x4 | (x1 ? (~x2 ^ x5) : (~x2 | ~x5)));
  assign n5844 = ~x1 & ((n742 & n5846) | (~x2 & ~n5845));
  assign n5845 = x0 ? ((~x5 | ~x6 | x3 | x4) & (x5 | x6 | ~x3 | ~x4)) : ((~x3 | x4 | ~x5 | ~x6) & (x3 | ~x4 | x5 | x6));
  assign n5846 = ~x4 & (x3 ? (~x5 & x6) : (x5 & ~x6));
  assign z308 = n5857 | ~n5861 | (x2 ? ~n5853 : ~n5848);
  assign n5848 = n5851 & (~x5 | n5849);
  assign n5849 = (x1 | n5850) & (~n873 | (~n1395 & ~n2724));
  assign n5850 = x0 ? ((x3 | ~x4 | ~x6 | x7) & (~x3 | x4 | x6 | ~x7)) : (x3 | x4 | (~x6 ^ x7));
  assign n5851 = (n5852 | n4910) & (n640 | n2528 | n2585);
  assign n5852 = x1 ? (~x5 | x7) : (x5 | ~x7);
  assign n5853 = ~n5854 & (x1 | (n5856 & (n3345 | n2129)));
  assign n5854 = ~n671 & ~n5855;
  assign n5855 = (~x3 | x5 | x6 | ~x0 | x1) & (x0 | ((~x5 | ~x6 | x1 | x3) & (~x1 | (x3 ? (~x5 | x6) : (x5 | ~x6)))));
  assign n5856 = (~n2857 | ~n658) & (~n1070 | ~n2094);
  assign n5857 = ~x1 & (n5859 | n5860 | (~x3 & ~n5858));
  assign n5858 = (~x0 | x2 | x4 | ~x5 | x7) & (x0 | ((x2 | ~x4 | ~x5 | ~x7) & (~x2 | (x4 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n5859 = ~n671 & (x0 ? (~x5 & ~n5064) : ~n1515);
  assign n5860 = ~n1337 & x3 & n995;
  assign n5861 = ~n5862 & (n1218 | (~n3464 & (~n622 | n753)));
  assign n5862 = x1 & ((n594 & n2209) | (~x0 & ~n5863));
  assign n5863 = ((~x4 ^ x7) | (x2 ? (~x3 ^ x5) : (~x3 | ~x5))) & (x2 | x3 | ~x4 | x5 | ~x7) & (~x2 | ((~x5 | ~x7 | ~x3 | ~x4) & (x5 | x7 | x3 | x4)));
  assign z309 = n5876 | ~n5878 | (x1 ? ~n5871 : ~n5865);
  assign n5865 = x3 ? n5868 : (x5 ? n5866 : n5867);
  assign n5866 = (~x4 | x6 | x7 | ~x0 | x2) & (x0 | ~x2 | x4 | ~x6 | ~x7);
  assign n5867 = x0 ? (x4 ? (~x6 | ~x7) : (x6 | x7)) : (x4 ? (x7 | (~x2 ^ ~x6)) : (x6 | ~x7));
  assign n5868 = (~x7 | n5869) & (~x5 | x7 | n5870);
  assign n5869 = (x4 | ((~x5 | ~x6 | ~x0 | x2) & (x0 | (x2 ? (~x5 | x6) : (x5 | ~x6))))) & (~x0 | ~x2 | ~x4 | (~x5 ^ ~x6));
  assign n5870 = (x0 | x2 | (~x4 ^ x6)) & (~x2 | (x0 ? (x4 | x6) : (~x4 | ~x6)));
  assign n5871 = ~n5872 & ~n5875 & (~n600 | ~n830);
  assign n5872 = ~x0 & ((x7 & ~n5873) | (n1379 & ~n5874));
  assign n5873 = (~x2 | x3 | x4 | x5 | ~x6) & (x6 | ((x2 | ~x3 | x4 | ~x5) & (~x2 | ~x4 | (~x3 ^ ~x5))));
  assign n5874 = (~x2 | x3 | ~x5 | x6) & (x2 | ~x6 | (~x3 ^ ~x5));
  assign n5875 = ~n765 & ((n742 & n1141) | (n743 & n1331));
  assign n5876 = x0 & (x1 ? (n1044 & n559) : ~n5877);
  assign n5877 = (~x2 | (x3 ? (x5 | ~x6) : (~x5 | x6))) & (x4 | ((x3 | ~x5) & (x2 | ~x3 | x5)));
  assign n5878 = (n1097 | n5879) & (x0 | (~n5880 & n5881));
  assign n5879 = (x2 | (x0 ? (x1 ? (x3 | x4) : (~x3 | ~x4)) : (~x1 | (~x3 ^ x4)))) & (x0 | ~x2 | (x1 ? (~x3 | ~x4) : (~x3 ^ x4)));
  assign n5880 = ~x4 & ((n1746 & n804) | (n4137 & ~n4336));
  assign n5881 = ~n5882 & (n1480 | n1100) & (n1954 | n5239);
  assign n5882 = x5 & x4 & ~x3 & ~x1 & ~x2;
  assign z310 = ~n5898 | n5896 | n5892 | n5884 | ~n5887;
  assign n5884 = n1167 & (n5885 | (~x5 & n570 & ~n871));
  assign n5885 = ~x2 & (n5886 | (n1317 & n2862));
  assign n5886 = x7 & x6 & ~x5 & ~x1 & x3;
  assign n5887 = ~n5890 & (n640 | (~x1 & n5888) | (x1 & n5889));
  assign n5888 = (x2 | ~x3 | x4 | ~x5) & (~x4 | ((~x0 | x3 | x5) & (~x2 | ((x3 | x5) & (x0 | ~x3 | ~x5)))));
  assign n5889 = (~x0 | x2 | x3 | x4 | x5) & (x0 | (~x3 ^ ~x5) | (~x2 ^ x4));
  assign n5890 = ~n3309 & ((~x1 & ~n5891) | (~x0 & x1 & ~n2077));
  assign n5891 = (x0 | x3 | x4 | ~x5 | ~x6) & (~x0 | ~x3 | ~x4 | (~x5 ^ ~x6));
  assign n5892 = ~n643 & (~n5894 | (~x2 & ~n5893));
  assign n5893 = (x0 | ~x1 | ~x3 | x4 | ~x5) & (~x0 | x3 | x5 | (~x1 ^ ~x4));
  assign n5894 = (~n639 | ~n1269) & (n877 | (~n1931 & ~n5895));
  assign n5895 = ~x0 & x4 & (x1 ^ ~x2);
  assign n5896 = ~x1 & ((n704 & n547) | ~n3424 | n5897);
  assign n5897 = ~n647 & ((~x2 & ~x6) | (x0 & x2 & x6));
  assign n5898 = ~n5899 & ~n5900 & (~n1121 | ~n622 | n5901);
  assign n5899 = ~n981 & ((n922 & n1084) | (~x0 & ~n4121));
  assign n5900 = ~n2075 & (n2955 | (n1723 & n543));
  assign n5901 = (x6 | ~x7 | ~x1 | x2) & (x1 | x7 | (x2 ^ ~x6));
  assign z311 = ~n5907 | (~x3 & (n5903 | n5905 | n5906));
  assign n5903 = ~x1 & ((n530 & n2058) | (~x2 & ~n5904));
  assign n5904 = (~x0 | ~x4 | ~x5 | x6 | ~x7) & (x4 | ((x5 | x6 | ~x7) & (x0 | ~x6 | (~x5 ^ ~x7))));
  assign n5905 = ~n1954 & ((n525 & n813) | (~n573 & ~n643));
  assign n5906 = n543 & ((n1518 & n978) | (x2 & ~n1113));
  assign n5907 = ~n5910 & ~n5912 & (x3 ? n5908 : n5913);
  assign n5908 = (x0 | n5909) & (~n2742 | (~n942 & ~n1383));
  assign n5909 = (~x1 | ~x4 | ~x5 | x6 | x7) & (x4 | ((x5 | ~x6 | ~x7) & (x1 | x6 | (~x5 ^ ~x7))));
  assign n5910 = x0 & ((n2296 & n676) | (n632 & ~n5911));
  assign n5911 = (x5 | x7 | ~x3 | x4) & (x3 | ((x5 | ~x7) & (x4 | ~x5 | x7)));
  assign n5912 = x3 & ~n765 & (~x0 ^ (~x1 & ~x4));
  assign n5913 = (x0 | x1 | ~x5 | x7) & ((x0 & x1) | (x4 ? (x5 | ~x7) : (~x5 | x7)));
  assign z312 = n5920 | ~n5923 | (~x2 & ~n5915);
  assign n5915 = x1 ? n5918 : (~n5917 & (~x0 | n5916));
  assign n5916 = (x3 | ~x5 | (x4 ? (~x6 | ~x7) : (x6 | x7))) & (x5 | (x3 ? (x6 | (~x4 ^ ~x7)) : (~x6 | (x4 ^ ~x7))));
  assign n5917 = n1380 & ((n828 & n1857) | (x6 & ~n671));
  assign n5918 = x6 ? (~n1310 | (~n2648 & ~n5212)) : n5919;
  assign n5919 = x0 ? (x5 | ((x4 | x7) & (x3 | ~x4 | ~x7))) : (~x5 | ((~x4 | ~x7) & (~x3 | x4 | x7)));
  assign n5920 = ~x0 & (n5922 | (~x2 & ~n5921));
  assign n5921 = (x1 | x3 | x4 | x5 | ~x6) & (~x4 | (x1 ? ((~x5 | ~x6) & (~x3 | x5 | x6)) : (x6 | (x3 & ~x5))));
  assign n5922 = x2 & x4 & (x1 ? (x5 ^ ~x6) : (x5 & ~x6));
  assign n5923 = ~n1225 & (~n560 | ~n3217) & (~x2 | n5924);
  assign n5924 = (n814 | ~n4199) & (n671 | n2290 | ~n1686);
  assign z313 = n5929 | n5932 | (x2 ? ~n1237 : ~n5926);
  assign n5926 = ~n1233 & (x3 | n5927);
  assign n5927 = x5 ? n5928 : (~n543 | (~n1479 & ~n3261));
  assign n5928 = ((~x4 ^ ~x6) | (x0 ? (x1 | ~x7) : (~x1 | x7))) & (x1 | x7 | (x0 ? (x4 | ~x6) : (~x4 | x6)));
  assign n5929 = ~x2 & ((x3 & ~n5930) | (n622 & ~n5931));
  assign n5930 = (x0 | ~x1 | (x5 ? (~x6 | x7) : (~x6 ^ ~x7))) & (x1 | ((~x5 | x6 | x7) & (~x0 | (x5 ? ~x6 : (x6 | ~x7)))));
  assign n5931 = (x5 | (x1 ? (x6 | ~x7) : (~x6 ^ ~x7))) & (~x1 | ~x5 | (~x6 & x7));
  assign n5932 = n1181 & ((x5 & ~x6 & x7) | (~x1 & (x5 ? x7 : (x6 & ~x7))));
  assign z314 = ~n5936 | (~x2 & (n5934 | (n699 & n1621)));
  assign n5934 = ~x5 & (x6 ? ~n5935 : (~n1246 & n2553));
  assign n5935 = (~x0 | ~x1 | ~x3 | x4 | x7) & (x0 | x3 | (x1 ? (~x4 | ~x7) : (x4 | x7)));
  assign n5936 = n1249 & (x2 | n1248) & (~n1250 | n5937);
  assign n5937 = (~x6 | ~x7 | ~x1 | x4) & (x6 | x7 | x1 | ~x4);
  assign z315 = n5939 | n5942 | ~n5943 | (n1080 & ~n2460);
  assign n5939 = ~x2 & ((n543 & n5940) | (~x4 & ~n5941));
  assign n5940 = ~x3 & x4 & (x5 ^ ~x7);
  assign n5941 = (x0 | x1 | x3 | x5 | ~x7) & (~x0 | ~x3 | x7 | (~x1 ^ x5));
  assign n5942 = ~x2 & (x0 ? (~x3 & (~x1 ^ ~x7)) : (x3 & (x1 ^ ~x7)));
  assign n5943 = ~n5944 & (n643 | n4317 | x4 | ~n804);
  assign n5944 = x2 & ((~x1 & ~x7) | (~x0 & x1 & x7));
  assign z316 = ~n5949 | ~n5948 | n5946 | n5947;
  assign n5946 = n653 & (n5162 | (x1 & x4 & ~n968));
  assign n5947 = n3517 & ((n1358 & n699) | (n704 & n712));
  assign n5948 = ~n1693 & ~n1270 & ~n3694 & (~n560 | ~n639);
  assign n5949 = (~n1145 | n815 | n4317) & (~n653 | n5950);
  assign n5950 = x1 ? (~x2 | x4) : (x2 | ~x4);
  assign z317 = n3829 | n5954 | ~n5956 | (~x0 & ~n5952);
  assign n5952 = ~n5953 & (~x1 | ~x2 | ~n1716) & (x1 | x2 | n647);
  assign n5953 = x5 & (x1 ? (x2 & ~n752) : (~x2 & n761));
  assign n5954 = x2 & (n5955 | (x4 & n543 & n719));
  assign n5955 = x6 & n1145 & (n4365 | (x0 & n1458));
  assign n5956 = ~n5957 & ~n5958 & n5959 & (~n639 | ~n841);
  assign n5957 = x4 & (x0 ? (~x1 & x3) : (~x5 & (x1 ^ ~x3)));
  assign n5958 = n1614 & x5 & n1167;
  assign n5959 = (~n880 | ~n830) & (~n774 | ~n1723 | ~n560);
  assign z318 = ~n5961 | n5970 | (x6 & (n5966 | n5968));
  assign n5961 = ~n5965 & ~n5964 & n5963 & n3844 & ~n5962;
  assign n5962 = n1084 & ~n1238;
  assign n5963 = ~n570 | (x0 ? ~n926 : ~n1643);
  assign n5964 = n1380 & ((x4 & x6 & x1 & x2) | (~x1 & ((x4 & ~x6) | (~x2 & ~x4 & x6))));
  assign n5965 = n1549 & (x1 ? (~x3 & n1479) : (x3 & ~n1408));
  assign n5966 = ~n671 & ~n5967;
  assign n5967 = (x0 | x1 | ~x2 | ~x3 | ~x5) & (~x0 | x5 | (x1 ? (x2 | x3) : ~x2));
  assign n5968 = n560 & n5969;
  assign n5969 = ~x7 & ~x5 & x3 & x4;
  assign n5970 = n706 & ((n560 & n2765) | (n2940 & ~n5971));
  assign n5971 = (~x3 | x4 | x7) & (~x4 | ~x7);
  assign z319 = n5977 | n5981 | n5984 | (~x3 & ~n5973);
  assign n5973 = x2 ? (~n543 | ~n5974) : (~n5975 & n5976);
  assign n5974 = ~x6 & ~x7 & (x4 ^ x5);
  assign n5975 = n1986 & ((x1 & x6 & (x4 ^ ~x5)) | (~x5 & ~x6 & ~x1 & x4));
  assign n5976 = (~x0 | x1 | x4 | ~x5 | ~x6) & (x0 | ~x1 | x6 | (~x4 ^ ~x5));
  assign n5977 = ~x1 & (~n5979 | (~x7 & ~n5978));
  assign n5978 = (x0 | ~x2 | x3 | ~x5 | ~x6) & (x2 | x6 | (x0 ? (~x3 ^ ~x5) : (~x3 | x5)));
  assign n5979 = n5980 & (~n594 | ~n1070);
  assign n5980 = x0 ? ((~x5 | x6 | ~x7) & (~x2 | (x5 ? x7 : (~x6 | ~x7)))) : (x5 ? (~x6 | (x2 & ~x7)) : (x6 | (~x2 & ~x7)));
  assign n5981 = x1 & (x5 ? ~n5983 : ~n5982);
  assign n5982 = (x0 | ~x2 | ~x3 | x6 | x7) & (~x0 | x2 | x3 | ~x6 | ~x7);
  assign n5983 = (~x0 & ~x2 & ~x3 & (~x6 | ~x7)) | (x0 & (x3 | (x6 & x7))) | (x2 & (x0 | (~x6 & ~x7)));
  assign n5984 = ~n5985 & n569 & n1188;
  assign n5985 = (x0 | ~x2 | ~x4 | x5) & (~x0 | x2 | (~x4 ^ ~x5));
  assign z320 = n5987 | ~n5990 | ~n5992 | (~n643 & ~n5989);
  assign n5987 = n2933 & ~n5988;
  assign n5988 = (~x3 | x5 | x6 | ~x0 | x2) & (x0 | x3 | ~x5 | (~x2 ^ ~x6));
  assign n5989 = ~n1613 & ~n3279 & (~n2940 | (~x3 & ~x4));
  assign n5990 = (~n560 | ~n1141) & (~n2315 | n5991);
  assign n5991 = (x0 | ~x2 | ~x3 | x4 | x5) & (~x0 | x2 | x3 | ~x4 | ~x5);
  assign n5992 = (x0 | n5995) & (n640 | (n5994 & (~x0 | n5993)));
  assign n5993 = x1 ? (x2 | x3) : (~x2 & (~x3 | ~x4));
  assign n5994 = ~n3377 & (~n1167 | (~n1195 & (~n1301 | ~n570)));
  assign n5995 = (x1 & x6) | (~x6 & (~x1 | (~x2 & ~x3 & ~x4))) | (x2 & (x3 | (x4 & ~x6)));
  assign z321 = n6000 | ~n6003 | (x4 ? ~n6002 : ~n5997);
  assign n5997 = ~n5998 & (~n742 | (~n5886 & (~n658 | ~n1317)));
  assign n5998 = ~x2 & ((n942 & n1244) | (x7 & ~n5999));
  assign n5999 = (x0 | ~x1 | x3 | ~x5 | x6) & (~x0 | ~x3 | (x1 ? (x5 | x6) : (~x5 | ~x6)));
  assign n6000 = n1167 & ~n6001;
  assign n6001 = (x1 | ~x2 | ~x3 | (~x5 ^ ~x7)) & (x3 | ((x1 | x2 | ~x5 | x7) & (~x1 | (x2 ? (~x5 ^ ~x7) : (x5 | ~x7)))));
  assign n6002 = (x3 | x7 | x0 | x2) & (~x7 | ((x2 | ~x3 | ~x0 | x1) & (x0 | ~x2 | (~x1 ^ x3))));
  assign n6003 = ~n6004 & ~n6005 & n6006 & (~n895 | ~n4293);
  assign n6004 = x1 & ((~x3 & x7 & x0 & ~x2) | (~x0 & x3 & (x2 ^ ~x7)));
  assign n6005 = ~x1 & (x0 ? (x2 & x7) : (~x7 & (x2 ^ x3)));
  assign n6006 = (~n1241 | ~n2144) & (~n560 | ~n2992);
  assign z322 = ~n6010 | (~x4 & (n6009 | (x5 & ~n6008)));
  assign n6008 = (~x0 | x1 | ~x3 | n785) & (x0 | ~x1 | x3 | n3929);
  assign n6009 = n1723 & ((n626 & n1413) | (n743 & ~n1605));
  assign n6010 = n6013 & (~n774 | n6011) & (x4 | n6012);
  assign n6011 = (~x0 | ~x1 | x2 | x5 | x6) & (x1 | ((~x0 | ~x5 | (~x2 ^ ~x6)) & (x5 | x6 | x0 | ~x2)));
  assign n6012 = (x0 | ~x1 | ~x2 | x3 | x5) & (x1 | x2 | (x0 ? (~x3 ^ x5) : (~x3 | ~x5)));
  assign n6013 = (x1 | ~x2 | (x0 ? (~x3 | ~x4) : x3)) & (x2 | ((~x1 | x3 | ~x4) & ((~x1 & ~x4) | (x0 ^ ~x3))));
  assign z323 = n6015 | n6019 | ~n6023 | (~x4 & ~n6022);
  assign n6015 = ~x1 & (n6016 | (n600 & n1621));
  assign n6016 = ~x4 & ((~x0 & ~n6017) | (n898 & ~n6018));
  assign n6017 = (x2 | x3 | ~x5 | x6 | ~x7) & (~x2 | ~x3 | x5 | ~x6 | x7);
  assign n6018 = (~x2 | ~x3 | ~x5 | x6) & (x2 | ~x6 | (~x3 ^ ~x5));
  assign n6019 = ~x4 & ((~x1 & ~n6020) | (n632 & ~n6021));
  assign n6020 = x0 ? ((~x2 | x3 | ~x5 | ~x6) & (x2 | x6 | (~x3 ^ ~x5))) : ((~x5 | ~x6 | x2 | x3) & (x5 | x6 | ~x2 | ~x3));
  assign n6021 = (x0 | x3 | (~x5 ^ x6)) & (~x3 | (x0 ? (x5 | x6) : (~x5 | ~x6)));
  assign n6022 = (~x0 | ~x1 | x2 | x3 | ~x5) & (x0 | ((x1 | x2 | ~x3 | x5) & (~x2 | (x1 ? (~x3 ^ ~x5) : (x3 | ~x5)))));
  assign n6023 = ~n6025 & n6026 & (~n2933 | n6024);
  assign n6024 = (~x0 | x2 | ~x3 | x5 | ~x6) & (x0 | x3 | ~x5 | (x2 ^ ~x6));
  assign n6025 = ~x0 & x4 & (x1 ^ ~x3);
  assign n6026 = ~n6027 & (~n1716 | ~n841) & (~n560 | ~n1202);
  assign n6027 = x0 & ~x3 & x4 & (~x1 ^ ~x2);
  assign z324 = ~n6037 | (x5 ? ~n6032 : (n6029 | n6030));
  assign n6029 = n837 & n774 & n569;
  assign n6030 = ~x1 & ((n550 & n2435) | (~x3 & ~n6031));
  assign n6031 = (x0 | ~x2 | ~x4 | ~x6 | ~x7) & (x2 | ((x6 | ~x7 | x0 | x4) & (~x0 | ~x6 | (~x4 ^ ~x7))));
  assign n6032 = ~n6036 & (x6 | (~n6034 & (x0 | n6033)));
  assign n6033 = x1 ? ((x2 | ~x3 | ~x4 | ~x7) & (~x2 | x3 | x4 | x7)) : (x2 | x3 | (~x4 ^ ~x7));
  assign n6034 = n841 & ((n1044 & n1379) | (x2 & n6035));
  assign n6035 = x3 & (x4 ^ ~x7);
  assign n6036 = ~n5971 & n841 & n778;
  assign n6037 = ~n6040 & ~n6041 & n6042 & (x2 | n6038);
  assign n6038 = (x4 | n6039) & (~n2024 | (~x1 & x3));
  assign n6039 = (x0 | x1 | x3 | x5 | ~x6) & (x6 | ((~x0 | ~x1 | ~x3 | x5) & ((~x3 ^ ~x5) | (~x0 ^ x1))));
  assign n6040 = ~n1134 & ((~x0 & ((x2 & ~x3) | (~x1 & ~x2 & x3))) | (x1 & (x0 ? (~x2 & ~x3) : x2)));
  assign n6041 = n570 & ((n536 & n559) | (~n1353 & ~n2924));
  assign n6042 = x3 ? n6043 : (~n681 | ~n1209);
  assign n6043 = (x0 | ((x1 | ~x2 | ~x4 | ~x5) & (~x1 | x2 | x4 | x5))) & (x4 | x5 | ~x0 | x1);
  assign z325 = n6050 | ~n6057 | (x2 ? ~n6055 : ~n6045);
  assign n6045 = x0 ? (~n6046 & (x1 | n6047)) : n6048;
  assign n6046 = ~n1353 & ((n750 & n1188) | (n757 & n1317));
  assign n6047 = x3 ? ((~x6 | ~x7 | x4 | x5) & (x6 | x7 | ~x4 | ~x5)) : (x5 | ((~x6 | x7) & (x4 | x6 | ~x7)));
  assign n6048 = (~n689 | ~n658) & (x5 | n6049);
  assign n6049 = (x6 | ~x7 | x3 | x4) & (~x1 | ~x3 | ~x4 | (~x6 ^ x7));
  assign n6050 = ~n1548 & (n6051 | n6052 | ~n6053);
  assign n6051 = ~x5 & (x0 ? (x1 ? (~x2 & ~x6) : (x2 & x6)) : ((~x1 & x2 & ~x6) | (x6 & (x1 | ~x2))));
  assign n6052 = n551 & ((x0 & ~x2 & (x6 ^ x7)) | (x2 & (x0 ? (~x6 & ~x7) : (x6 & x7))));
  assign n6053 = (x2 | ~x5 | x6 | ~n543) & (x5 | n6054);
  assign n6054 = (x0 | x1 | (x2 ? (~x6 | x7) : (x6 | ~x7))) & (~x1 | ((x6 | ~x7 | x0 | ~x2) & (~x0 | x2 | ~x6 | x7)));
  assign n6055 = ~n6056 & (x4 | x5 | ~n841 | n3315);
  assign n6056 = ~n1205 & ((n841 & n1358) | (n1167 & ~n5699));
  assign n6057 = ~n6058 & ~n6061 & ~n6062 & (n2527 | n6060);
  assign n6058 = ~x5 & (x6 ? ~n6059 : (n689 & ~n2185));
  assign n6059 = x0 ? ((x1 | ~x2 | ~x3 | ~x4) & (~x1 | x2 | x3 | x4)) : (~x3 | ~x4 | (~x1 ^ ~x2));
  assign n6060 = (x5 | ((x0 | (x1 & ~x2)) & (x1 | ~x2 | ~x7))) & (x2 | ~x5 | (x0 ? (x1 | ~x7) : (~x1 | x7)));
  assign n6061 = ~n1967 & ~n5422;
  assign n6062 = n4240 & (n6063 | (n1835 & n622));
  assign n6063 = x6 & x4 & ~x0 & x3;
  assign z326 = n6065 | n6070 | ~n6076 | (~x0 & ~n6075);
  assign n6065 = ~x2 & (n6066 | n6068);
  assign n6066 = x0 & ((~x4 & ~n6067) | (~x1 & n2724));
  assign n6067 = (x5 | x7 | ((~x3 | ~x6) & (~x1 | x3 | x6))) & (x1 | (~x6 ^ x7));
  assign n6068 = ~x0 & ((~n640 & ~n5765) | (n1145 & n6069));
  assign n6069 = ~x5 & (x3 ? (~x6 & ~x7) : (x6 & x7));
  assign n6070 = x2 & (n6074 | (~x0 & (n6071 | ~n6072)));
  assign n6071 = ~n643 & ((x3 & (x1 ? (x4 & x5) : (~x4 & ~x5))) | (~x1 & ~x3 & (x4 | x5)));
  assign n6072 = (~n6073 | ~n943) & (~n1317 | (~n2723 & ~n2402));
  assign n6073 = ~x4 & ~x1 & x3;
  assign n6074 = x0 & ~x1 & x3 & (x6 ^ ~x7);
  assign n6075 = (~x3 | x4 | x6 | ~x1 | x2) & (~x2 | ((~x4 | x6 | x1 | ~x3) & (~x1 | ~x6 | (~x3 ^ x4))));
  assign n6076 = ~n6077 & ~n6078 & (~n1723 | ~n742 | n905);
  assign n6077 = ~x3 & ((~x0 & x1 & ~x2 & ~x6) | (x0 & (x1 ? (~x2 & x6) : (x2 & ~x6))));
  assign n6078 = x6 & x3 & ~x2 & ~x0 & ~x1;
  assign z327 = n6080 | ~n6086 | (~x0 & (n6083 | n6085));
  assign n6080 = ~x1 & ((n547 & n830) | (x3 & ~n6081));
  assign n6081 = (~x5 | n6082) & (x4 | x5 | ~n1181 | n640);
  assign n6082 = (x0 | ~x2 | x4 | x6 | x7) & (~x0 | x2 | ~x4 | ~x6 | ~x7);
  assign n6083 = n1145 & (n6084 | (x5 & ~n835));
  assign n6084 = x2 & ~x5 & (x3 ^ x7);
  assign n6085 = x4 & n1133 & (x3 ? (x5 ^ x7) : (x5 & x7));
  assign n6086 = ~n6087 & ~n6090 & (x0 ? n6088 : n6089);
  assign n6087 = n837 & n526 & n828;
  assign n6088 = (x2 | ((x1 | x7) & (~x4 | ~x7 | ~x1 | x3))) & (x1 | ((~x3 | x7) & (~x2 | x3 | ~x7)));
  assign n6089 = (~x4 | ((~x1 | x2 | ~x3 | x7) & (x1 | (~x3 ^ ~x7)))) & (~x1 | (x3 ? (x4 | ~x7) : (x2 ? (x4 | x7) : ~x7)));
  assign n6090 = n1093 & ((~n5194 & n2302) | (n594 & n1395));
  assign z328 = ~n6099 | n6092 | n6094;
  assign n6092 = x2 & ((n727 & n993) | (x7 & ~n6093));
  assign n6093 = (x0 | ~x1 | x4 | ~n1520) & (~x0 | x1 | n4302);
  assign n6094 = ~x2 & (n6095 | (n689 & n1479 & ~n6098));
  assign n6095 = x6 & (x0 ? ~n6097 : ~n6096);
  assign n6096 = (x1 | ~x3 | ~x4 | x5 | ~x7) & (~x1 | x3 | x4 | ~x5 | x7);
  assign n6097 = (x1 | ~x3 | ~x4 | ~x5 | x7) & (~x1 | x5 | (x3 ? (x4 | x7) : (~x4 | ~x7)));
  assign n6098 = x0 ? (~x5 | x7) : (x5 | ~x7);
  assign n6099 = n6101 & ~n6100 & ~n5227 & ~n1120 & ~n5225;
  assign n6100 = n934 & ((n922 & n761) | (n626 & ~n752));
  assign n6101 = ~n6102 & (~n959 | ~n837) & (n1934 | n1119);
  assign n6102 = (x2 ^ ~x5) & (x0 ? (~x1 & x4) : (x1 & ~x4));
  assign z329 = n6112 | ~n6113 | (x0 ? ~n6104 : ~n6108);
  assign n6104 = ~n6105 & ~n6106;
  assign n6105 = x4 & ((~n765 & ~n2499) | (n804 & ~n3925));
  assign n6106 = ~x4 & (x3 ? ~n6107 : (n570 & n881));
  assign n6107 = (~x1 | x2 | x5 | ~x6 | x7) & (x1 | x6 | ~x7 | (~x2 ^ ~x5));
  assign n6108 = x3 ? (~n6109 & (~n702 | n5950)) : n6110;
  assign n6109 = ~x6 & ((n632 & n717) | (n570 & n2317));
  assign n6110 = (x2 | n6111) & (~x1 | ~x2 | x4 | ~n813);
  assign n6111 = x1 ? (~x6 | (x4 ? (x5 | ~x7) : (~x5 | x7))) : (x6 | (x4 ? (x5 | x7) : (~x5 | ~x7)));
  assign n6112 = ~n1548 & (x6 ? ~n5236 : (n632 & ~n791));
  assign n6113 = n6118 & (~n841 | n6114) & (x0 | n6115);
  assign n6114 = (x4 | x5 | x2 | x3) & (~x5 | ((x2 | ~x3 | x4 | x6) & (~x2 | (x3 ? (~x4 | ~x6) : x6))));
  assign n6115 = n6117 & (n623 | n4477) & (~n2371 | n6116);
  assign n6116 = (~x4 | ~x6 | ~x1 | ~x3) & (x1 | x3 | (~x4 ^ x6));
  assign n6117 = (~x1 | ~x2 | ~x3 | x5 | x6) & (x1 | x2 | x3 | ~x5 | ~x6);
  assign n6118 = x5 ? (x6 ? n5235 : n6119) : (x6 ? n6119 : n5235);
  assign n6119 = (~x0 | x1 | x2 | ~x3 | ~x4) & (x0 | ((x1 | ~x2 | ~x3 | ~x4) & (~x1 | x2 | x3 | x4)));
  assign z330 = ~n6135 | ~n6130 | n6128 | n6121 | n6123;
  assign n6121 = ~x3 & ((n662 & n1269) | (~x2 & ~n6122));
  assign n6122 = (~x4 | ~n530 | x0 | ~x1) & (~x0 | (x1 ? (~x4 | ~n813) : (x4 | ~n530)));
  assign n6123 = ~n643 & (~n6125 | (~x2 & ~n6124));
  assign n6124 = (x0 | ~x1 | x3 | x4 | ~x5) & (~x0 | ~x3 | (x1 ? (x4 | x5) : (~x4 | ~x5)));
  assign n6125 = ~n6126 & (n905 | ~n6127) & (~n825 | n5950);
  assign n6126 = ~x3 & ((x1 & ~x2 & x4) | (x0 & ~x1 & x2 & ~x4));
  assign n6127 = ~x5 & ~x0 & x2;
  assign n6128 = n841 & ~n6129;
  assign n6129 = (x2 | ~x3 | ~x4 | x5 | x6) & (x4 | ((~x2 | ~x3 | x5 | ~x6) & (x2 | (x3 ? (~x5 | x6) : (x5 | ~x6)))));
  assign n6130 = ~n6131 & ~n6133 & n6134 & (x3 | n6132);
  assign n6131 = n825 & ((~x4 & x6 & x1 & ~x2) | (~x1 & ~x6 & (x2 ^ ~x4)));
  assign n6132 = (x0 | ~x1 | ~x2 | ~x4 | x6) & (~x0 | ((x1 | ~x2 | ~x4 | ~x6) & (~x1 | x2 | x4 | x6)));
  assign n6133 = ~n905 & n1300 & n1310;
  assign n6134 = (~n610 | ~n712) & (~n588 | ~n2534);
  assign n6135 = (n640 | ~n6139) & (x0 | (n6136 & (n640 | n6138)));
  assign n6136 = (~n559 | ~n2135) & (x3 | n6137);
  assign n6137 = (x1 | ~x4 | (x2 ? (x5 | ~x6) : (~x5 | x6))) & (x4 | ((x1 | ~x2 | ~x5 | ~x6) & (~x1 | x6 | (~x2 ^ ~x5))));
  assign n6138 = x1 ? ((x2 | ~x3 | ~x4 | ~x5) & (~x2 | x3 | x4 | x5)) : (x2 ? (~x3 | x4) : (x3 | (~x4 ^ x5)));
  assign n6139 = n841 & (x2 ? n1909 : n1392);
  assign z331 = n6141 | n6145 | (x2 ? ~n6153 : ~n6149);
  assign n6141 = x0 & (n6142 | (n576 & n931));
  assign n6142 = ~x1 & ((~x2 & ~n6143) | (n885 & ~n6144));
  assign n6143 = (~x3 | ~x4 | ~x5 | ~x6 | x7) & (x4 | (x3 ? (x5 | (~x6 ^ ~x7)) : (~x5 | (~x6 ^ x7))));
  assign n6144 = (x4 | x5 | x6 | ~x7) & (~x4 | ~x5 | (~x6 ^ ~x7));
  assign n6145 = ~x0 & (n6146 | (n3151 & ~n6148));
  assign n6146 = ~x5 & ((~n905 & ~n6147) | (n576 & n1395));
  assign n6147 = x2 ? (~x6 | ~x7) : (x6 ^ ~x7);
  assign n6148 = x1 ? ((x2 | ~x4 | ~x6 | ~x7) & (~x2 | x4 | x6 | x7)) : (~x4 | x7 | (~x2 ^ ~x6));
  assign n6149 = ~n6150 & n6151 & ~n6152 & (n1605 | n4758);
  assign n6150 = ~n714 & ((n841 & n2438) | (~x0 & n683));
  assign n6151 = (~x1 | x3 | ~n674) & (x0 | x1 | ~x3 | ~n4089);
  assign n6152 = (x1 ? (~x4 & x7) : (x4 & ~x7)) & (~x0 ^ ~x3);
  assign n6153 = ~n6154 & (x1 ? (x0 | n3266) : n6155);
  assign n6154 = ~n714 & ((x0 & ~x1 & x3 & ~x7) | (~x0 & ((~x3 & x7) | (x1 & x3 & ~x7))));
  assign n6155 = (~x0 & ~x3 & (x5 | x7)) | (x0 & x3) | (~x4 & x7) | (x4 & ~x7);
  assign z332 = ~n6157 | n6164 | (~x3 & (n6166 | n6168));
  assign n6157 = ~n6158 & (n1198 | n6161) & (~x3 | n6162);
  assign n6158 = ~x1 & (x0 ? ~n6159 : ~n6160);
  assign n6159 = (~x5 | ((x2 | x4 | ~x6) & (~x3 | (~x6 & (~x2 | x4))))) & (x3 | x5 | ((~x4 | x6) & (~x2 | (~x4 & x6))));
  assign n6160 = x3 ? (x5 | (x6 & (x2 | ~x4))) : (~x5 | (x4 ? ~x6 : ~x2));
  assign n6161 = (x0 | ~x2 | ~x3 | (x1 ^ ~x4)) & (x2 | (x0 ? (x1 ? (x3 | ~x4) : (~x3 | x4)) : (x1 ? (~x3 | ~x4) : (x3 | x4))));
  assign n6162 = (~x0 | x1 | ~x7 | n4781) & (x0 | (x1 ? n6163 : (x7 | n4781)));
  assign n6163 = (x2 | x4 | ~x5 | x6 | x7) & (~x2 | ~x4 | x5 | ~x6 | ~x7);
  assign n6164 = x1 & (x0 ? (n1044 & n696) : ~n6165);
  assign n6165 = x4 ? (x3 ? (~x5 | (~x2 & ~x6)) : (x5 | x6)) : ((x2 | (~x3 ^ x5)) & (x3 | ~x5 | ~x6) & (~x3 | x5 | x6));
  assign n6166 = ~x2 & ((~n1850 & ~n2929) | (x6 & ~n6167));
  assign n6167 = (~x4 | x5 | x7 | ~x0 | x1) & (x0 | ~x1 | ~x7 | (~x4 ^ ~x5));
  assign n6168 = x2 & (x0 ? (n772 & n658) : ~n6169);
  assign n6169 = x1 ? ((~x4 | x5 | ~x6 | x7) & (x4 | ~x5 | x6 | ~x7)) : (~x7 | (x4 ? (~x5 | x6) : (x5 | ~x6)));
  assign z333 = ~n6180 | n6176 | n6171 | n6174;
  assign n6171 = ~x2 & (n6172 | (n588 & n1234));
  assign n6172 = ~x3 & ((n529 & n1070) | (x4 & ~n6173));
  assign n6173 = (~x1 | ((x6 | ~x7 | ~x0 | x5) & (x0 | ~x5 | (~x6 ^ ~x7)))) & (~x0 | x1 | x7 | (~x5 ^ ~x6));
  assign n6174 = ~n671 & (x6 ? ~n6175 : (~n2227 & n1411));
  assign n6175 = (~x0 | ~x1 | x2 | x3 | x5) & (x1 | ((~x2 | ~x3 | x5) & (x0 | (x2 ? x5 : (x3 | ~x5)))));
  assign n6176 = ~x0 & (n6178 | ~n6179 | (~x5 & ~n6177));
  assign n6177 = x1 ? ((~x4 | ~x6 | x2 | x3) & (~x2 | x4 | x6)) : (~x3 | (x2 ? (~x4 | x6) : (x4 | ~x6)));
  assign n6178 = ~n2227 & ((n1445 & n1364) | (~x1 & n3795));
  assign n6179 = (n1408 | n2889) & (~n576 | ~n728);
  assign n6180 = ~n6181 & n6185 & (n1353 | n6184);
  assign n6181 = ~n1218 & ((n841 & ~n6182) | (~x0 & ~n6183));
  assign n6182 = (~x2 | x3 | ~x5 | x6) & (x2 | (x3 ? (~x5 | x6) : (x5 | ~x6)));
  assign n6183 = (~x1 | ~x2 | x5 | ~x6) & (x1 | ~x5 | x6 | (x2 & x3));
  assign n6184 = (x1 | ~x2 | ~x3 | ~x5) & (~x1 | x2 | (x0 ? (x3 | ~x5) : (~x3 | x5)));
  assign n6185 = ~n841 | (n6186 & (~n596 | ~n931));
  assign n6186 = ((~x4 ^ ~x5) | (x2 ? (x3 | ~x6) : (~x3 ^ ~x6))) & (x2 | x3 | x4 | ~x5 | ~x6) & (~x4 | x5 | x6 | (~x2 & ~x3));
  assign z334 = n6192 | ~n6195 | (~x5 & (n6188 | n6190));
  assign n6188 = x0 & ((n548 & n1439) | (~x4 & ~n6189));
  assign n6189 = (x1 | ~x2 | x3 | ~x6 | x7) & (x2 | x6 | ((x3 | x7) & (~x1 | ~x3 | ~x7)));
  assign n6190 = ~x0 & ((n558 & n3790) | (x1 & ~n6191));
  assign n6191 = (~x2 | ~x3 | ~x4 | x6 | ~x7) & (x2 | x3 | (x4 ? (~x6 | x7) : ~x7));
  assign n6192 = ~x7 & ((~x0 & ~n6193) | (n841 & ~n6194));
  assign n6193 = (~x2 | (~x5 ^ ~x6)) & (x3 | x5 | (x1 ? x6 : (x2 | ~x6)));
  assign n6194 = (~x2 | (~x5 ^ ~x6)) & (x2 | x3 | ~x5 | x6);
  assign n6195 = n6199 & (~x7 | n6196) & (x2 | n6198);
  assign n6196 = (n710 | n2227 | ~x5 | x6) & (~x6 | (n6197 & (x5 | n710 | n2227)));
  assign n6197 = (~x0 | x1 | ~x2 | ~x3 | x5) & (x0 | ~x1 | (x2 ? (~x3 | x5) : (x3 | ~x5)));
  assign n6198 = x3 ? (x5 | x7 | (x0 & x1)) : ((x0 | x1 | ~x5 | ~x7) & (~x0 | ((x5 | ~x7) & (~x1 | ~x5 | x7))));
  assign n6199 = (~n1269 | ~n2476) & (~n1586 | n6200);
  assign n6200 = x0 ? (x1 | (x4 ? ~x7 : (~x6 | x7))) : (~x1 | (x4 ? (x6 | ~x7) : x7));
  assign z335 = n6206 | ~n6207 | ~n6209 | (~x6 & ~n6202);
  assign n6202 = ~n6205 & (x4 | (~n6204 & (x7 | n6203)));
  assign n6203 = x0 ? ((x1 | ~x2 | ~x3 | ~x5) & (~x1 | x2 | x3 | x5)) : (~x2 | ~x3 | (~x1 ^ ~x5));
  assign n6204 = n619 & ((~x2 & x3 & x5) | (~x0 & (x2 ? (~x3 & ~x5) : x3)));
  assign n6205 = n1029 & ((~x0 & x1 & x2 & ~x7) | (~x1 & ((~x2 & x7) | (x0 & x2 & ~x7))));
  assign n6206 = ~n3309 & ((~x0 & (n3903 | (x1 & n846))) | (~x1 & (n3903 | (x0 & n846))));
  assign n6207 = (n1994 | n6208) & (~n830 | ~n4632);
  assign n6208 = (~x0 | x3 | x4 | x5 | ~x6) & (x0 | ~x3 | x6 | (~x4 & ~x5));
  assign n6209 = (n823 | n6210) & (x3 | (~n6211 & n6212));
  assign n6210 = x2 ? (x6 | (~x3 ^ (x4 | x5))) : (x3 | ~x6);
  assign n6211 = n2332 & ((n922 & n778) | (n626 & n3431));
  assign n6212 = (~x0 | ~x1 | x2 | ~x4 | ~x6) & (x0 | x1 | (x2 ? (~x4 | x6) : ~x6));
  assign z336 = ~n6216 | (n681 & (x7 ? ~n6214 : ~n6215));
  assign n6214 = (~x0 & (~x1 | (~x2 & x6))) | (x0 & x1 & x2) | (~x3 & ~x6) | (x3 & x6);
  assign n6215 = (~x0 | x1 | x2 | x3 | x6) & (x0 | (x3 ? ~x6 : (x6 | (~x1 & ~x2))));
  assign n6216 = n6220 & (x4 ? (n1205 | n710) : n6217);
  assign n6217 = (n1954 | n6218) & (~x5 | n6219);
  assign n6218 = (x0 | ~x3 | ~x5 | x7) & (~x0 | x3 | (~x5 ^ ~x7));
  assign n6219 = (x0 | ~x1 | ~x2 | (~x3 ^ x7)) & (x1 | ((x2 | ~x3 | x7) & (~x0 | ((~x3 | x7) & (x2 | x3 | ~x7)))));
  assign n6220 = (~n626 | ~n2647) & (~n632 | ~n1465 | n1010);
  assign z337 = ~n6223 | (~x2 & (n6222 | (n922 & n959)));
  assign n6222 = ~x5 & ((~n1246 & ~n4910) | (n550 & n712));
  assign n6223 = n6226 & (~x4 | n6224) & (n1954 | n6225);
  assign n6224 = (~x2 | ((~x0 | x1 | ~x5) & (x0 | ~x1 | x5 | ~x6))) & (x0 | x1 | x2 | (~x5 & ~x6));
  assign n6225 = (x0 | ~x4 | (~x5 & ~x6)) & (x4 | x5 | ((x6 | x7) & (~x0 | (x6 & x7))));
  assign n6226 = (n4226 | ~n6227) & (n1957 | (~n1121 & ~n696));
  assign n6227 = x7 & ~x5 & ~x1 & x4;
  assign z338 = ~n6233 | (~x2 & (~n6229 | (~x3 & ~n6232)));
  assign n6229 = (x3 | n6230) & (~n922 | ~n779 | ~x3 | x4);
  assign n6230 = x0 ? (~n1145 | ~n978) : (x6 | n6231);
  assign n6231 = (x5 | x7 | x1 | ~x4) & (~x1 | ~x7 | (x4 ^ ~x5));
  assign n6232 = (~x0 | x1 | ~x5 | ~x6 | ~x7) & (x0 | x6 | (x1 ? (x5 | x7) : (~x5 | ~x7)));
  assign n6233 = n6236 & (n1794 | ~n6234) & (n765 | n6235);
  assign n6234 = ~x6 & ~x5 & x1 & ~x2;
  assign n6235 = (~x0 | ~x1 | x2 | x3 | ~x6) & (x1 | (~x2 & ~x3) | (~x0 ^ ~x6));
  assign n6236 = (x5 | x6 | ~x0 | x1) & (x0 | ((~x5 | ~x6) & (x5 | x6 | ~x1 | ~x2)));
  assign z341 = ~x2 & (n6239 | ~n6240 | (~x1 & ~n6238));
  assign n6238 = x3 ? ((x4 & (~x0 | (x5 & x6))) | (~x0 & (x5 | x6))) : ((x0 & (~x5 | ~x6)) | (~x4 & (x0 | (~x5 & ~x6))));
  assign n6239 = n543 & ((n1029 & n813) | (n530 & n828));
  assign n6240 = (x1 | n573 | n871) & (x0 | ~x1 | n1548);
  assign z342 = n6242 | n6246 | ~n6247 | (~x0 & ~n6245);
  assign n6242 = x3 & (n6243 | (n1291 & ~n5214));
  assign n6243 = ~x1 & (x0 ? n6244 : (n1070 & n1084));
  assign n6244 = x4 & ((~x6 & ~x7 & x2 & ~x5) | (x6 & x7 & ~x2 & x5));
  assign n6245 = (~x1 | x2 | ~x3 | ~x4 | ~x5) & (x1 | ((~x2 | x3 | ~x4 | x5) & (x2 | ~x3 | x4 | ~x5)));
  assign n6246 = x2 & ((~x0 & x1 & ~x3) | (~x1 & ((~x3 & ~x4) | (x0 & (~x3 | ~x4)))));
  assign n6247 = ~n2330 & (~n5433 | n1977) & (~n610 | ~n5198);
  assign z343 = n6253 | ~n6255 | (x7 & (n6249 | n6252));
  assign n6249 = ~x1 & ((x4 & ~n6250) | (~x0 & n6251));
  assign n6250 = (~x0 | x2 | ~x3 | ~x5 | ~x6) & (x6 | ((x0 | ~x2 | x3 | ~x5) & (~x0 | (x2 ? (~x3 | x5) : (x3 | ~x5)))));
  assign n6251 = ~x2 & ~x4 & ~x5 & (x3 ^ ~x6);
  assign n6252 = n543 & ((n704 & n885) | (~x2 & ~n4302));
  assign n6253 = ~x0 & (x1 ? ~n3424 : ~n6254);
  assign n6254 = x2 ? (~x4 | (x3 ? (x5 | x6) : (~x5 | ~x6))) : (x3 | x4 | (~x5 ^ x6));
  assign n6255 = ~n6260 & ~n6259 & ~n6258 & ~n5363 & ~n6256;
  assign n6256 = x0 & ((n576 & n728) | (~x1 & ~n6257));
  assign n6257 = (~x2 | ~x3 | ~x4 | x5 | ~x6) & (x2 | ((x3 | ~x4 | ~x5 | ~x6) & (~x3 | x4 | x5 | x6)));
  assign n6258 = ~n877 & (x0 ? (~x1 & n859) : (x1 & ~n1532));
  assign n6259 = ~x0 & x3 & (x1 ? (x2 & x4) : (x2 ^ x4));
  assign n6260 = n1084 & ((n1451 & n922) | (n1301 & n626));
  assign z344 = n6262 | n6264 | ~n6271 | (~x2 & ~n6267);
  assign n6262 = x0 & ((n576 & n577) | (~x1 & ~n6263));
  assign n6263 = (x3 | x4 | ~x5 | x6) & (~x3 | x5 | (x2 ? (~x4 ^ ~x6) : (x4 | ~x6)));
  assign n6264 = x2 & (n6265 | (~x0 & x1 & ~n4164));
  assign n6265 = ~x1 & ((n943 & n1074) | (n876 & ~n6266));
  assign n6266 = (x4 | ~x6 | x7) & (~x0 | ~x4 | x6 | ~x7);
  assign n6267 = ~n6268 & (~x3 | (~n6269 & (~n529 | ~n942)));
  assign n6268 = ~n5129 & ((n757 & n825) | (n750 & n622));
  assign n6269 = n772 & (n6270 | (x0 & ~n2063));
  assign n6270 = ~x7 & ~x6 & ~x0 & ~x5;
  assign n6271 = (x0 & n6272) | (~n6274 & n6275 & ~x0 & n6273);
  assign n6272 = (x2 | ((x4 | ~x5 | x1 | ~x3) & (~x1 | x3 | ~x4 | x5))) & (x1 | ((x3 | x4 | x5) & (~x2 | ~x4 | ~x5)));
  assign n6273 = ((~x1 ^ ~x2) | (x3 ? (x4 | ~x5) : (~x4 | x5))) & (~x4 | ~x5 | ~x1 | x2) & (x1 | ~x2 | (x3 ? (~x4 | ~x5) : (x4 | x5)));
  assign n6274 = ~n1353 & (x1 ? (~x2 & n876) : (x2 & ~n1566));
  assign n6275 = x1 ? ~n6276 : (~n1044 | ~n577);
  assign n6276 = x2 & ((x5 & x6 & ~x3 & ~x4) | (~x5 & ~x6 & x3 & x4));
  assign z345 = n6287 | n6288 | (x3 ? ~n6278 : ~n6281);
  assign n6278 = n6280 & (~x7 | (~n1208 & (x2 | n6279)));
  assign n6279 = (~x0 | x1 | ~x4 | ~x5 | ~x6) & (x5 | ((x1 | ~x4 | x6) & (x0 | ((~x4 | x6) & (~x1 | x4 | ~x6)))));
  assign n6280 = (x1 | ~x2 | n990) & (x0 | ((~x2 | n990) & (x1 | (n990 & (~x2 | ~n2758)))));
  assign n6281 = ~n6282 & n6286 & (n1408 | n6285);
  assign n6282 = ~x2 & (x6 ? ~n6283 : (n1310 & ~n6284));
  assign n6283 = (x0 | ~x1 | x4 | ~x5 | ~x7) & (x7 | ((~x4 | ~x5 | x0 | ~x1) & (~x0 | x1 | (~x4 ^ ~x5))));
  assign n6284 = x1 ? (~x4 | x7) : (x4 | ~x7);
  assign n6285 = (x0 | ~x1 | ~x2 | x5 | x7) & (x1 | ((~x0 | (x2 ? (x5 | x7) : (~x5 | ~x7))) & (x5 | x7 | x0 | x2)));
  assign n6286 = (~n746 & n4040) | (~n1621 & (~n830 | n4040));
  assign n6287 = x3 & ((~n710 & ~n1100) | (n704 & n560));
  assign n6288 = ~x3 & (n6290 | ~n6291 | (~x2 & ~n6289));
  assign n6289 = (x0 | ~x5 | (x1 ? (~x4 | x6) : (x4 | ~x6))) & (x5 | x6 | ~x0 | x1);
  assign n6290 = ~n1097 & (~n4040 | (x2 & ~x4 & ~n823));
  assign n6291 = ~n3915 & ~n6292 & (~n559 | ~n746);
  assign n6292 = ~x0 & ~x2 & (x1 ? (~x4 & ~x5) : (x4 & x5));
  assign z346 = ~n6303 | (x0 ? ~n6294 : ~n6298);
  assign n6294 = (~x4 | n6295) & (x1 | x4 | n6297);
  assign n6295 = (x6 | ~x7 | ~n1467 | n2737) & (~x6 | n6296);
  assign n6296 = (x2 | (x1 ? (x3 | x7) : (~x5 | ~x7))) & (x1 | x5 | x7 | (~x2 & ~x3));
  assign n6297 = (x2 | ~x5 | ~x6 | (x3 ^ ~x7)) & (x5 | ((~x3 | x6 | x7) & (~x2 | ((x6 | x7) & (x3 | ~x6 | ~x7)))));
  assign n6298 = x2 ? n6301 : (x1 ? n6299 : n6300);
  assign n6299 = (x3 | ~x5 | (x4 ? (~x6 | ~x7) : (x6 | x7))) & (x5 | ((~x3 | x4 | (~x6 ^ ~x7)) & (~x4 | (~x6 ^ x7))));
  assign n6300 = x6 ? (x4 ? (x5 | x7) : ((x5 | ~x7) & (x3 | ~x5 | x7))) : ((~x4 | x5 | ~x7) & (~x3 | (x4 ? ~x7 : (x5 | x7))));
  assign n6301 = x7 ? n6302 : (~n846 & (~n597 | n4493));
  assign n6302 = (~x4 | x5 | x6 | ~x1 | x3) & (x1 | ~x3 | x4 | ~x5 | ~x6);
  assign n6303 = ~n6304 & ~n6308 & n6310 & (~n772 | n6307);
  assign n6304 = ~x4 & ((~x2 & ~n6305) | (n742 & ~n6306));
  assign n6305 = x0 ? ((~x1 | x3 | ~x5 | ~x6) & (x1 | x5 | (~x3 ^ ~x6))) : ((~x3 | ~x5 | ~x6) & (~x1 | x3 | x5 | x6));
  assign n6306 = (~x3 | x5 | x6) & (x1 | x3 | ~x5 | ~x6);
  assign n6307 = (x0 | x2 | x3 | ~x5 | x6) & (~x0 | ((~x2 | x3 | ~x5 | x6) & (x2 | (x3 ? (~x5 | x6) : (x5 | ~x6)))));
  assign n6308 = ~n6309 & (n1621 | (~x4 & ~n1701));
  assign n6309 = (~x0 | x2 | x3) & (~x2 | (x0 & (x1 | ~x3)));
  assign n6310 = x4 ? (~n706 | ~n733) : n6311;
  assign n6311 = (x0 | ~x1 | ~x2 | ~x5 | ~x6) & (~x0 | ((x1 | ~x2 | ~x5 | ~x6) & (~x1 | x2 | x5 | x6)));
  assign z347 = n6317 | ~n6323 | (x0 ? ~n6320 : ~n6313);
  assign n6313 = x1 ? (~n6316 & (~n949 | ~n951)) : n6314;
  assign n6314 = (~x2 | x4 | ~x7 | n3349) & (~x4 | n6315);
  assign n6315 = (x2 | ~x3 | ~x5 | ~x6 | x7) & (~x7 | ((x5 | x6 | x2 | x3) & (~x2 | ((x5 | ~x6) & (x3 | ~x5 | x6)))));
  assign n6316 = x2 & ((~x7 & ~n4302) | (x3 & x7 & ~n1198));
  assign n6317 = ~n1097 & ((n572 & ~n6319) | (~x7 & ~n6318));
  assign n6318 = x0 ? ((x1 | ~x2 | ~x3) & (~x1 | x2 | x3 | x4)) : (~x2 | ((x3 | (x1 & ~x4)) & (~x1 | ~x3 | x4)));
  assign n6319 = x0 ? (x1 | ~x3) : (x3 | (~x1 ^ ~x4));
  assign n6320 = x1 ? ~n6321 : (~n6322 & (~x3 | n3656));
  assign n6321 = ~x2 & ~x3 & x7 & (x5 ^ x6);
  assign n6322 = x7 & n1044 & (x4 ? (x5 & x6) : (~x5 ^ ~x6));
  assign n6323 = ~n6324 & ~n6327 & n6329 & (x1 | n6326);
  assign n6324 = x7 & ((n543 & n2775) | (n570 & ~n6325));
  assign n6325 = x3 ? (~x4 | (x0 ^ ~x5)) : (x4 | x5);
  assign n6326 = (~x0 | x3 | x7 | (~x2 ^ ~x5)) & (~x3 | ((~x0 | x2 | ~x5 | x7) & (x0 | x5 | (x2 ^ ~x7))));
  assign n6327 = ~n6328 & ~x7 & n1181;
  assign n6328 = (~x1 | (x3 ? (~x4 | ~x5) : (x4 | x5))) & (x1 | x3 | x4 | ~x5);
  assign n6329 = (~n746 | ~n1460) & (n1548 | n6330);
  assign n6330 = (~x0 | x5 | (x1 ? (x2 | x7) : (~x2 | ~x7))) & (x0 | x2 | ~x5 | x7);
  assign z348 = ~n6340 | (x1 ? (n2581 | n6332) : ~n6335);
  assign n6332 = ~x0 & ((~x4 & ~n6333) | (n1379 & ~n6334));
  assign n6333 = (x2 | ~x3 | x5 | ~x6 | ~x7) & (x3 | ((~x6 | ~x7 | x2 | ~x5) & (~x2 | x7 | (~x5 ^ ~x6))));
  assign n6334 = (x2 | x3 | ~x5 | x6) & (~x2 | ~x3 | (~x5 ^ x6));
  assign n6335 = x5 ? n6338 : (x4 ? n6337 : n6336);
  assign n6336 = (x0 | ~x2 | x3 | x6 | ~x7) & (~x0 | x2 | ~x3 | ~x6 | x7);
  assign n6337 = (x0 | x2 | ~x3 | x6 | x7) & (~x7 | (~x2 ^ ~x3) | (x0 ^ ~x6));
  assign n6338 = (~n1786 | ~n2435) & (x3 | n6339);
  assign n6339 = (x0 | x4 | (x2 ? (~x6 | ~x7) : (x6 | x7))) & (~x4 | ((x0 | x2 | x6 | ~x7) & (~x0 | ~x6 | (x2 & x7))));
  assign n6340 = x2 ? n6343 : (x7 ? n6342 : n6341);
  assign n6341 = x6 ? ((x0 | x1 | ~x3 | ~x4) & (x3 | x4 | ~x0 | ~x1)) : ((x0 | ((~x3 | x4) & (~x1 | (~x3 & x4)))) & (x1 | x3 | ~x4) & (~x0 | ((x3 | ~x4) & (x1 | (x3 & ~x4)))));
  assign n6342 = (~x6 | ((x3 | (~x1 ^ ~x4)) & (~x0 | (x3 ? x1 : x4)))) & (x0 | x6 | ((~x1 | x3 | x4) & (~x3 | (x1 & ~x4))));
  assign n6343 = n6346 & (~n2320 | ~n6344) & (x1 | n6345);
  assign n6344 = ~x7 & (x3 ^ x4);
  assign n6345 = (x0 | x3 | ~x4 | ~x6 | ~x7) & (~x3 | ((x6 | x7 | x0 | ~x4) & (~x7 | (x0 ? (~x4 ^ ~x6) : (x4 | ~x6)))));
  assign n6346 = (x0 | ~x1 | ~x7 | (~x3 ^ ~x6)) & (x1 | ((x0 | x3 | ~x6 | x7) & (~x0 | (x3 ? (~x6 | x7) : x6))));
  assign z349 = ~n6349 | ~n6353 | ~n6356 | (~x0 & ~n6348);
  assign n6348 = x1 ? (x2 ? (x3 ? (x4 | x7) : (~x4 | ~x7)) : (x7 | (~x3 ^ ~x4))) : ((~x2 | x3 | ~x4 | x7) & (x2 | (x3 ? (~x4 ^ ~x7) : (x4 | ~x7))));
  assign n6349 = (n981 | n6350) & (n6351 | ~n6352);
  assign n6350 = (x0 | x1 | ~x2 | x4 | x7) & (~x0 | ~x7 | (x1 ? (x2 | x4) : (~x2 | ~x4)));
  assign n6351 = x2 ? ((x5 | ~x6 | ~x3 | ~x4) & (x3 | (x4 ? (~x5 | x6) : (x5 | ~x6)))) : ((~x3 | x4 | ~x5 | x6) & (x3 | ~x4 | x5 | ~x6));
  assign n6352 = ~x7 & x0 & ~x1;
  assign n6353 = x0 ? n6354 : (~x1 | n6355);
  assign n6354 = (x1 | ~x2 | ~x3 | x4 | ~x7) & (x2 | ((~x4 | ~x7 | x1 | ~x3) & (x3 | (x1 ? (~x4 ^ ~x7) : (x4 | ~x7)))));
  assign n6355 = (~x7 | ((x4 | x5 | x2 | ~x3) & (~x5 | (x2 ? (~x3 ^ ~x4) : (x3 | ~x4))))) & (~x2 | x5 | x7 | (~x3 ^ ~x4));
  assign n6356 = ~n6357 & (x0 | (~n6360 & (~n4089 | n6363)));
  assign n6357 = ~x1 & (x3 ? ~n6359 : ~n6358);
  assign n6358 = x2 ? ((x5 | ~x7 | x0 | x4) & (~x0 | x7 | (~x4 ^ x5))) : (~x4 | ((~x5 | x7) & (x0 | x5 | ~x7)));
  assign n6359 = (~x0 | x2 | x4 | (~x5 ^ ~x7)) & (~x2 | ((~x0 | ~x4 | ~x5 | x7) & (x0 | ~x7 | (~x4 ^ x5))));
  assign n6360 = x4 & ((n570 & n6361) | (n934 & ~n6362));
  assign n6361 = x3 & x5 & (x6 ^ x7);
  assign n6362 = (x6 | x7 | x1 | ~x3) & (~x1 | x3 | (~x6 ^ ~x7));
  assign n6363 = (~x1 | ((x2 | ~x3 | ~x5 | x6) & (~x2 | x3 | x5 | ~x6))) & (x1 | ~x2 | ~x3 | x5 | ~x6);
  assign z350 = ~n6370 | (~x4 & ~n6365) | (n543 & ~n6369);
  assign n6365 = x7 ? (x2 | n6368) : (~n6366 & n6367);
  assign n6366 = n922 & ~n1566 & ~x2 & x6;
  assign n6367 = (~n1519 | ~n1269) & (n800 | n1916);
  assign n6368 = (x0 | x1 | ~x3 | x5 | ~x6) & (x3 | ((~x0 | x5 | (x1 ^ ~x6)) & (x0 | ~x1 | ~x5 | x6)));
  assign n6369 = x4 ? ((~x2 | (~x3 ^ x5)) & (x2 | x3 | x5 | x6)) : ((~x2 | ~x3 | ~x5 | ~x6) & (x2 | (x3 ? x5 : (~x5 | ~x6))));
  assign n6370 = n6377 & (x1 | n6371) & (~n1518 | n6375);
  assign n6371 = ~n6372 & ~n6373 & ~n6374 & (n1794 | n2760);
  assign n6372 = ~x6 & x5 & x4 & x2 & ~x3;
  assign n6373 = ~x5 & ~x4 & x3 & x0 & ~x2;
  assign n6374 = (x2 ^ x4) & (x0 ? (x3 & x5) : (~x3 & ~x5));
  assign n6375 = x6 ? (~n1188 | ~n6376) : (n1794 | n5786);
  assign n6376 = x7 & (x0 ^ x5);
  assign n6377 = (n1353 | n6378) & (n627 | n6379);
  assign n6378 = (x3 | ~x5 | ~x0 | x2) & (x0 | ((x1 | ~x2 | ~x3 | x5) & (~x1 | (x2 ? (x3 | x5) : (~x3 | ~x5)))));
  assign n6379 = x0 ? (x5 | (x1 ? (x2 | x4) : (~x2 | ~x4))) : (x1 | ~x5 | (~x2 ^ ~x4));
  assign z351 = n6395 | n6392 | ~n6388 | n6381 | n6385;
  assign n6381 = ~x3 & ((~x1 & ~n6382) | (n543 & ~n6384));
  assign n6382 = x2 ? (n3098 | (x0 ^ ~x5)) : (x5 | n6383);
  assign n6383 = (x0 | x4 | ~x6 | ~x7) & (~x0 | x7 | (x4 ^ ~x6));
  assign n6384 = (x2 | ~x4 | ~x5 | x6 | ~x7) & (x4 | ((~x2 | x5 | ~x6 | x7) & (x2 | ~x5 | (~x6 ^ ~x7))));
  assign n6385 = x2 & ((~n1097 & ~n6386) | (~x1 & ~n6387));
  assign n6386 = (~x3 | ~x4 | ~x0 | x1) & (x0 | (x1 ? x3 : (~x3 | x4)));
  assign n6387 = x3 ? ((~x5 | x6 | x0 | ~x4) & (x5 | ~x6 | ~x0 | x4)) : (x0 ? (~x5 | (x4 & x6)) : (x5 | (~x4 & ~x6)));
  assign n6388 = ~n4679 & (n6389 | n6390) & (n1097 | n6391);
  assign n6389 = x0 ? (x2 | x7) : (~x2 | ~x7);
  assign n6390 = x1 ? ((x3 | ~x4 | ~x5 | x6) & (~x3 | x4 | x5 | ~x6)) : (~x3 | (x4 ? (x5 | ~x6) : (~x5 | x6)));
  assign n6391 = (~x0 | x4 | n3827) & (~x4 | n1205 | ~n3828);
  assign n6392 = ~x2 & ((~x0 & ~n4438) | n6393 | (x0 & ~n6394));
  assign n6393 = ~n1097 & ((~x0 & x1 & ~x3 & x4) | (~x1 & (x0 ? (x3 ^ ~x4) : (x3 & ~x4))));
  assign n6394 = (~x1 | ~x3 | x4 | x5 | x6) & (x1 | ((x3 | ~x4 | ~x5 | x6) & (~x3 | x4 | x5 | ~x6)));
  assign n6395 = n825 & (x1 ? ~n6396 : (n942 & n1084));
  assign n6396 = (~x2 | ~x4 | x5 | x6 | ~x7) & (x2 | ~x5 | x7 | (~x4 ^ x6));
  assign z352 = n6406 | ~n6411 | (x1 ? ~n6403 : ~n6398);
  assign n6398 = ~n6401 & (~x7 | (~n6400 & (~x2 | n6399)));
  assign n6399 = x0 ? ((~x5 | ~x6 | x3 | x4) & (x5 | x6 | ~x3 | ~x4)) : (x4 ? (x3 ? (~x5 | x6) : (x5 | ~x6)) : (x5 | x6));
  assign n6400 = n878 & (x0 ? (x3 ? (~x4 & ~x5) : x5) : (~x4 & x5));
  assign n6401 = n1986 & ~n6402;
  assign n6402 = (~x4 | x5 | ~x6 | (~x2 & ~x3)) & (x2 | ~x5 | ((~x4 | ~x6) & (x3 | x4 | x6)));
  assign n6403 = ~n3926 & (x0 | (~x3 & n6404) | (x3 & n6405));
  assign n6404 = (x6 | ~x7 | x2 | x5) & (~x5 | (x2 ? (x4 ? (~x6 | x7) : (x6 | ~x7)) : (x4 | x7)));
  assign n6405 = (x2 | x4 | x5 | ~x6 | ~x7) & (~x2 | ~x5 | (x4 ? ~x6 : (x6 | ~x7)));
  assign n6406 = ~n640 & (n6408 | ~n6409 | (~x1 & ~n6407));
  assign n6407 = (x0 | ~x2 | x3 | x4 | ~x5) & (x2 | ((x3 | ((~x4 | x5) & (~x0 | x4 | ~x5))) & (x0 | ((~x3 | x4 | ~x5) & (~x4 | x5)))));
  assign n6408 = ~n1134 & ((x0 & ~x1 & x2) | (x1 & ~x2 & ~x3));
  assign n6409 = ~n914 & ~n6410 & (~n746 | ~n1641);
  assign n6410 = ~x0 & ((~x1 & x2 & x3 & ~x4) | (x1 & x4 & (x2 ^ x3)));
  assign n6411 = ~n6414 & (n643 | (~n6413 & (x4 | n6412)));
  assign n6412 = (x0 | ~x1 | ~x2 | ~x3 | x5) & (x2 | ((x0 | (x1 ? (~x3 | ~x5) : x5)) & (x3 | ((x1 | x5) & (~x0 | ~x1 | ~x5)))));
  assign n6413 = n772 & ((~x0 & x2 & ~x3 & x5) | (x0 & ~x5 & (~x2 ^ ~x3)));
  assign n6414 = ~n1850 & (n3463 | (~n2227 & ~n3394));
  assign z353 = ~n6421 | ~n6427 | (~x2 & ~n6416);
  assign n6416 = x5 ? n6419 : (x0 ? n6417 : n6418);
  assign n6417 = x1 ? (x6 | (x3 ? (x4 | ~x7) : (~x4 | x7))) : (~x6 | (x3 ^ ~x7));
  assign n6418 = (~x1 | x3 | x4 | x6 | ~x7) & (~x6 | ((x3 | x4 | x7) & (x1 | ~x7 | (~x3 & ~x4))));
  assign n6419 = (~n699 | ~n1786) & (x1 | n6420);
  assign n6420 = (~x7 | (x0 ? (x3 | (~x4 ^ ~x6)) : (x6 | (~x3 & ~x4)))) & (~x3 | x7 | (x0 ? x6 : (x4 | ~x6)));
  assign n6421 = x1 ? n6424 : (x0 ? n6422 : n6423);
  assign n6422 = (~x2 | x4 | (x3 ? (x5 | x7) : (~x5 | ~x7))) & (x3 | ~x4 | x5 | x7) & (x2 | ((x3 | x5 | x7) & (~x5 | ~x7 | ~x3 | ~x4)));
  assign n6423 = (x7 | (x3 ^ ~x4) | (x2 ^ x5)) & (x3 | ~x7 | (x2 ? x5 : (x4 | ~x5)));
  assign n6424 = n6426 & (x2 | n6425);
  assign n6425 = (~x0 | x3 | ~x4 | ~x5 | x7) & (x0 | x5 | ~x7 | (x3 ^ ~x4));
  assign n6426 = (~x0 | x2 | x3 | x5 | ~x7) & (x0 | ~x3 | ~x5 | (~x2 ^ ~x7));
  assign n6427 = ~n6428 & (~x2 | (~n6431 & ~n6432));
  assign n6428 = ~n1097 & (x1 ? ~n6430 : ~n6429);
  assign n6429 = (x0 | ~x2 | x3 | x4 | x7) & (~x3 | (x0 ? (x2 ? (~x4 | x7) : (x4 | ~x7)) : (x2 ? ~x7 : (~x4 | x7))));
  assign n6430 = (~x0 | x2 | x3 | x4 | x7) & (x0 | (x2 ? (x3 | ~x7) : (~x4 | (~x3 ^ ~x7))));
  assign n6431 = ~n1198 & ((n841 & n2492) | (~n1548 & ~n3134));
  assign n6432 = ~x7 & ((~x1 & ~n6434) | (~x0 & x1 & ~n6433));
  assign n6433 = (x3 | x4 | ~x5 | x6) & (~x3 | ~x4 | x5 | ~x6);
  assign n6434 = (x0 | ~x3 | ~x4 | ~x5 | x6) & (~x0 | x4 | ~x6 | (~x3 ^ ~x5));
  assign z354 = ~n6440 | (~x2 & (x0 ? ~n6436 : ~n6438));
  assign n6436 = (x5 | x7 | n6437) & (~x5 | ~x7 | ~n1145 | n1026);
  assign n6437 = (~x1 | (x3 ? (x4 | ~x6) : (~x4 | x6))) & (x1 | x3 | ~x4 | ~x6);
  assign n6438 = x5 ? n6439 : (~n569 | ~n6073);
  assign n6439 = (x1 | ~x3 | x4 | x6 | x7) & (~x7 | (x1 ? (x3 ? (~x4 | x6) : (x4 | ~x6)) : (~x4 | (~x3 ^ ~x6))));
  assign n6440 = ~n6441 & ~n6443 & n6447 & (n640 | n6446);
  assign n6441 = ~x0 & (x1 ? ~n3284 : ~n6442);
  assign n6442 = (x2 | x3 | ~x4 | ~x6 | x7) & (~x3 | ((x6 | ~x7 | x2 | x4) & (~x2 | (x4 ? (x6 | ~x7) : (~x6 | x7)))));
  assign n6443 = x2 & ((~n3266 & ~n6444) | (n825 & ~n6445));
  assign n6444 = (x0 | ~x1 | x3 | ~x6) & (~x0 | x1 | (~x3 ^ ~x6));
  assign n6445 = (~x1 | ~x4 | x5 | x6 | x7) & (x1 | ((~x4 | x5 | ~x6 | x7) & (x4 | ~x5 | x6 | ~x7)));
  assign n6446 = (x2 | ((~x0 | (x1 ? (x3 | x4) : (~x3 | ~x4))) & (x0 | ~x1 | x3 | ~x4))) & (x0 | ~x2 | x4 | (~x1 ^ ~x3));
  assign n6447 = (~x1 | n6450) & (~n841 | n6448) & (x1 | n6449);
  assign n6448 = x2 ? ((x3 | ~x4 | ~x6 | x7) & (~x3 | x4 | x6 | ~x7)) : (x3 | (x4 ? (x6 | ~x7) : (~x6 | x7)));
  assign n6449 = (~x3 | x4 | x6 | ~x0 | x2) & (x0 | ~x2 | x3 | ~x4 | ~x6) & ((~x0 ^ ~x2) | (x3 ? (~x4 | x6) : (x4 | ~x6)));
  assign n6450 = (~x0 | x2 | x3 | ~x4 | ~x6) & (x0 | (~x3 ^ ~x6) | (~x2 ^ ~x4));
  assign z355 = ~n6461 | n6458 | n6452 | n6455;
  assign n6452 = x1 & ((n1693 & n931) | (~x6 & ~n6453));
  assign n6453 = x2 ? (x0 | (~n5969 & ~n4414)) : n6454;
  assign n6454 = (x0 | x3 | x4 | ~x5 | ~x7) & (x5 | ((x0 | ~x3 | ~x4 | ~x7) & (~x0 | (x3 ? (x4 | ~x7) : (~x4 | x7)))));
  assign n6455 = ~x1 & (n6457 | (~n877 & ~n6456));
  assign n6456 = (~x0 | ~x2 | x6 | (~x4 ^ ~x7)) & (x2 | ((x6 | ~x7 | ~x0 | x4) & (x0 | ~x4 | (~x6 ^ x7))));
  assign n6457 = ~x6 & ((n674 & n600) | (~n524 & n1988));
  assign n6458 = ~x0 & (x2 ? ~n6460 : ~n6459);
  assign n6459 = x1 ? ((~x3 | ~x4 | ~x5 | x7) & (x5 | ~x7 | x3 | x4)) : ((~x4 | (x3 ? (x5 | ~x7) : (~x5 | x7))) & (~x3 | x4 | (~x5 ^ ~x7)));
  assign n6460 = (x1 | ~x3 | x4 | ~x5 | x7) & (~x1 | x3 | ~x4 | x5 | ~x7) & ((x1 ? (x3 | x4) : (~x3 | ~x4)) | (~x5 ^ ~x7));
  assign n6461 = n6462 & (~n841 | n6464) & (x1 | n6463);
  assign n6462 = (n1218 | n4075) & (x2 | ~n543 | n3972);
  assign n6463 = (x0 | x2 | x3 | x4 | ~x7) & (~x0 | ((x2 | ~x3 | ~x4 | x7) & (~x2 | x3 | x4 | ~x7)));
  assign n6464 = ((x2 ? (~x3 | x4) : (x3 | ~x4)) | (~x5 ^ ~x7)) & ((x3 ? (x5 | ~x7) : (~x5 | x7)) | (x2 ^ x4));
  assign z356 = ~n6483 | n6479 | n6476 | n6466 | n6473;
  assign n6466 = x1 & (n6471 | (~x2 & (n6467 | n6469)));
  assign n6467 = ~x5 & ~n6468;
  assign n6468 = (~x0 | x7 | (x3 ? (x4 | ~x6) : (~x4 | x6))) & (x0 | x3 | ~x4 | ~x6 | ~x7);
  assign n6469 = n1380 & (n3684 | (x3 & n6470));
  assign n6470 = x7 & (x4 ^ ~x6);
  assign n6471 = ~n6472 & ~x7 & n742;
  assign n6472 = (x5 | x6 | ~x3 | ~x4) & (x3 | ~x5 | (~x4 ^ ~x6));
  assign n6473 = x2 & ((~x1 & ~n6474) | (n3488 & ~n6475));
  assign n6474 = x0 ? ((~x5 | ~x6 | x3 | x4) & (x6 | (x3 ? (~x4 ^ ~x5) : (~x4 | x5)))) : ((x3 | x4 | ~x5 | x6) & (x5 | ~x6 | ~x3 | ~x4));
  assign n6475 = x3 ? (x4 | ~x5) : (~x4 ^ ~x5);
  assign n6476 = ~x2 & (x4 ? ~n6478 : ~n6477);
  assign n6477 = x1 ? (x0 ? (x6 | (~x3 ^ x5)) : (~x6 | (~x3 ^ ~x5))) : ((x5 | ~x6 | ~x0 | ~x3) & (x0 | (x3 ? (x5 | x6) : (~x5 | ~x6))));
  assign n6478 = (x0 | ~x1 | (x3 ? (x5 | x6) : (~x5 | ~x6))) & (x1 | (~x3 ^ ~x5) | (~x0 ^ ~x6));
  assign n6479 = ~x1 & (n6481 | n6482 | (~n1353 & ~n6480));
  assign n6480 = (~x0 | ~x2 | x7 | (~x3 ^ ~x5)) & (x0 | x2 | x3 | ~x5 | ~x7);
  assign n6481 = ~n1040 & (x0 ? (~x2 & n683) : (x2 & ~n1205));
  assign n6482 = n902 & ((n566 & n951) | (n564 & n978));
  assign n6483 = n6484 & (~x6 | n4077 | ~n626);
  assign n6484 = (n1682 | n2291) & (n623 | n2373);
  assign z357 = n6486 | ~n6497 | (x2 ? ~n6493 : ~n6489);
  assign n6486 = ~n643 & (x0 ? ~n6488 : ~n6487);
  assign n6487 = x2 ? ((~x4 | ~x5 | ~x1 | x3) & (x4 | ((~x3 | x5) & (x1 | (~x3 & x5))))) : ((~x4 | ~x5 | x1 | x3) & (~x1 | (x3 ? (~x4 | ~x5) : (~x4 ^ x5))));
  assign n6488 = (~x3 | x4 | x5 | ~x1 | x2) & (x1 | ((x2 | x4 | (~x3 ^ ~x5)) & (~x4 | (~x2 ^ (x3 & ~x5)))));
  assign n6489 = n6492 & (n1701 | n3541) & (x1 | n6490);
  assign n6490 = (~x0 | n6491) & (x0 | x3 | ~x5 | n3945);
  assign n6491 = x3 ? ((~x4 | x5 | ~x6 | ~x7) & (x4 | ~x5 | x6 | x7)) : ((~x6 | ~x7 | ~x4 | ~x5) & (x6 | x7 | x4 | x5));
  assign n6492 = (~x0 | ~x1 | x3 | n1282) & (x0 | (x1 ? (x3 | ~n993) : (~x3 | n1282)));
  assign n6493 = x1 ? (x0 | n6496) : (~n6494 & n6495);
  assign n6494 = ~n640 & ((n1121 & n825) | (n681 & n622));
  assign n6495 = x0 ? (x3 ? (x4 | n1701) : (~x4 | n2063)) : (x3 ? (x4 | n2063) : (~x4 | n1701));
  assign n6496 = x3 ? (x5 | ((~x6 | ~x7) & (~x4 | x6 | x7))) : (~x5 | ((x6 | x7) & (x4 | ~x6 | ~x7)));
  assign n6497 = (x2 & n6501) | (~x2 & ~n6498 & ~n6499 & n6500);
  assign n6498 = n1310 & (x1 ? (x3 & n1479) : (~x3 & ~n1408));
  assign n6499 = ~n2819 & ~n1682;
  assign n6500 = (x0 | x1 | ~x3 | n1040) & (~x0 | x3 | (x1 ? n1040 : ~n577));
  assign n6501 = (n3133 | ~n6502) & (~n543 | n877 | n1408);
  assign n6502 = ~x1 & (~x0 ^ ~x6);
  assign z358 = n6512 | ~n6514 | (~x2 & (~n6504 | ~n6509));
  assign n6504 = n6507 & (x3 | (~n6506 & (x0 | n6505)));
  assign n6505 = x1 ? ((x6 | x7 | ~x4 | ~x5) & (x4 | (x5 ? ~x6 : (x6 | x7)))) : ((~x4 | ~x5 | ~x6 | x7) & (x6 | ~x7 | x4 | x5));
  assign n6506 = ~x7 & n2061 & (x1 ? (~x4 & ~x6) : x6);
  assign n6507 = (n1337 | n6508) & (~n727 | ~n1621);
  assign n6508 = (~x0 | x3 | (~x1 ^ ~x6)) & (~x3 | ((x1 | ~x6) & (x0 | ~x1 | x6)));
  assign n6509 = (n671 | n6510) & (x1 | n6511);
  assign n6510 = (x3 | x5 | x0 | ~x1) & (~x0 | x1 | (~x3 ^ x5));
  assign n6511 = (x0 | x4 | (x3 ? (x5 | ~x7) : (~x5 | x7))) & (~x0 | ~x3 | ~x4 | ~x5 | ~x7);
  assign n6512 = x2 & (~n6513 | (~n1008 & ~n1721));
  assign n6513 = (~x3 | ~n717 | x0 | ~x1) & (x1 | x3 | ~n2209);
  assign n6514 = ~n6518 & (n1205 | n6516) & (n6515 | n6517);
  assign n6515 = (x1 | x6) & (x0 | ~x1 | ~x6);
  assign n6516 = x1 ? ((x4 | x5 | ~x0 | x2) & (x0 | ~x4 | (~x2 ^ x5))) : ((~x2 | x4 | ~x5) & (x0 | x2 | ~x4 | x5));
  assign n6517 = x2 ? ((x3 | ~x4 | ~x5 | x7) & (~x3 | x4 | x5 | ~x7)) : (~x3 | x4 | (~x5 ^ ~x7));
  assign n6518 = ~n765 & ((n1331 & n837) | (n5101 & ~n6519));
  assign n6519 = (x1 | ~x6) & (x0 | ~x1 | x6);
  assign z359 = ~n6529 | (x5 ? (n6521 | n6524) : ~n6525);
  assign n6521 = ~x2 & ((x4 & ~n6522) | (n828 & ~n6523));
  assign n6522 = (x0 | (x3 ? ((x6 | x7) & (x1 | ~x6 | ~x7)) : (~x6 ^ x7))) & (x1 | ~x3 | x6 | x7) & (x3 | ((x1 | (~x6 ^ x7)) & (~x0 | ~x1 | ~x6 | ~x7)));
  assign n6523 = (x6 | ~x7 | (~x0 & ~x1)) & (x0 | x7 | (~x1 ^ ~x6));
  assign n6524 = n1156 & ~n710 & (x3 ? (x6 ^ ~x7) : (x6 & ~x7));
  assign n6525 = x3 ? (~n6527 & ~n6528) : n6526;
  assign n6526 = (~n816 | ~n2834) & (n643 | n1918);
  assign n6527 = ~x0 & ((~x6 & ~x7 & x2 & x4) | (~x2 & x7 & (x4 ^ ~x6)));
  assign n6528 = n743 & ((n1445 & n1857) | (~x1 & n6470));
  assign n6529 = ~n6531 & (x3 | n6530) & (~n841 | n6532);
  assign n6530 = (x0 | ~x2 | (x4 ? (~x5 | ~x6) : x6)) & (x2 | ((x5 | x6 | x0 | ~x4) & (~x0 | ~x6 | (~x4 ^ x5))));
  assign n6531 = n825 & (x2 ? ~n1040 : n2359);
  assign n6532 = (~x2 | (x3 ? (~x4 | x6) : (x4 ? (~x5 | ~x6) : x6))) & (~x3 | x4 | ~x6 | (x2 & x5));
  assign z360 = n6546 | n6544 | n6541 | n6534 | n6538;
  assign n6534 = ~x2 & (~n6536 | (n757 & ~n6535));
  assign n6535 = x1 ? (x0 ? (x4 | x6) : (x3 ? ~x4 : (x4 | ~x6))) : ((~x0 | (~x3 ^ ~x4)) & (~x3 | ~x4 | x6));
  assign n6536 = x0 ? (~n550 | ~n1188) : (n6537 & (~n1188 | ~n2758));
  assign n6537 = (x6 | ~x7 | x3 | x4) & (~x3 | ~x6 | (x1 ? (x4 | x7) : (~x4 | ~x7)));
  assign n6538 = ~n1008 & (x1 ? ~n6540 : ~n6539);
  assign n6539 = (x0 | ((~x2 | ~x3 | ~x4 | x6) & (x4 | ~x6 | x2 | x3))) & (x2 | ~x3 | x4 | x6) & (~x2 | x3 | ~x4 | (~x0 & ~x6));
  assign n6540 = (~x0 | x2 | x3 | x4 | ~x6) & (x0 | ((x2 | ~x3 | x4 | x6) & (~x2 | ~x4 | (~x3 ^ x6))));
  assign n6541 = x2 & ((~x0 & ~n6542) | (n6352 & ~n6543));
  assign n6542 = (~x3 | ~x4 | ~x5 | ~x6 | x7) & (x3 | x6 | (x4 ? (x5 | ~x7) : x7));
  assign n6543 = x3 ? (~x4 | ~x5) : (x4 | x6);
  assign n6544 = ~n765 & (n2369 | (~n710 & (~n6545 | ~n920)));
  assign n6545 = (x2 | ~x3 | ~x4 | x6) & (x4 | ~x6 | ~x2 | x3);
  assign n6546 = ~n671 & (~n6547 | (n1322 & n1209));
  assign n6547 = (x0 | ~x2 | ~x3 | x5 | ~x6) & (~x0 | x2 | x3 | ~x5 | x6);
  assign z361 = n6555 | ~n6562 | (x3 ? ~n6549 : ~n6558);
  assign n6549 = (x1 & n6553) | (~n6551 & ~n6552 & ~x1 & ~n6550);
  assign n6550 = x2 & (n3333 | (n525 & n943));
  assign n6551 = n3476 & x0 & ~x2;
  assign n6552 = ~n1408 & (x0 ? (x2 & n1429) : (x2 ? n526 : n1429));
  assign n6553 = x0 ? (~n942 | ~n1084) : n6554;
  assign n6554 = x2 ? ((x4 | x5 | ~x6 | x7) & (x6 | ~x7 | ~x4 | ~x5)) : (~x4 | x7 | (~x5 ^ ~x6));
  assign n6555 = ~x0 & ((~x1 & ~n6556) | (n927 & ~n6557));
  assign n6556 = (x5 | ((x2 | x3 | x4 | ~x6) & (~x2 | ~x3 | ~x4 | x6))) & (~x3 | ~x5 | ((~x4 | ~x6) & (x2 | (~x4 & ~x6))));
  assign n6557 = (~x5 | ((x4 | ~x6) & (x2 | ~x4 | x6))) & (~x2 | ((~x5 | ~x6) & (~x4 | x5 | x6)));
  assign n6558 = ~n6560 & n6561 & (~n841 | n6559);
  assign n6559 = (x2 | x4 | ~x5 | ~x6 | x7) & (~x7 | ((~x5 | ~x6 | x2 | ~x4) & (~x2 | x5 | (~x4 ^ x6))));
  assign n6560 = x7 & n566 & ((~x5 & ~x6) | (~x2 & x5 & x6));
  assign n6561 = (~n733 | ~n2758) & (n990 | n1998);
  assign n6562 = (~n1365 | ~n6563) & (n2133 | (n710 & ~n837));
  assign n6563 = x5 & ((~x2 & x4 & ~x6) | (x6 & (x2 | ~x4)));
  assign z362 = ~n6576 | (x4 ? (n6569 | ~n6572) : ~n6565);
  assign n6565 = ~n6566 & (~n837 | ~n2888) & (n823 | n6568);
  assign n6566 = ~x0 & ((n676 & n951) | (~x2 & ~n6567));
  assign n6567 = (~x5 | ((x3 | ~x6 | ~x7) & (x1 | x6 | x7))) & (~x7 | (x1 ? (x3 | ~x6) : (x6 | (x3 & x5))));
  assign n6568 = (x6 | ((~x2 | ((x5 | ~x7) & (x3 | ~x5 | x7))) & (~x3 | (x5 ? x2 : ~x7)))) & (x2 | ~x5 | (x3 ? ~x7 : (~x6 | x7)));
  assign n6569 = ~x3 & ((~x2 & ~n6570) | (n1966 & ~n6571));
  assign n6570 = (~x0 | ~x7 | (x1 ? (x5 | ~x6) : (~x5 | x6))) & (x7 | (x0 ? (~x5 | (~x1 ^ x6)) : (x5 | (x1 & ~x6))));
  assign n6571 = (x1 | ~x6 | ~x7) & (x0 | (~x6 ^ ~x7));
  assign n6572 = (n1008 | n6573) & (~x3 | (~n6574 & ~n6575));
  assign n6573 = (x1 | ((~x6 | (~x2 ^ x3)) & (~x0 | ((~x3 | ~x6) & (x2 | x3 | x6))))) & (x0 | ((x3 | ~x6) & (~x2 | (x6 ? ~x1 : ~x3))));
  assign n6574 = ~n605 & ((n1857 & n841) | (n1300 & n543));
  assign n6575 = n2315 & ((~x5 & ~x7 & x0 & ~x2) | (x7 & ((x2 & x5) | (~x0 & (x2 | x5)))));
  assign n6576 = ~n6577 & (n6579 | (x0 ? (x3 | ~x7) : (~x3 | x7)));
  assign n6577 = ~n6578 & (n2402 | (~x4 & ~n1116));
  assign n6578 = (x0 & (x2 ? x1 : x3)) | (~x2 & ((x1 & x3) | (~x0 & ~x1 & ~x3)));
  assign n6579 = (x1 | ~x2 | x4 | ~x5 | ~x6) & (~x1 | x2 | ~x4 | (~x5 ^ ~x6));
  assign z365 = n6585 | n6584 | ~n2545 | n6581;
  assign n6581 = x6 & (n6582 | (n525 & ~n6583));
  assign n6582 = ~x0 & ((n809 & n979) | (~n697 & ~n2798));
  assign n6583 = (x1 | ~x2 | ~x3 | ~x5 | ~x7) & (x3 | ((x5 | x7 | ~x1 | x2) & (x1 | ((x5 | ~x7) & (x2 | ~x5 | x7)))));
  assign n6584 = ~n1218 & ((n560 & n624) | (n742 & ~n1262));
  assign n6585 = ~x6 & (n6586 | (n750 & n774 & n816));
  assign n6586 = ~x3 & ((n733 & n867) | (n1477 & ~n6587));
  assign n6587 = (~x0 | x1 | x7) & (~x2 | ~x7 | x0 | ~x1);
  assign z366 = ~n2567 | n6589 | (x4 & ~n6591);
  assign n6589 = n1835 & ((n560 & n2575) | (~x0 & ~n6590));
  assign n6590 = (~x5 | ((~x2 | ~x3 | ~x7) & (~x1 | (~x3 ^ ~x7)))) & (x1 | x5 | ((x3 | ~x7) & (x2 | ~x3 | x7)));
  assign n6591 = x5 ? (~x6 | n6594) : (~n6592 & ~n6593);
  assign n6592 = ~n2341 & ((n632 & n1465) | (n570 & n1903));
  assign n6593 = n1686 & ((~x1 & x2 & n1465) | (~x2 & n1903));
  assign n6594 = (x0 | ~x1 | ~x2 | ~x3 | ~x7) & (~x0 | x1 | ((~x3 | ~x7) & (~x2 | x3 | x7)));
  assign z367 = n6596 | n6600 | ~n6604 | (x1 & ~n6602);
  assign n6596 = ~x2 & (n6597 | (n1005 & ~n6599));
  assign n6597 = ~x3 & (x0 ? (n1145 & n978) : ~n6598);
  assign n6598 = (x1 | ~x4 | x5 | x6 | x7) & (~x7 | ((~x1 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (x5 | x6 | x1 | x4)));
  assign n6599 = (~x0 | ~x1 | x4 | x5 | x7) & ((~x4 ^ x7) | (x0 ? (x1 | ~x5) : (~x1 ^ ~x5)));
  assign n6600 = ~n1218 & ((n3848 & n837) | (x6 & ~n6601));
  assign n6601 = (x0 | ~x3 | ((x2 | x5) & (~x1 | ~x2 | ~x5))) & (x1 | (x0 ? (~x5 | (~x2 & ~x3)) : (~x2 | x5)));
  assign n6602 = (~x4 | n6603) & (x2 | x4 | ~x5 | n4925);
  assign n6603 = (x0 | ((x2 | x3 | ~x5 | x6) & (~x2 | x5 | ~x6))) & (~x0 | x2 | x3 | ~x6);
  assign n6604 = ~n2598 & ~n6605 & ~n6608 & (x4 | n6610);
  assign n6605 = n3431 & ((n566 & n6606) | (x7 & ~n6607));
  assign n6606 = x5 & ~x7 & (x1 | x3);
  assign n6607 = (x1 | x5 | (x0 ? (~x3 | ~x4) : (x3 | x4))) & (x0 | x4 | ~x5 | (~x1 & ~x3));
  assign n6608 = ~x1 & ((n704 & n547) | (n1005 & ~n6609));
  assign n6609 = (~x0 | ~x2 | x4 | ~x5) & (x0 | (x2 ? (x4 | x5) : (~x4 | ~x5)));
  assign n6610 = (x1 | (x0 ? (x6 | (x3 & x5)) : (~x5 | ~x6))) & (x0 | ((x3 | ~x5 | ~x6) & (~x1 | x5 | x6)));
  assign z368 = (~x3 | ~n6620) & (x3 | n6612 | n6614 | ~n6615);
  assign n6612 = ~x5 & ((n548 & n733) | (~x7 & ~n6613));
  assign n6613 = (~x1 | x2 | x4 | ~x6) & (x1 | x6 | (x0 ? x4 : (~x2 | ~x4)));
  assign n6614 = n691 & (x0 ? (~x1 & n2834) : (x1 & ~n3319));
  assign n6615 = ~n6616 & ~n6617 & n6618 & (n1431 | n2357);
  assign n6616 = x6 & ((~x0 & (x1 ? (x2 & ~x5) : (~x2 & x5))) | (x0 & x1 & ~x2 & x5));
  assign n6617 = ~n1008 & ((n922 & n878) | (n626 & ~n784));
  assign n6618 = ~n6619 & (~x7 | ~n1310 | n1185);
  assign n6619 = ~x6 & x5 & x0 & ~x1;
  assign n6620 = ~n6622 & ~n6623 & n6624 & (n643 | n6621);
  assign n6621 = (~x0 | x1 | ~x2 | ~x4 | x5) & (x0 | ~x5 | (x1 ^ ~x2));
  assign n6622 = ~n640 & ((n841 & n1966) | (~x0 & n2849));
  assign n6623 = n5017 & ((n569 & n570) | (n1769 & n632));
  assign n6624 = (x0 | x1 | x2 | (~x5 ^ x7)) & ((x0 ? (x1 | x2) : (~x1 | ~x2)) | (~x5 ^ ~x7));
  assign z369 = n6626 | n6631 | ~n6636 | (~n643 & ~n6634);
  assign n6626 = ~x1 & (n6627 | n6630);
  assign n6627 = x0 & ((~n3929 & ~n6628) | (~x3 & ~n6629));
  assign n6628 = x3 ? (x4 | x5) : (x4 ^ ~x5);
  assign n6629 = x6 ? (~x7 | (~x2 & (x4 | x5))) : (x7 | ((~x4 | ~x5) & (x2 | (~x4 & ~x5))));
  assign n6630 = ~x3 & n742 & (n3687 | (~n640 & ~n3754));
  assign n6631 = n543 & (x5 ? (n1044 & ~n6633) : ~n6632);
  assign n6632 = (~x2 | ~x3 | x4 | ~x6 | ~x7) & (x3 | ((x4 | x6 | x7) & (x2 | ((x6 | x7) & (~x4 | ~x6 | ~x7)))));
  assign n6633 = (~x4 | x6 | x7) & (~x6 | ~x7);
  assign n6634 = x2 ? (~n543 | (x3 & ~n1716)) : n6635;
  assign n6635 = (~x0 | ((~x3 | x4 | x5) & (~x1 | x3 | ~x4))) & (x3 | ((~x5 | (~x1 ^ x4)) & (x0 | (x1 & x4))));
  assign n6636 = (~n837 | ~n846) & (~x3 | (~n6637 & ~n6638));
  assign n6637 = ~x1 & ~n815 & (~x0 | n525 | n2332);
  assign n6638 = n543 & ((x2 & x6 & (x4 | n1364)) | (~x6 & (~x2 | (~x4 & n1364))));
  assign z370 = ~n6642 | (n681 & (x1 ? ~n6640 : ~n6641));
  assign n6640 = (~x0 | x2 | x3 | x6 | ~x7) & (x0 | (x3 ? ((x6 | x7) & (~x2 | ~x6 | ~x7)) : (~x6 | x7)));
  assign n6641 = x3 ? ((x0 | ~x2 | x6 | x7) & (~x0 | ((~x6 | ~x7) & (x2 | x6 | x7)))) : ((~x6 | x7) & (~x0 | x6 | ~x7));
  assign n6642 = n6646 & (~n632 | n6643) & (x4 | n6644);
  assign n6643 = (~x0 | x3 | ~x4 | x7) & (x0 | ~x3 | x4 | ~x7);
  assign n6644 = x7 ? (~n1301 | (~n841 & ~n746)) : n6645;
  assign n6645 = (x3 & x5) | (x0 & x1 & x2) | (~x5 & (~x0 | ~x3 | (~x1 & ~x2)));
  assign n6646 = (x0 | x1 | ~x3 | ~x7) & (~x4 | (x0 & x1) | (~x3 ^ ~x7));
  assign z371 = ~n6650 | (~x4 & (n4313 | n6648));
  assign n6648 = ~x5 & (x3 ? (n1857 & n816) : ~n6649);
  assign n6649 = (~x0 | ~x6 | (x1 ? (x2 | ~x7) : (~x2 | x7))) & (x0 | ~x1 | ~x2 | x6 | ~x7);
  assign n6650 = n6652 & (x5 | (n4986 & n6651));
  assign n6651 = (~n816 | ~n1395) & (n671 | n2530);
  assign n6652 = ~n6653 & (~n841 | ~n926) & (~n779 | ~n6654);
  assign n6653 = ~x4 & ((~x1 & x5) | (~x0 & (x5 | x6)));
  assign n6654 = x4 & ~x3 & ~x2 & x0 & x1;
  assign z372 = ~n6659 | (~x3 & ~n6656) | (~n1008 & ~n6658);
  assign n6656 = (~n845 | ~n746) & (x1 | x7 | n6657);
  assign n6657 = (x0 | x2 | ~x4 | x5 | x6) & (~x0 | ~x2 | ~x6 | (~x4 ^ ~x5));
  assign n6658 = x0 ? (~x6 | (x1 ? (x2 | x3) : (~x2 | ~x3))) : (x6 | (x1 ^ ~x2));
  assign n6659 = n6660 & ~n6661 & ~n6662 & (~n878 | n3095);
  assign n6660 = x0 ? (x1 | x2 | (~x5 ^ x6)) : (~x1 | ((x5 | ~x6) & (~x2 | ~x5 | x6)));
  assign n6661 = n757 & n689 & (x0 ? n865 : n878);
  assign n6662 = ~x1 & ((x0 & x2 & x5 & ~x6) | (~x0 & ~x5 & x6));
  assign z373 = ~n6667 | (~x5 & ~n6664);
  assign n6664 = x0 ? n6665 : (~n6666 & (~n558 | ~n1395));
  assign n6665 = (~n1786 | ~n979) & (~n676 | ~n1668);
  assign n6666 = ~n643 & ((n828 & n1133) | n676 | n979);
  assign n6667 = ~n6668 & n6669 & ~n6672 & (x3 | n6671);
  assign n6668 = ~n4282 & x5 & n939;
  assign n6669 = n6670 & (n3152 | (n3275 & (~n570 | ~n959)));
  assign n6670 = (x0 | ~x3 | (x1 ? (~x2 | ~x6) : (x2 | x6))) & (~x0 | x1 | x2 | ~x6);
  assign n6671 = (x0 | ~x4 | (x1 ? (~x2 | ~x6) : (x2 | x6))) & (~x0 | x1 | ~x2 | x4 | ~x6);
  assign n6672 = n1380 & ((n669 & n1585) | (~n643 & ~n6673));
  assign n6673 = (~x1 | x2 | ~x3) & (x3 | x4 | x1 | ~x2);
  assign z374 = ~n6676 | ~n6679 | (~x7 & ~n6675);
  assign n6675 = (x0 | x1 | x2 | ~x3 | x4) & (x3 | ((~x0 | x1 | ~x2 | x4) & (x0 | ~x4 | (~x1 ^ ~x2))));
  assign n6676 = ~n2507 & n6677 & n6678 & (~n841 | ~n1080);
  assign n6677 = (~n1209 | ~n5802) & (~n543 | ~n1413);
  assign n6678 = ~x7 | ((x1 | ~x2 | ~x3) & (~x1 | x2 | x3) & (x0 | (x1 ^ ~x2)));
  assign n6679 = (x1 | n6681) & (x0 | (~n6680 & (x1 | ~n911)));
  assign n6680 = n828 & (x1 ? (x2 & ~n1008) : (~x2 & n750));
  assign n6681 = (~n1693 | ~n610) & (~n1451 | n6682);
  assign n6682 = (x0 | x2 | x4 | ~x6 | x7) & (~x0 | ~x2 | ~x4 | (~x6 ^ ~x7));
  assign z375 = n6684 | n6687 | ~n6689 | (~x0 & ~n6688);
  assign n6684 = ~x2 & (n6685 | (n830 & n1234));
  assign n6685 = x5 & ((n3261 & n873) | (n527 & ~n6686));
  assign n6686 = (~x0 | (x3 ? (x4 | ~x7) : (~x4 | x7))) & (x0 | ~x3 | ~x4 | x7);
  assign n6687 = ~x4 & ((n1322 & n1269) | (~x2 & ~n5999));
  assign n6688 = (x4 | x5 | ~x1 | x3) & (x1 | ~x3 | (x2 ? (x4 | ~x5) : (~x4 | x5)));
  assign n6689 = n6691 & ~n6690 & n5322 & ~n3279 & ~n5363;
  assign n6690 = ~x2 & x4 & (x0 ? (x1 ^ x3) : (x1 ^ ~x3));
  assign n6691 = (~n1209 | ~n3217) & (~n662 | ~n1644);
  assign z376 = ~n6698 | (~x2 & (~n6693 | ~n6697));
  assign n6693 = x5 ? (~n6696 & (~n699 | ~n1585)) : n6694;
  assign n6694 = (~n550 | ~n1234) & (~x7 | n6695);
  assign n6695 = (x0 | x1 | x3 | x4 | x6) & ((x0 ^ ~x3) | (x1 ? (~x4 | x6) : (x4 | ~x6)));
  assign n6696 = n1188 & ((n1857 & n566) | (x0 & ~n3098));
  assign n6697 = (~x0 | ((~x1 | x3 | ~x4 | ~x5) & (x1 | ~x3 | x4 | x5))) & (x4 | ~x5 | x1 | x3) & (x0 | ((x1 | x4 | ~x5) & (~x4 | (x1 ? (~x3 ^ ~x5) : (~x3 | x5)))));
  assign n6698 = ~n6699 & ~n6703 & n6704 & (~x2 | n6702);
  assign n6699 = ~x5 & ((~x1 & ~n6700) | (n632 & ~n6701));
  assign n6700 = (~x0 | ~x2 | x3 | ~x4 | x6) & (x0 | x4 | (x2 ? (~x3 | x6) : (x3 | ~x6)));
  assign n6701 = (~x4 | ~x6 | x0 | ~x3) & (~x0 | (x3 ? (x4 | x6) : (~x4 | ~x6)));
  assign n6702 = (x0 | ~x1 | x3 | x4 | x5) & (x1 | ~x3 | (x0 ? (~x4 ^ x5) : (~x4 | ~x5)));
  assign n6703 = ~x3 & ((~x0 & x1 & ~x2 & ~x4) | (~x1 & (x0 ? (x2 ^ x4) : (x2 & x4))));
  assign n6704 = ~n932 & (~n1121 | (n6705 & (~n569 | ~n1644)));
  assign n6705 = (~x0 | x1 | ~x2 | ~x3 | x6) & (x0 | ~x1 | x3 | (~x2 ^ ~x6));
  assign z377 = n6707 | ~n6711 | ~n6716 | (n3034 & ~n6710);
  assign n6707 = ~x1 & (~n6709 | (~x3 & ~n6708));
  assign n6708 = (x0 | ~x2 | x4 | x5 | ~x6) & (~x0 | ((~x2 | (x4 ? (x5 | x6) : (~x5 | ~x6))) & (x2 | ~x4 | x5 | ~x6)));
  assign n6709 = (x0 | x3 | x4 | ~x5 | x6) & (~x3 | ((x5 | ~x6 | x0 | ~x4) & (~x0 | x6 | (~x4 ^ ~x5))));
  assign n6710 = (x3 | x4 | ~x5 | x6 | ~x7) & (~x4 | ((~x6 | ~x7 | x3 | ~x5) & (~x3 | (x5 ? (~x6 | x7) : (x6 | ~x7)))));
  assign n6711 = ~n6712 & ~n6714 & ~n6715 & (n615 | n6713);
  assign n6712 = ~x0 & ((~x1 & x3 & ~x5 & ~x6) | (x6 & (x1 ? (x3 ^ ~x5) : (~x3 & x5))));
  assign n6713 = (x0 | ~x2 | ~x7 | (~x1 ^ x5)) & (~x0 | ~x1 | x2 | x5 | x7);
  assign n6714 = x6 & ~x5 & x3 & x0 & ~x1;
  assign n6715 = n1044 & ((n543 & n706) | (x0 & ~n623));
  assign n6716 = (~n4137 | n6717) & (x2 | (~n6718 & ~n6720));
  assign n6717 = (x0 | ~x2 | x3 | ~x4 | ~x5) & (x4 | (x0 ? (x2 | (~x3 ^ x5)) : ((~x3 | ~x5) & (~x2 | x3 | x5))));
  assign n6718 = ~x0 & ((n2980 & ~n5129) | (n750 & ~n6719));
  assign n6719 = (x1 | ~x3 | ~x4 | x6) & (~x1 | x3 | ~x6);
  assign n6720 = n6352 & (n1228 | (x5 & (n1331 | n5072)));
  assign z378 = n6726 | n6729 | ~n6731 | (~x1 & ~n6722);
  assign n6722 = x0 ? (~n6725 & (~n1044 | ~n1668)) : n6723;
  assign n6723 = ~n6724 & (~n813 | ~n949) & (~n1518 | ~n1070);
  assign n6724 = x2 & (x4 ? (x6 & (~x5 | x7)) : (~x5 & ~x6));
  assign n6725 = n4817 & (n629 | (~x2 & n4604));
  assign n6726 = ~n643 & (~n6728 | (~x2 & ~n6727));
  assign n6727 = (x3 | x4 | ~x0 | x1) & (x0 | ((x1 | ~x3 | x4 | ~x5) & (~x1 | (x3 ? (x4 | x5) : ~x5))));
  assign n6728 = x0 ? ((x1 | ~x4 | ~x5) & (~x1 | x2 | x4 | x5)) : (x4 | (x1 ? (~x2 | x5) : (~x2 ^ ~x5)));
  assign n6729 = n543 & ((n658 & n1556) | (~x5 & ~n6730));
  assign n6730 = (~x6 | ~x7 | ~x2 | ~x4) & (x2 | x3 | x6 | (x4 & x7));
  assign n6731 = (n2803 | n6732) & (n1850 | n6733);
  assign n6732 = (~x5 & ((x1 & x2 & x3) | (~x1 & ~x2 & ~x3) | (~x0 & (~x1 | (~x2 & ~x3))))) | (~x0 & ~x1 & x2 & x3) | (x0 & ((~x2 & x3 & x5) | (x1 & (x2 | x3))));
  assign n6733 = (~x2 | ((x0 | ~x1 | ~x5) & (x3 | x5 | ~x0 | x1))) & (x0 | ~x1 | ~x3 | ~x5) & (x2 | ((x0 | x1 | x3 | ~x5) & (~x0 | (x1 ? (x3 | ~x5) : (~x3 | x5)))));
  assign z379 = n6735 | ~n6738 | n6749 | (~x4 & ~n6744);
  assign n6735 = ~n1198 & ((x4 & ~n6736) | (n1084 & ~n6737));
  assign n6736 = x1 ? ((x2 | x3 | ~x7) & (x0 | (x2 ? (~x3 | x7) : ~x7))) : ((x2 | x3 | x7) & (~x3 | ~x7 | ~x0 | ~x2));
  assign n6737 = (x0 & x3) | (x1 & ~x7) | (x7 & (~x1 | (~x0 & ~x3)));
  assign n6738 = ~n6739 & (n1548 | n6742) & (~n543 | n6743);
  assign n6739 = ~x1 & ((x2 & ~n6740) | (n691 & ~n6741));
  assign n6740 = (x0 | ~x3 | ~x4 | x5 | ~x7) & (x3 | x4 | ((~x5 | x7) & (~x0 | x5 | ~x7)));
  assign n6741 = (x0 | x3 | ~x7) & (~x3 | x7 | (~x0 & ~x4));
  assign n6742 = (~x0 | ~x1 | x2 | x5 | x7) & (~x2 | ((x1 | x5 | ~x7) & (x0 | (x1 ? (~x5 ^ ~x7) : (~x5 | x7)))));
  assign n6743 = (~x2 | ~x5 | ~x7 | (~x3 ^ ~x4)) & (x5 | ((x4 | x7 | ~x2 | x3) & (x2 | (x3 ? (~x4 | x7) : (x4 | ~x7)))));
  assign n6744 = x0 ? n6747 : (~n6745 & (~x1 | n6746));
  assign n6745 = ~n1097 & ((~x3 & ~x7 & x1 & ~x2) | (~x1 & x7 & (~x2 ^ ~x3)));
  assign n6746 = (x2 | ~x3 | x5 | x6 | x7) & (~x2 | ((~x6 | ~x7 | x3 | x5) & (x6 | x7 | ~x3 | ~x5)));
  assign n6747 = (~n576 | ~n813) & (~n6748 | (~n572 & ~n1413));
  assign n6748 = ~x1 & (x5 ^ ~x6);
  assign n6749 = x4 & (n6751 | (~n1097 & ~n6750));
  assign n6750 = (x0 | ~x1 | x2 | x3 | x7) & (x1 | ((~x3 | ~x7 | x0 | x2) & (~x0 | (x2 ? (~x3 | x7) : (x3 | ~x7)))));
  assign n6751 = ~x1 & ((n852 & n2264) | (x0 & ~n1635));
  assign z380 = n6753 | n6757 | ~n6760 | (~n643 & ~n6756);
  assign n6753 = x0 & (n6754 | (n676 & n2402));
  assign n6754 = ~x2 & ((n943 & n3194) | (~x7 & ~n6755));
  assign n6755 = (x1 | ~x3 | ~x4 | ~x5 | x6) & (~x1 | x4 | x5 | (x3 ^ ~x6));
  assign n6756 = (~x2 | (x0 ? (x1 | (~x3 ^ x4)) : (~x3 | (~x1 & ~x4)))) & (x0 | x2 | x3 | (x1 & x4));
  assign n6757 = ~x0 & ~n6758;
  assign n6758 = x1 ? ((~n1966 | n1967) & (x4 | n6759)) : (~x4 | n6759);
  assign n6759 = (x2 | ~x3 | x5 | ~x6 | x7) & (~x2 | x6 | (x3 ? (x5 | x7) : (~x5 | ~x7)));
  assign n6760 = ~n6764 & ~n6766 & n6767 & (n640 | n6761);
  assign n6761 = ~n6762 & (~n626 | ~n1780) & (x5 | n6763);
  assign n6762 = ~x2 & ((~x0 & x1 & x3 & x4) | (x0 & (x1 ? (~x3 & x4) : (x3 & ~x4))));
  assign n6763 = (x0 | ~x1 | ~x2 | x3 | x4) & (~x0 | x1 | x2 | ~x3 | ~x4);
  assign n6764 = ~n6765 & x7 & n778;
  assign n6765 = (x3 | x4 | ~x0 | ~x1) & (x0 | ~x3 | (~x1 ^ x4));
  assign n6766 = ~n815 & ~n3495;
  assign n6767 = (~n1269 | ~n1525) & (~x6 | n2726 | ~n2742);
  assign z381 = n6770 | ~n6772 | ~n6779 | (n825 & ~n6769);
  assign n6769 = (x1 | x2 | ~x4 | x5 | x7) & (~x1 | ((x5 | x7 | x2 | x4) & (~x2 | ~x7 | (~x4 ^ x5))));
  assign n6770 = ~x3 & ((~n1538 & n5463) | (x0 & ~n6771));
  assign n6771 = (~x1 | x2 | x4 | x5 | x7) & (x1 | ~x2 | ~x4 | ~x5 | ~x7);
  assign n6772 = ~n6773 & ~n6775 & n6776 & (n1008 | n6763);
  assign n6773 = x7 & ~n6774;
  assign n6774 = (~x0 | ~x1 | x2 | x3 | ~x4) & (x0 | ((x3 | ~x4 | x1 | x2) & ((~x3 ^ ~x4) | (x1 ^ ~x2))));
  assign n6775 = ~x1 & ~x4 & (x0 ? (x3 ^ ~x7) : (x3 & ~x7));
  assign n6776 = ~n6777 & (~n587 | ~n2402) & (~n2742 | ~n6778);
  assign n6777 = ~x7 & x4 & ~x3 & ~x0 & x1;
  assign n6778 = ~x7 & (x2 ^ ~x3);
  assign n6779 = ~n6780 & (~x7 | (~n6782 & ~n6783));
  assign n6780 = ~n640 & ((n622 & ~n1284) | (~x0 & n6781));
  assign n6781 = x3 & ((x1 & ~x4 & (~x2 ^ ~x5)) | (~x1 & ~x2 & x4 & x5));
  assign n6782 = ~x2 & (x0 ? ~n897 : (n704 & n689));
  assign n6783 = ~n5565 & n742 & n1479;
  assign z382 = n6789 | n6792 | (x7 ? ~n6785 : ~n6796);
  assign n6785 = x1 ? (~x4 | n6788) : (x4 ? n6786 : n6787);
  assign n6786 = (x0 | x2 | x3 | x5 | x6) & (~x0 | ~x2 | ~x3 | ~x5 | ~x6);
  assign n6787 = (x0 | x2 | ~x3 | ~x5 | ~x6) & (x5 | ((x0 | x2 | x3 | x6) & (~x0 | ~x2 | (~x3 ^ x6))));
  assign n6788 = (~x0 | x2 | x3 | ~x5 | x6) & (x0 | (~x2 ^ x5) | (~x3 ^ x6));
  assign n6789 = ~x1 & (~n6791 | (~x2 & ~n6790));
  assign n6790 = x0 ? ((x4 | ~x5 | ~x6) & (x3 | ~x4 | x5 | x6)) : (~x4 | ~x5 | (x3 ^ ~x6));
  assign n6791 = (~x3 | (x2 ? (x4 | ~x6) : (~x4 | x5))) & (~x2 | ((x4 | ~x5) & (x3 | ~x4 | x5 | x6))) & (x2 | ~x4 | ((x5 | ~x6) & (x3 | ~x5 | x6)));
  assign n6792 = x1 & (n6793 | n6794 | ~n6795);
  assign n6793 = ~x0 & ((x2 & ~x3 & x4 & x5) | (~x4 & ((~x3 & ~x5) | (~x2 & (~x3 | ~x5)))));
  assign n6794 = ~n1353 & ((~x3 & x5 & x0 & ~x2) | (~x0 & x3 & (x2 ^ x5)));
  assign n6795 = ~n730 & (~n1005 | n1426);
  assign n6796 = (~n1269 | ~n1748) & (~x6 | n6797);
  assign n6797 = (x0 | ~x2 | ~x4 | n5565) & (~x0 | x2 | n6798);
  assign n6798 = (x1 | x3 | ~x4 | ~x5) & (x4 | x5 | ~x1 | ~x3);
  assign z383 = ~n6810 | n6800 | ~n6803;
  assign n6800 = x1 & (n3926 | (~x0 & (n6801 | n6802)));
  assign n6801 = ~n627 & ((n750 & n1518) | (x2 & ~n1014));
  assign n6802 = x6 & ((n674 & n885) | (~x2 & n2296));
  assign n6803 = ~n6804 & ~n6807 & ~n6809 & (x3 | n6808);
  assign n6804 = x4 & (x2 ? ~n6805 : ~n6806);
  assign n6805 = (x0 | x1 | x3 | x5 | x6) & (~x5 | (~x0 ^ x1) | (~x3 ^ x6));
  assign n6806 = (~x0 | x1 | x3 | x5 | ~x6) & (x0 | ((~x3 | x5 | ~x6) & (x1 | x3 | ~x5 | x6)));
  assign n6807 = ~n1008 & ((n1141 & n816) | (n525 & ~n1009));
  assign n6808 = (x6 | (~x0 ^ x1) | (~x2 ^ x5)) & (x2 | ~x6 | (x0 ? (~x1 | x5) : (x1 | ~x5)));
  assign n6809 = n1188 & ((~x5 & x6 & x0 & ~x2) | (~x0 & x5 & (x2 ^ ~x6)));
  assign n6810 = ~n6811 & (x1 | (~x2 & n6815) | (x2 & n6814));
  assign n6811 = ~x4 & (x1 ? ~n6812 : ~n6813);
  assign n6812 = (x0 | ~x2 | (x3 ? (~x5 ^ ~x6) : (x5 | ~x6))) & (x2 | ((~x5 | ~x6 | x0 | x3) & (x6 | (x0 ? (~x3 ^ x5) : (~x3 | ~x5)))));
  assign n6813 = (x0 | ~x2 | x3 | x5 | ~x6) & (~x3 | ((x0 | ~x2 | x5 | x6) & (~x0 | ~x5 | (~x2 ^ ~x6))));
  assign n6814 = (~n5168 | ~n951) & (n765 | n627 | n807);
  assign n6815 = (x3 | n6816) & (~x4 | ~n951 | ~x0 | ~x3);
  assign n6816 = x0 ? (~x6 | (x4 ? (~x5 | x7) : (x5 | ~x7))) : (x6 | (x4 ? (x5 | x7) : ~x7));
  assign z384 = n6823 | ~n6826 | (~x1 & ~n6818);
  assign n6818 = x5 ? (x2 ? n6820 : n6819) : n6821;
  assign n6819 = (x0 | ~x3 | x4 | (~x6 ^ x7)) & (~x4 | (x0 ? (x3 ? (~x6 | ~x7) : (x6 | x7)) : (x3 | ~x6)));
  assign n6820 = (~x0 | ~x3 | ~x4 | x6 | ~x7) & (x0 | x3 | (x4 ? (x6 | ~x7) : ~x6));
  assign n6821 = (~n1693 | ~n3790) & (x4 | n6822);
  assign n6822 = (~x0 | x2 | x3 | ~x6 | x7) & (x6 | (x0 ? (x2 | (~x3 & ~x7)) : (~x2 | ~x3)));
  assign n6823 = n543 & (x7 ? ~n6825 : ~n6824);
  assign n6824 = (x2 | ~x3 | x4 | (~x5 ^ x6)) & (x3 | ~x4 | ((x5 | ~x6) & (~x2 | ~x5 | x6)));
  assign n6825 = (x2 | ~x3 | ~x4 | x5 | x6) & (x3 | ((~x5 | ~x6 | x2 | x4) & (x5 | (x2 ? (~x4 ^ x6) : (~x4 | ~x6)))));
  assign n6826 = ~n6827 & ~n6831 & n6834 & (n3319 | n6833);
  assign n6827 = ~n640 & ((~x1 & ~n6828) | ~n6830 | (x1 & ~n6829));
  assign n6828 = x2 ? ((~x4 | ~x5 | ~x0 | x3) & (x0 | x4 | (~x3 ^ ~x5))) : ((~x0 | ((~x3 | x4 | ~x5) & (~x4 | x5))) & (x3 | ~x4 | x5) & (x0 | ~x5 | (~x3 ^ ~x4)));
  assign n6829 = (x0 | ~x2 | ~x3 | ~x4 | x5) & (~x0 | x2 | x3 | x4 | ~x5);
  assign n6830 = x0 ? ((x1 | ~x2 | ~x3 | x4) & (~x1 | x2 | x3 | ~x4)) : (~x3 | (x1 ? (~x2 ^ x4) : (~x2 | ~x4)));
  assign n6831 = ~x3 & ((n543 & n550) | (~x1 & ~n6832));
  assign n6832 = (x0 | ~x2 | ~x4 | ~x6 | x7) & (~x0 | ((~x2 | x4 | ~x6 | x7) & (x2 | ~x4 | x6 | ~x7)));
  assign n6833 = (x0 | ~x2 | ~x3 | (x1 ^ ~x5)) & (x2 | ~x5 | (x1 ? x3 : ~x0));
  assign n6834 = (n871 | n6836) & (~x7 | n2208 | ~n6835);
  assign n6835 = ~x6 & x3 & ~x0 & ~x2;
  assign n6836 = x0 ? ((~x1 | x2 | x4 | x5) & (x1 | ~x2 | (~x4 & ~x5))) : ((~x4 | ~x5 | ~x1 | ~x2) & (x4 | x5 | x1 | x2));
  assign z385 = n6854 | n6851 | n6848 | n6838 | n6845;
  assign n6838 = ~x6 & (n6839 | ~n6841);
  assign n6839 = ~x2 & ((n2296 & n727) | (~x3 & ~n6840));
  assign n6840 = (~x0 | x1 | (x4 ? (x5 | ~x7) : (~x5 | x7))) & (~x1 | ((~x0 | ~x4 | ~x5 | x7) & (x0 | ~x7 | (~x4 ^ ~x5))));
  assign n6841 = (n807 | n6843) & (~n6842 | n6844);
  assign n6842 = x2 & x7;
  assign n6843 = (~x1 | x2 | ~x3 | x5 | ~x7) & (x1 | ((x2 | ~x3 | ~x5 | ~x7) & (~x2 | (x3 ? (~x5 | x7) : (x5 | ~x7)))));
  assign n6844 = (~x0 | x1 | ~x3 | ~x4 | x5) & (x0 | x4 | (x1 ? (~x3 ^ x5) : (~x3 | ~x5)));
  assign n6845 = ~n765 & (~n6847 | (~x6 & ~n6846));
  assign n6846 = (x0 | ~x1 | ~x2 | ~x3 | ~x4) & (~x0 | x3 | (x1 ? (x2 | x4) : (~x2 | ~x4)));
  assign n6847 = x0 ? ((~x1 | x2 | x3 | ~x4) & (x1 | (x2 ? (~x3 | x4) : (~x3 ^ ~x4)))) : (x1 ? (x2 ? (x3 | ~x4) : (~x3 | x4)) : (x2 ? (~x3 ^ ~x4) : (x3 | ~x4)));
  assign n6848 = n569 & ((n543 & ~n6850) | (~x1 & ~n6849));
  assign n6849 = (x0 | x4 | (x2 ? (~x3 | ~x5) : (~x3 ^ x5))) & ((x0 ^ ~x4) | (x2 ? (x3 | x5) : (~x3 | ~x5)));
  assign n6850 = (x4 | ~x5 | ~x2 | x3) & (x2 | ~x4 | (~x3 ^ x5));
  assign n6851 = ~x1 & (n6852 | ~n6853 | (~n2466 & ~n1337));
  assign n6852 = ~n1998 & ~n4754;
  assign n6853 = (~n2296 | ~n547) & (~n674 | ~n549);
  assign n6854 = x1 & (x0 ? (n2296 & n1044) : ~n6855);
  assign n6855 = (x2 | ~x3 | ~x4 | ~x5 | x7) & (~x2 | x3 | x4 | x5 | ~x7) & ((~x2 ^ ~x3) | (x4 ? (x5 | ~x7) : (~x5 | x7)));
  assign z386 = n6868 | n6866 | ~n6862 | n6857 | n6859;
  assign n6857 = ~x2 & ((n1358 & n727) | (~x5 & ~n6858));
  assign n6858 = (~x0 | ~x1 | ~x3 | x4 | x6) & (x1 | x3 | ~x6 | (x0 & x4));
  assign n6859 = ~n1408 & ((n742 & ~n6861) | (~x2 & ~n6860));
  assign n6860 = (x0 | ~x1 | ~x3 | ~x5 | ~x7) & (~x0 | ((~x1 | x3 | ~x5 | x7) & (x1 | ~x3 | x5 | ~x7)));
  assign n6861 = (x1 | x3 | ~x5 | ~x7) & (~x1 | x5 | (~x3 ^ x7));
  assign n6862 = ~n6863 & ~n6864 & n6865 & (n1097 | n5015);
  assign n6863 = ~n752 & (n769 | (x7 & n1181 & ~n2290));
  assign n6864 = n742 & ((n1358 & n927) | (n704 & n689));
  assign n6865 = (n1036 | n2077) & (n1100 | ~n3416);
  assign n6866 = ~n1026 & ((n837 & n2209) | (~x1 & ~n6867));
  assign n6867 = (x0 | ~x2 | x4 | x5 | ~x7) & (~x4 | ((~x0 | (x2 ? (x5 | x7) : (~x5 | ~x7))) & (x0 | x2 | x5 | ~x7)));
  assign n6868 = ~x7 & ((~n6869 & n2320) | (~x1 & ~n6870));
  assign n6869 = (x4 | x5 | x2 | x3) & (~x4 | ~x5 | ~x2 | ~x3);
  assign n6870 = (~n1358 | ~n2435) & (~n1044 | (~n2820 & ~n5036));
  assign z387 = n6872 | n6876 | ~n6882 | (~n3319 & ~n6881);
  assign n6872 = ~n640 & (n6874 | n6875 | (~x0 & ~n6873));
  assign n6873 = (~x4 | (x1 ? (~x2 | x5) : (x2 ? ~x3 : (x3 | x5)))) & (x1 | x2 | ~x3 | x4) & (~x5 | ((x2 | x3 | x4) & (~x1 | (x2 ? (~x3 | x4) : x3))));
  assign n6874 = ~n1134 & (n880 | (~x0 & (n676 | n979)));
  assign n6875 = n841 & ((x2 & (x3 ? ~x4 : (x4 & ~x5))) | (~x3 & ~x4 & x5) | (~x2 & (x3 ? (x4 & ~x5) : ~x4)));
  assign n6876 = ~x2 & (x1 ? (n6877 | n6880) : ~n6878);
  assign n6877 = n942 & n2204;
  assign n6878 = (~x6 | n6879) & (x0 | ~n1029 | ~n658);
  assign n6879 = (~x0 | ((x3 | ~x4 | ~x5 | ~x7) & (~x3 | x4 | x5 | x7))) & (x0 | x3 | ~x4 | ~x5 | x7);
  assign n6880 = ~n3754 & n653 & ~x6 & x7;
  assign n6881 = (~x0 & ((~x2 & x5) | (~x1 & (x5 ? ~x3 : x2)))) | (x2 & ((x0 & x3 & x5) | (x1 & ~x3 & ~x5))) | (x0 & (x1 | (~x2 & x3 & ~x5))) | (~x2 & (x3 ? x1 : x5));
  assign n6882 = ~n6883 & ~n6885 & ~n6886 & (~n1209 | ~n1621);
  assign n6883 = n742 & ((n942 & n6073) | (n4972 & ~n6884));
  assign n6884 = (~x1 | ~x5 | (~x3 ^ x6)) & (x5 | x6 | x1 | ~x3);
  assign n6885 = ~n2128 & (x0 ? (x1 ? (~x2 & ~x3) : (x2 & x3)) : ((~x2 & x3) | (~x1 & x2 & ~x3)));
  assign n6886 = ~x0 & (n6887 | (~x1 & n1518 & n943));
  assign n6887 = ~x7 & x6 & ~x5 & x1 & ~x4;
  assign z388 = n6898 | ~n6903 | (x5 ? ~n6894 : ~n6889);
  assign n6889 = (x1 | n6890) & (x0 | ~x1 | n6893);
  assign n6890 = (~x6 | x7 | ~n1029 | n6891) & (~x7 | n6892);
  assign n6891 = ~x0 & x2;
  assign n6892 = (x0 | x2 | x3 | x4 | ~x6) & (x6 | ((x3 | ~x4 | (x0 & ~x2)) & (~x0 | x4 | (~x2 ^ ~x3))));
  assign n6893 = (~x2 | ~x3 | x4 | ~x6 | x7) & (x3 | (x2 ? (x4 ? (~x6 | x7) : (x6 | ~x7)) : (x7 | (x4 & x6))));
  assign n6894 = ~n6897 & (x3 | (~n6896 & (~x4 | n6895)));
  assign n6895 = x0 ? (x7 | (x1 ? (x2 | ~x6) : (~x2 | x6))) : (~x1 | ~x7 | (~x2 & x6));
  assign n6896 = ~x4 & n1181 & (x1 ? x7 : (x6 & ~x7));
  assign n6897 = n6063 & (x1 ? ~x7 : (~x2 & x7));
  assign n6898 = ~n640 & (~n6900 | (~x0 & ~n6899));
  assign n6899 = (x1 | x2 | x3 | ~x4) & (~x5 | ((x1 | x2 | ~x3 | x4) & (~x1 | (x2 ? (x3 | x4) : (~x3 | ~x4)))));
  assign n6900 = ~n6901 & ~n6902 & (~n560 | ~n639);
  assign n6901 = ~x5 & (x1 ? (x0 ? (~x2 & ~x3) : x3) : (x2 & ~x3));
  assign n6902 = ~x1 & x5 & ((x2 & x3) | (x0 & ~x2 & ~x3));
  assign n6903 = ~n6905 & (n3315 | n6904);
  assign n6904 = (x2 | ((x0 | ~x1 | ~x4 | x5) & (~x0 | (x1 ? (x4 | x5) : ~x5)))) & (x1 | ((~x4 | ~x5) & (x4 | x5 | x0 | ~x2)));
  assign n6905 = ~n643 & ((~n2373 & ~n1148) | (~x4 & ~n6906));
  assign n6906 = (x0 | ~x1 | x2 | ~x3 | ~x5) & (x1 | (x2 ? (x3 | ~x5) : (~x3 | x5)));
  assign z389 = n6914 | ~n6920 | (x6 ? ~n6916 : ~n6908);
  assign n6908 = x1 ? n6911 : (~n6910 & (~x5 | n6909));
  assign n6909 = (x4 | (x0 ? (x2 ? (x3 | ~x7) : (~x3 | x7)) : (x2 ? (x3 | x7) : (~x3 | ~x7)))) & (~x0 | ~x4 | (x2 ? (~x3 | x7) : x3));
  assign n6910 = n757 & ((~x0 & x2 & (x3 ^ ~x4)) | (~x2 & ((x3 & ~x4) | (x0 & ~x3 & x4))));
  assign n6911 = (x2 | n6913) & (x0 | ~x2 | n6912);
  assign n6912 = (x3 | x4 | ~x5 | x7) & (~x3 | ~x4 | (~x5 ^ x7));
  assign n6913 = (~x4 | ((x0 | ~x3 | x5 | x7) & (~x0 | x3 | (x5 & x7)))) & (x0 | ~x3 | x4 | (~x5 & ~x7));
  assign n6914 = x4 & ((n804 & n2862) | (x2 & ~n6915));
  assign n6915 = (x0 | ((~x6 | ~x7 | ~x1 | ~x5) & (x6 | x7 | (x1 & x5)))) & (x1 | ((~x0 | ~x6 | ~x7) & (x5 | (~x6 ^ ~x7))));
  assign n6916 = ~n6919 & (x2 | (~x1 & n6917) | (x1 & n6918));
  assign n6917 = (~x0 | x4 | ~x5 | (~x3 ^ ~x7)) & (~x4 | ((~x3 | x5 | ~x7) & (x0 | (x3 ? ~x7 : (x5 | x7)))));
  assign n6918 = (x0 | x7 | (x3 ? (~x4 | x5) : (x4 | ~x5))) & (~x0 | x3 | ~x4 | ~x7);
  assign n6919 = n4240 & ((x4 & x7 & ~x0 & x3) | (~x3 & ((x4 & ~x7) | (x0 & ~x4 & x7))));
  assign n6920 = n6923 & (n1116 | n6921) & (n1008 | n6922);
  assign n6921 = (x0 | ((~x1 | x2 | x3) & (~x2 | x4))) & (x4 | ((x1 | ~x2 | ~x3) & (~x0 | x2 | x3)));
  assign n6922 = (~x2 | x4 | x6 | ~x0 | x1) & (x0 | ~x1 | ~x4 | ~x6);
  assign n6923 = (n6924 | n6925) & (~n1167 | n6926);
  assign n6924 = x0 ? (~x3 | x7) : (x3 | ~x7);
  assign n6925 = (~x1 | x2 | x4 | x5 | ~x6) & (x1 | ((~x5 | ~x6 | ~x2 | ~x4) & (x2 | x5 | (~x4 ^ ~x6))));
  assign n6926 = (~x1 | ~x2 | x5 | x6 | ~x7) & (x2 | ~x5 | ((~x6 | ~x7) & (x1 | x6 | x7)));
  assign z390 = n6932 | ~n6935 | (x7 & (n6928 | n6930));
  assign n6928 = ~n6929 & ~x1 & ~n1134;
  assign n6929 = x0 ? (x2 ? (x3 | ~x6) : (~x3 | x6)) : (x2 | (~x3 ^ ~x6));
  assign n6930 = x1 & (x0 ? (n902 & n696) : ~n6931);
  assign n6931 = (~x2 | x3 | x4 | ~x5 | ~x6) & (x2 | ((~x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (x3 | ~x4 | x5 | x6)));
  assign n6932 = ~n765 & (x1 ? ~n6933 : ~n6934);
  assign n6933 = (x2 | ((~x4 | x6 | x0 | ~x3) & (x4 | ~x6 | ~x0 | x3))) & (x0 | ~x2 | (x6 ? (~x3 & ~x4) : x3));
  assign n6934 = (x0 | (x2 ? (x3 | ~x6) : (~x3 | x6))) & (~x2 | ((~x0 | x4 | x6) & ((~x3 ^ ~x6) | (~x0 & x4))));
  assign n6935 = ~n6940 & n6942 & (n1008 | (~n6936 & n6937));
  assign n6936 = n543 & ((~x2 & ~x4 & (x3 ^ ~x6)) | (x2 & x3 & x4 & ~x6));
  assign n6937 = ~n6938 & ~n6939 & (~n560 | ~n2352);
  assign n6938 = ~x2 & (x0 ? ((~x3 & ~x6) | (~x1 & x3 & x6)) : (~x3 & x6));
  assign n6939 = ~x6 & x3 & x2 & ~x0 & ~x1;
  assign n6940 = ~x2 & ((n592 & n727) | (~x3 & ~n6941));
  assign n6941 = (x0 | x1 | ~x4 | x5 | x6) & (~x0 | ~x5 | ~x6 | (~x1 ^ ~x4));
  assign n6942 = (n1580 | n6943) & (~x4 | ~n1885 | ~n2431);
  assign n6943 = (x5 | x6 | x2 | ~x3) & (~x2 | (x3 ? (~x5 | x6) : (x5 | ~x6)));
  assign z391 = n6953 | ~n6957 | (x2 ? ~n6945 : ~n6948);
  assign n6945 = ~n6946 & (~n659 | (~n936 & (x0 | n1820)));
  assign n6946 = x5 & ((n866 & n2834) | (~x1 & ~n6947));
  assign n6947 = x0 ? ((~x6 | ~x7 | ~x3 | ~x4) & (x6 | x7 | x3 | x4)) : (x3 | (x4 ? (x6 | x7) : (~x6 | ~x7)));
  assign n6948 = x4 ? n6951 : (~n6950 & (~n689 | ~n6949));
  assign n6949 = ~x5 & (x0 ? (~x6 & ~x7) : (x6 & x7));
  assign n6950 = ~n640 & ((n1301 & n841) | (~x0 & ~n1221));
  assign n6951 = x5 ? (~n1857 | ~n699) : n6952;
  assign n6952 = (~x0 | ((x1 | ~x3 | ~x6 | ~x7) & (~x1 | x3 | x6 | x7))) & (x0 | x1 | x3 | x6 | x7);
  assign n6953 = ~n643 & (n6955 | ~n6956 | (~x2 & ~n6954));
  assign n6954 = (x0 | ~x3 | ~x5 | (~x1 ^ ~x4)) & (x5 | ((x0 | x1 | ~x3 | ~x4) & (~x0 | (x1 ? (~x3 | x4) : (x3 | ~x4)))));
  assign n6955 = x2 & ((~x3 & x4 & x0 & ~x1) | (~x0 & (x1 ? (~x3 & ~x4) : (x3 & x4))));
  assign n6956 = (~n1209 | ~n1311) & (x3 | ~n743 | n1164);
  assign n6957 = ~n6958 & n6960 & ~n6963 & (x1 | n6962);
  assign n6958 = ~n5269 & ~n6959;
  assign n6959 = (x0 | ~x1 | ~x2 | x4 | ~x5) & (~x4 | ((x0 | ~x1 | x2 | ~x5) & (~x0 | x1 | (~x2 ^ ~x5))));
  assign n6960 = (x4 | n6961) & (~x2 | ~x4 | ~n543 | n627);
  assign n6961 = x0 ? ((x1 | ~x2 | ~x3 | ~x6) & (~x1 | x2 | x3 | x6)) : ((x1 | ~x2 | ~x3 | x6) & (~x1 | x2 | x3 | ~x6));
  assign n6962 = x0 ? ((x6 | n646) & (x2 | ~x6 | n647)) : ((~x6 | n646) & (x2 | x6 | n647));
  assign n6963 = n1283 & (n960 | (x3 & n6964));
  assign n6964 = ~x6 & (x4 ^ x5);
  assign z392 = n6966 | ~n4489 | (~x0 & x1 & ~n668);
  assign n6966 = ~x3 & ((~n1218 & ~n4488) | (n527 & ~n6967));
  assign n6967 = (x0 | x2 | ~x4 | x5 | x7) & (~x0 | ~x2 | x4 | ~x5 | ~x7);
  assign z393 = n6976 | n6972 | n4504 | n6969;
  assign n6969 = ~x2 & (n3181 | ~n6971 | (x5 & ~n6970));
  assign n6970 = (~x0 | x1 | x3 | ~x4 | ~x6) & (x6 | ((x1 | ~x3 | x4) & (x0 | ((~x3 | x4) & (~x1 | x3 | ~x4)))));
  assign n6971 = (~n704 | ~n699) & (~x6 | ~n1301 | n710);
  assign n6972 = ~x6 & (n6973 | n6975 | (n837 & n1598));
  assign n6973 = ~x7 & ((n733 & n1311) | (~x1 & ~n6974));
  assign n6974 = (x0 | ~x2 | x3 | x4 | x5) & (~x0 | ~x3 | ~x4 | (~x2 ^ ~x5));
  assign n6975 = ~n1920 & ((~x1 & ~x2 & x7) | (~x0 & ((~x2 & x7) | (x1 & x2 & ~x7))));
  assign n6976 = x6 & ((n4413 & n1269) | (n1392 & ~n6977));
  assign n6977 = x2 ? ((x0 | ~x5 | ~x7) & (x1 | ((~x5 | ~x7) & (~x0 | x5 | x7)))) : ((~x1 | ~x5 | x7) & (x0 | ((~x5 | x7) & (~x1 | x5 | ~x7))));
  assign z394 = n6979 | ~n6984 | ~n6991 | (~n1138 & ~n6990);
  assign n6979 = x4 & (n6980 | (n1451 & ~n6983));
  assign n6980 = x5 & ((x6 & ~n6981) | (n527 & ~n6982));
  assign n6981 = (x1 | ((x2 | ~x3 | x7) & (x3 | ~x7 | ~x0 | ~x2))) & (x0 | ~x1 | x3 | ~x7);
  assign n6982 = (x0 | x2 | ~x3 | ~x7) & (x3 | x7 | ~x0 | ~x2);
  assign n6983 = (~x2 | x6 | x7 | ~x0 | x1) & (x0 | ~x1 | x2 | (~x6 ^ ~x7));
  assign n6984 = ~n6985 & ~n6987 & ~n6989 & (n524 | n6986);
  assign n6985 = ~n3234 & ((~x0 & x1 & ~x4 & x5) | (~x1 & ((x4 & ~x5) | (x0 & ~x4 & x5))));
  assign n6986 = (x0 | x1 | ~x2 | ~x3 | ~x6) & (x3 | x6 | ((~x1 | x2) & (x0 | (~x1 & x2))));
  assign n6987 = ~n5496 & ~n6988;
  assign n6988 = (~x1 | x2 | x3 | ~x5 | ~x7) & (x1 | ((~x3 | x5 | x7) & (~x2 | (x3 ? x7 : (x5 | ~x7)))));
  assign n6989 = ~n4587 & ((x3 & x4 & x5) | (~x2 & (x3 ? x4 : (~x4 & ~x5))));
  assign n6990 = (~x0 | x2 | x4 | x5 | x7) & (x0 | ((~x4 | ~x5 | ~x7) & (~x2 | x4 | x5 | x7)));
  assign n6991 = x0 ? n6995 : (n6993 & (~x2 | n6992));
  assign n6992 = (x1 | ~x3 | ~x4 | ~x5 | x6) & (~x1 | x5 | (x3 ? (~x4 | x6) : (x4 | ~x6)));
  assign n6993 = (n714 | n1143) & (~n1084 | n6994);
  assign n6994 = (x5 | x6 | ~x1 | ~x3) & (x1 | x3 | ~x6);
  assign n6995 = x4 ? (~n1723 | ~n576) : n6996;
  assign n6996 = (x2 | (x1 ? (x3 | ~x6) : (~x3 | x6))) & (x1 | ((~x3 | x5 | x6) & (~x2 | x3 | ~x6)));
  assign z395 = n7006 | ~n7008 | (x1 ? ~n7003 : ~n6998);
  assign n6998 = x3 ? n6999 : (~n7001 & (~n658 | ~n3176));
  assign n6999 = (x4 | n7000) & (n640 | n791 | ~x2 | ~x4);
  assign n7000 = (x0 | x6 | ~x7 | (~x2 ^ ~x5)) & (~x6 | ((x0 | ~x2 | ~x5 | x7) & (~x0 | (x2 ? (x5 | x7) : (~x5 | ~x7)))));
  assign n7001 = ~x2 & ((n1310 & ~n4773) | (x0 & n7002));
  assign n7002 = x5 & (x4 ? ~x6 : (x6 & ~x7));
  assign n7003 = ~n7004 & (~n547 | ~n1725);
  assign n7004 = ~x5 & ((n3261 & ~n917) | (~x6 & ~n7005));
  assign n7005 = (x4 | ~x7 | ~x0 | x2) & (x0 | ((x2 | ~x3 | ~x4 | x7) & (~x2 | x4 | ~x7)));
  assign n7006 = ~x5 & ((n543 & n5758) | (~x1 & ~n7007));
  assign n7007 = x0 ? (x2 | x3 | (~x4 ^ x7)) : (~x2 | ((x4 | ~x7) & (~x3 | ~x4 | x7)));
  assign n7008 = ~n7010 & (~n5802 | ~n733) & (n1218 | n7009);
  assign n7009 = (~x0 | x1 | ~x2 | x3) & (~x3 | ((x0 | ~x1 | x2 | ~x5) & (~x0 | x1 | (x2 & ~x5))));
  assign n7010 = ~n1176 & (n880 | (~x0 & (n676 | ~n3802)));
  assign z396 = n7020 | ~n7022 | (x5 ? ~n7012 : ~n7015);
  assign n7012 = ~n7013 & (~n1300 | ~n1029 | ~n560);
  assign n7013 = ~x3 & ((n560 & n1585) | (~x6 & ~n7014));
  assign n7014 = (x0 | ~x1 | x2 | x4 | x7) & (x1 | ((~x4 | x7 | x0 | ~x2) & (~x0 | (x2 ? (x4 | x7) : (~x4 | ~x7)))));
  assign n7015 = x4 ? n7018 : (~n7017 & (x6 | n7016));
  assign n7016 = x0 ? (x2 | (x1 ? ~x3 : (x3 | x7))) : (x1 | ~x2 | (~x3 ^ ~x7));
  assign n7017 = n778 & ((n543 & n1465) | (n536 & ~n1543));
  assign n7018 = (~x6 | n7019) & (x3 | x6 | x7 | ~n816);
  assign n7019 = (~x0 | ~x1 | x2 | x3 | x7) & (x0 | ~x3 | ~x7 | (~x1 ^ ~x2));
  assign n7020 = ~x1 & ((n594 & n978) | (n1051 & ~n7021));
  assign n7021 = (x0 | x5 | ~x7) & (x2 | ((x5 | ~x7) & (~x0 | ~x5 | x7)));
  assign n7022 = ~n7023 & ~n7026 & n7027 & (x1 | n7025);
  assign n7023 = ~n714 & ((n1209 & n684) | (~x0 & ~n7024));
  assign n7024 = (~x1 | ((~x2 | x3 | ~x6 | x7) & (x2 | ~x3 | x6 | ~x7))) & (x1 | x2 | x3 | ~x6 | x7);
  assign n7025 = (x0 | ~x2 | ~x3 | ~x5 | x6) & (x2 | ((~x0 | (x3 ? (~x5 | x6) : (x5 | ~x6))) & (x5 | x6 | x0 | ~x3)));
  assign n7026 = ~n3924 & ((x0 & ~x1 & x2 & ~x6) | (~x0 & (x1 ? (x2 ^ ~x6) : (~x2 & x6))));
  assign n7027 = ~n7028 & ~n7029 & (~n837 | (~n3848 & ~n2904));
  assign n7028 = ~x0 & ((x1 & (x2 ? (~x5 & ~x6) : (x5 & x6))) | (~x1 & x2 & ~x5 & x6));
  assign n7029 = x6 & x5 & x2 & x0 & ~x1;
  assign z397 = n7031 | ~n7039 | ~n7044 | (~n643 & ~n7036);
  assign n7031 = ~x1 & (n7032 | (~x0 & (n2384 | n7035)));
  assign n7032 = x0 & (x2 ? (n7033 | n7034) : n4449);
  assign n7033 = x7 & x6 & ~x5 & ~x3 & x4;
  assign n7034 = ~x7 & ~x6 & x5 & x3 & ~x4;
  assign n7035 = n4089 & (x2 ? (~x3 & n1364) : (n3848 | (x3 & n1364)));
  assign n7036 = ~n7037 & n7038 & (~n743 | n2208 | n1566);
  assign n7037 = ~x2 & ((~x1 & x3 & ~x4) | (~x3 & (x0 ? (x1 & x4) : (~x1 ^ ~x4))));
  assign n7038 = (~n1716 | ~n746) & (~n543 | ~n1489);
  assign n7039 = (n640 | n7040) & (~n4248 | n7043);
  assign n7040 = x0 ? (x1 | (~n7041 & ~n2537)) : n7042;
  assign n7041 = ~x2 & ~x3 & (x4 ^ x5);
  assign n7042 = x1 ? (x2 | (x3 ? x4 : (~x4 | ~x5))) : (~x2 | (x3 ? (x4 | x5) : ~x4));
  assign n7043 = (x0 | ~x4 | x5 | ~x6 | ~x7) & (x4 | ((x6 | x7 | ~x0 | ~x5) & (x0 | (x5 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n7044 = x1 ? n7047 : (x6 ? n7045 : n7046);
  assign n7045 = (x2 | ~x3 | ~x4 | (x0 & ~x5)) & (x3 | x4 | ((~x2 | x5) & (~x0 | (~x2 & x5))));
  assign n7046 = (~x2 | ~x3 | ~x4) & (x0 | ~x5 | (x2 ? ~x3 : (x3 | x4)));
  assign n7047 = (~n696 | ~n600) & (x0 | n7048);
  assign n7048 = (x4 | x6 | ~x2 | x3) & (~x3 | (x2 ? (~x6 | (~x4 & ~x5)) : (~x4 | x6)));
  assign z398 = n7050 | ~n7053 | n7058 | (x6 & ~n7060);
  assign n7050 = ~x1 & ((~x4 & ~n7051) | (n1121 & ~n7052));
  assign n7051 = (x0 | ~x2 | ~x3 | (~x5 ^ ~x7)) & (x3 | ((x0 | ~x2 | x5 | ~x7) & (~x0 | x2 | (~x5 ^ x7))));
  assign n7052 = (x3 | x7 | x0 | x2) & (~x0 | (x2 ? (x3 | x7) : (~x3 | ~x7)));
  assign n7053 = ~n7055 & n7057 & (x1 | n7054);
  assign n7054 = (x0 | x2 | x3 | x4 | ~x7) & (~x0 | ((~x3 | x4 | x7) & (~x2 | ~x7 | (~x3 ^ ~x4))));
  assign n7055 = ~x6 & ((n560 & n5969) | (n543 & ~n7056));
  assign n7056 = x2 ? (x4 | ~x5 | (x3 ^ ~x7)) : (x5 | (x3 ? (~x4 | x7) : ~x7));
  assign n7057 = (~x4 | ~x7 | x0 | ~x3) & (x7 | ((x3 | ~x4 | ~x0 | x2) & (x0 | (x2 ? (x3 | ~x4) : (~x3 | x4)))));
  assign n7058 = x1 & ((n674 & n547) | (~x4 & ~n7059));
  assign n7059 = (x0 | ~x5 | (x2 ? (~x3 | ~x7) : (x3 | x7))) & (x5 | (~x0 ^ x2) | (~x3 ^ x7));
  assign n7060 = ~n7062 & (x1 | (n7061 & (n882 | n5085)));
  assign n7061 = (~n809 | ~n1783) & (~n594 | ~n635);
  assign n7062 = n4248 & ((x0 & ~x4 & x5 & ~x7) | (~x0 & ((~x5 & ~x7) | (~x4 & x5 & x7))));
  assign z399 = ~n7075 | n7072 | n7064 | n7067;
  assign n7064 = ~x7 & ((n733 & n1643) | (~x1 & ~n7065));
  assign n7065 = (~x6 | n1548 | ~n1549) & (~x2 | n7066);
  assign n7066 = (~x0 | x3 | x4 | x5 | x6) & (x0 | ~x4 | (x3 ? (x5 | ~x6) : (~x5 | x6)));
  assign n7067 = x7 & (x0 ? ~n7070 : ~n7068);
  assign n7068 = x6 ? (~n2332 | n1480) : n7069;
  assign n7069 = x1 ? (~x3 | (x2 ? (x4 | ~x5) : (~x4 | x5))) : (x3 | (x2 ? (x4 | ~x5) : x5));
  assign n7070 = (~n706 | ~n1044 | ~x1 | x4) & (x1 | (~n7071 & (~x4 | ~n706 | ~n1044)));
  assign n7071 = x2 & ((x3 & ~x4 & x5 & x6) | (~x3 & x4 & ~x5 & ~x6));
  assign n7072 = ~x2 & ((x1 & ~n7073) | (n841 & ~n7074));
  assign n7073 = (x0 | ~x5 | (x3 ? (~x4 | ~x6) : (x4 | x6))) & (x3 | ~x4 | x5 | ~x6);
  assign n7074 = (x3 | x4 | ~x5 | x6) & (~x3 | (x4 ? ~x6 : (x5 | x6)));
  assign n7075 = n7078 & (x2 | n7076) & (n627 | n7077);
  assign n7076 = (x0 | ~x3 | ~x4 | x5 | ~x6) & (x3 | ((~x5 | x6 | x0 | ~x4) & (~x0 | (x4 ? (x5 | x6) : (~x5 | ~x6)))));
  assign n7077 = (x0 | ((x1 | ((~x2 | x4 | ~x5) & (~x4 | x5))) & (~x2 | ~x4 | x5) & (x2 | ((~x4 | ~x5) & (~x1 | x4 | x5))))) & (x1 | ~x4 | (x5 ? ~x0 : ~x2));
  assign n7078 = (~n859 | ~n1323) & (x0 | ~n7071);
  assign z400 = ~n7081 | ~n7086 | ~n7089 | (~n1097 & ~n7080);
  assign n7080 = x0 ? ((x1 | ~x2 | ~x3 | ~x4) & (~x1 | x2 | x3 | x4)) : ((~x3 | ~x4 | x1 | x2) & (~x2 | (x1 ? (~x3 ^ x4) : (x3 | x4))));
  assign n7081 = n7084 & ~n7082 & n7083;
  assign n7082 = ~x2 & ((n1716 & n626) | (x0 & n959));
  assign n7083 = (~n731 | ~n746) & (~n895 | n6433);
  assign n7084 = (~n1283 | n7085) & (~n2534 | ~n4900);
  assign n7085 = (x5 | ~x6) & (x3 | ~x5 | x6);
  assign n7086 = ~n7088 & (x1 | (~x0 & n3838) | (x0 & n7087));
  assign n7087 = (x2 | ~x3 | ~x5 | x6) & (x5 | ~x6 | ~x2 | x3);
  assign n7088 = x2 & ((n696 & n712) | (n653 & ~n1335));
  assign n7089 = n7093 & (~x2 | (~n7091 & (~n1365 | ~n7090)));
  assign n7090 = ~x4 & x6 & (x5 ^ ~x7);
  assign n7091 = ~x3 & (x0 ? (n1145 & n951) : ~n7092);
  assign n7092 = (x1 | ~x4 | ~x5 | x6 | ~x7) & (~x1 | x4 | x5 | ~x6 | x7);
  assign n7093 = (n1014 | n7094) & (n1337 | n7095);
  assign n7094 = (~x0 | ~x1 | x2 | x3 | x6) & (x0 | ((~x3 | ~x6 | x1 | x2) & (~x2 | (x1 ? (~x3 ^ x6) : (x3 | x6)))));
  assign n7095 = (x0 | ~x1 | x2 | ~x3 | x6) & (x1 | ((~x3 | ~x6 | x0 | ~x2) & (x3 | (x0 ? (~x2 ^ x6) : (x2 | x6)))));
  assign z401 = ~n7099 | n7105 | ~n7107 | (~x1 & ~n7097);
  assign n7097 = (x2 | n7098) & (x0 | ~x2 | ~x6 | n1920);
  assign n7098 = (x0 | ~x3 | ~x4 | ~x5 | ~x6) & (x3 | ((x5 | ~x6 | x0 | x4) & (~x0 | x6 | (~x4 ^ ~x5))));
  assign n7099 = ~n7100 & ~n7102 & n7104 & (~x6 | n7103);
  assign n7100 = ~n643 & (n5363 | (~n714 & (n880 | n7101)));
  assign n7101 = ~x0 & (x1 ^ ~x3);
  assign n7102 = ~n647 & ((x2 & x6 & ~x0 & x1) | (~x6 & (x0 ? (~x1 ^ ~x2) : (~x1 & ~x2))));
  assign n7103 = (~x3 | ~x4 | ~x0 | x1) & (x2 | x3 | x0 | ~x1);
  assign n7104 = (~n761 | ~n1269) & (~x4 | ~n658 | ~n1922);
  assign n7105 = ~n640 & (n7106 | (~n714 & (n935 | n2144)));
  assign n7106 = n1188 & ((~x0 & x2 & x4 & ~x5) | (x0 & ~x4 & (~x2 | x5)));
  assign n7107 = ~n7109 & (x5 | n7108) & (n615 | n7110);
  assign n7108 = (~n2359 | ~n1317 | n6389) & (~n3790 | ~n1365);
  assign n7109 = n3488 & ((n1121 & n902) | (x2 & ~n1920));
  assign n7110 = (~x0 | x1 | ~x2 | x5 | ~x7) & (x0 | ((x1 | ~x2 | ~x5 | ~x7) & (~x1 | x2 | x5 | x7)));
  assign z402 = n7112 | n7121 | n7125 | (~x5 & ~n7117);
  assign n7112 = ~x7 & (n7113 | n7114);
  assign n7113 = ~n752 & ((n841 & n2371) | (~x0 & ~n753));
  assign n7114 = ~x1 & (x0 ? ~n7115 : ~n7116);
  assign n7115 = (x5 | ~x6 | ~x3 | ~x4) & (x3 | ((x5 | x6 | ~x2 | x4) & (x2 | ~x5 | (~x4 ^ ~x6))));
  assign n7116 = (~x5 | ~x6 | ~x3 | ~x4) & (x3 | x4 | (x2 ? (~x5 | x6) : (x5 | ~x6)));
  assign n7117 = n7119 & (x2 ? (x0 | n1218) : n7118);
  assign n7118 = (~x0 | x1 | x3 | ~x4 | ~x7) & (x4 | ((x0 | ~x1 | x3 | x7) & (x1 | (x0 ? (~x3 ^ ~x7) : (~x3 | x7)))));
  assign n7119 = ~n7120 & (~n1209 | ~n2647);
  assign n7120 = ~x2 & ((~x0 & ~x1 & x4 & x7) | (x0 & x1 & ~x4 & ~x7));
  assign n7121 = x5 & (n7122 | n7124 | (~x0 & ~n7123));
  assign n7122 = n560 & n2647;
  assign n7123 = (x3 | x7 | ~x1 | x2) & (x1 | x4 | ~x7 | (x2 ^ ~x3));
  assign n7124 = ~n671 & (x0 ? (x1 ? n1044 : ~n2737) : (x1 ? ~n2737 : n1044));
  assign n7125 = x7 & (n7126 | (~n1408 & ~n3208));
  assign n7126 = ~x3 & (x2 ? ~n7127 : (n543 & ~n2259));
  assign n7127 = (~x4 | x5 | x6 | ~x0 | x1) & (x0 | ((x1 | ~x4 | ~x5 | x6) & (~x1 | x4 | x5 | ~x6)));
  assign z403 = ~n7129 | (~x6 & ~n7138) | (~x2 & ~n7140);
  assign n7129 = ~n7130 & n7134 & (n835 | n7133);
  assign n7130 = x6 & (x2 ? ~n7132 : ~n7131);
  assign n7131 = (~x0 | x5 | (x1 ? (x3 | ~x7) : ~x3)) & (~x5 | ((~x0 | ~x1 | x3 | x7) & (x0 | ((~x3 | x7) & (x1 | x3 | ~x7)))));
  assign n7132 = (~x5 | x7 | x0 | ~x3) & (x1 | ((~x5 | ~x7 | x0 | x3) & (~x0 | x5 | (~x3 ^ x7))));
  assign n7133 = x0 ? (x1 | (x2 ? (~x5 ^ x6) : (x5 | x6))) : ((~x1 | (x2 ? ~x5 : (x5 | ~x6))) & (~x2 | ~x5 | ~x6) & (x1 | (x2 ? (x5 | x6) : ~x5)));
  assign n7134 = (n7135 | n7136) & (~x7 | ~n596 | n7137);
  assign n7135 = (x5 | x6 | x2 | x4) & (~x5 | ~x6 | ~x2 | ~x4);
  assign n7136 = (~x0 | x1 | ~x3 | x7) & (x0 | ~x1 | x3 | ~x7);
  assign n7137 = (x0 | ~x1 | x4 | x5 | ~x6) & (x1 | x6 | (x0 ? (~x4 ^ ~x5) : (x4 | ~x5)));
  assign n7138 = (~x5 | n7139) & (x7 | ~n1269 | ~x3 | x5);
  assign n7139 = x0 ? (x1 ? (x2 | x3) : (~x3 | x7)) : ((~x1 | ((~x2 | x3 | ~x7) & (~x3 | x7))) & (x2 | (x1 ? ~x3 : (x3 | ~x7))));
  assign n7140 = ~n7142 & (x3 | (~n7141 & (~n841 | ~n3853)));
  assign n7141 = n543 & (n588 | (x4 & (n706 | n1070)));
  assign n7142 = ~n7143 & ~x7 & n825;
  assign n7143 = (x5 | ~x6 | ~x1 | x4) & (x1 | x6 | (x4 ^ ~x5));
  assign z404 = n7145 | n7147 | ~n7152 | (n876 & ~n7151);
  assign n7145 = n619 & (x0 ? ~n7146 : (n596 & n926));
  assign n7146 = x2 ? ((~x5 | ~x6 | ~x3 | ~x4) & (x3 | x4 | x6)) : (~x3 | x6 | (~x4 & ~x5));
  assign n7147 = ~x7 & ((~x5 & ~n7148) | (n551 & ~n7150));
  assign n7148 = x1 ? (x6 | n7149) : (~x6 | (~n600 & n4477));
  assign n7149 = (~x0 | x2 | ~x3 | x4) & (x0 | ~x2 | x3 | ~x4);
  assign n7150 = (x3 | x4 | ~x6 | (~x0 & ~x2)) & (x2 | ((~x3 | ~x6) & (x0 | x4 | x6)));
  assign n7151 = (x0 | ~x1 | x2 | x4 | ~x6) & (x1 | ((x2 | x4 | x6) & (~x4 | ~x6 | ~x0 | ~x2)));
  assign n7152 = ~n7153 & n7156 & (~x2 | n7155);
  assign n7153 = ~n7154 & (x1 ? (x6 ^ ~x7) : (~x6 & x7));
  assign n7154 = (x3 | (x0 ? x2 : x4)) & (x0 | x2 | (x4 ? ~x3 : ~x5));
  assign n7155 = (x1 | ~x6 | (~x3 ^ x4)) & (x0 | (x1 ? (~x3 | x6) : (~x4 | ~x6)));
  assign n7156 = (~n2021 | n1312) & (~n746 | ~n1759);
  assign z405 = ~n7163 | ~n7167 | (x7 ? ~n7158 : ~n7161);
  assign n7158 = ~n7160 & (~x3 | (~n7159 & (~n841 | ~n5627)));
  assign n7159 = x1 & ((n743 & n696) | (n742 & n559));
  assign n7160 = ~x6 & n653 & (n5526 | (x1 & ~n1934));
  assign n7161 = ~n3196 & (x1 | (~n7162 & (n1932 | n2184)));
  assign n7162 = x6 & n1392 & (x0 ? n691 : n2371);
  assign n7163 = ~n7164 & ~n7165 & n7166 & (~n733 | ~n1598);
  assign n7164 = n841 & (x3 ? (x2 ? (~x4 & ~x7) : (x4 & x7)) : (~x4 & x7));
  assign n7165 = ~x0 & ((x2 & ~x3 & ~x4 & x7) | (~x2 & x4 & (x3 ^ ~x7)));
  assign n7166 = (~x3 | x7 | x0 | ~x2) & (~x0 | ~x1 | x2 | x3 | ~x7);
  assign n7167 = ~n7169 & (x1 | (~n808 & (~n525 | ~n7168)));
  assign n7168 = ~x5 & (x2 ? (x3 & ~x7) : (~x3 & x7));
  assign n7169 = ~n710 & (x2 ? (~x3 & n674) : (x3 & n2705));
  assign z406 = n7171 | ~n7173 | n7178 | (n1301 & ~n7177);
  assign n7171 = x2 & ~n7172;
  assign n7172 = (~x3 | ((~x0 | x1 | ~x4 | x5) & (x0 | ~x5 | (~x1 ^ x4)))) & (~x0 | x1 | x4 | (x3 & ~x5));
  assign n7173 = n7176 & (x5 ? (~n825 | n7175) : n7174);
  assign n7174 = (x0 | ~x2 | x3 | ~x4 | x6) & (x2 | ((x3 | ~x4 | ~x6) & (x4 | x6 | ~x0 | ~x3)));
  assign n7175 = x1 ? (~x4 | ~x6 | (x2 ^ ~x7)) : (x4 | x6 | (~x2 ^ ~x7));
  assign n7176 = (~x4 | ~x5 | x2 | x3) & (x0 | ((x2 | ~x3 | x4 | x5) & (~x2 | (x3 ? (~x4 | x5) : x4))));
  assign n7177 = (x0 | ~x1 | ~x2 | ~x4 | x6) & (x1 | ((x4 | ~x6 | x0 | ~x2) & (~x0 | ~x4 | (~x2 ^ x6))));
  assign n7178 = n2061 & ((~x2 & ~n7179) | (~x1 & x2 & ~n1862));
  assign n7179 = (~x3 | x4 | ~x6 | x7) & (~x1 | x3 | ~x4 | x6 | ~x7);
  assign z407 = n7181 | n7183 | ~n7186 | (~x1 & ~n7185);
  assign n7181 = ~n1205 & (x4 ? (n1364 & n543) : ~n7182);
  assign n7182 = (x0 | x1 | ~x5 | x6) & (~x0 | x5 | ~x6 | (x1 ^ ~x2));
  assign n7183 = ~x6 & ((n3034 & n4873) | (~x2 & ~n7184));
  assign n7184 = (~n699 | ~n867) & (x5 | ~n525 | n5144);
  assign n7185 = (x0 | x3 | (x4 ? (x5 | x6) : (~x5 | ~x6))) & (~x3 | ((~x0 | x5 | (~x4 ^ ~x6)) & (~x4 | ~x5 | (x0 & x6))));
  assign n7186 = ~n7187 & n7188 & (~n543 | (~n2794 & ~n2145));
  assign n7187 = ~x6 & ((n746 & n1311) | (n1549 & ~n1820));
  assign n7188 = (~n830 | ~n2534) & (n7189 | (x4 & ~x6));
  assign n7189 = x0 ? (x3 | ~x5 | (x1 & x2)) : (~x3 | x5);
  assign z408 = n7194 | ~n7196 | (x5 & ~n7191);
  assign n7191 = x0 ? (~n804 | ~n4897) : (~n7192 & ~n7193);
  assign n7192 = ~n2737 & (x1 ? ~n2803 : ~n3098);
  assign n7193 = n1044 & ((n1857 & n4894) | (~x1 & ~n3098));
  assign n7194 = ~n640 & (x2 ? (n1477 & n841) : ~n7195);
  assign n7195 = (x0 | ~x1 | x3 | x4 | ~x5) & (~x0 | ~x4 | x5 | (x1 ^ ~x3));
  assign n7196 = ~n1758 & (n1408 | n7197) & (n643 | n7198);
  assign n7197 = (x2 | x3 | ((x1 | x5) & (~x0 | ~x1 | ~x5))) & (x0 | x5) & (~x0 | x1 | ~x5 | (~x2 & ~x3));
  assign n7198 = ~n7199 & (n1954 | n4758) & (~n1716 | ~n560);
  assign n7199 = ~x0 & x4 & x5 & (x1 ^ ~x2);
  assign z409 = n4618 | n7201 | ~n7204 | (x0 & ~n7203);
  assign n7201 = ~x2 & (n7202 | (~x3 & n543 & ~n1337));
  assign n7202 = x0 & ((n927 & n2209) | (n689 & n717));
  assign n7203 = (x1 | x2 | x3 | x5 | ~x7) & ((~x5 ^ ~x7) | (x1 ^ (~x2 & ~x3)));
  assign n7204 = (~n904 | ~n1044 | n2223) & (x0 | n7205);
  assign n7205 = x1 ? (x5 | ~x7 | (~x2 & ~x3)) : (~x5 | x7);
  assign z410 = ~n7209 | (n1044 & ~n7207) | (~x2 & ~n7208);
  assign n7207 = (x0 | ~x1 | ~x4 | x6 | ~x7) & (x7 | ((x4 | ~x6 | ~x0 | x1) & (x0 | (x1 ? (~x4 ^ ~x6) : (~x4 | x6)))));
  assign n7208 = (x1 | ~x3 | x6 | x7) & (~x1 | (x0 ? (x3 | x6) : (~x3 | (~x6 ^ x7))));
  assign n7209 = n7212 & (x2 | (~n7210 & (~n661 | ~n931)));
  assign n7210 = ~x4 & ((n658 & n1244) | (n1093 & ~n7211));
  assign n7211 = (~x0 | ~x3 | x6) & (x0 | x3 | ~x6 | ~x7);
  assign n7212 = (x0 | (x1 ? (~x2 | (~x6 ^ x7)) : (~x6 | ~x7))) & (x1 | x6 | (x7 ? ~x0 : ~x2));
  assign z411 = n5782 | ~n7215 | (n743 & (n7214 | n1253));
  assign n7214 = ~x7 & (x1 ^ x3);
  assign n7215 = (x0 | ~x7) & (x1 | ((x2 | ~x7 | ~n2647) & (~x0 | x7 | (~x2 & ~n2647))));
  assign z412 = ~n2877 | (n560 & n1268) | (n1586 & ~n7217);
  assign n7217 = (~x4 | x6 | x7 | ~x0 | x1) & (x0 | ~x1 | x4 | ~x6 | ~x7);
  assign z413 = ~x0 & ~n7219;
  assign n7219 = n7221 & (x5 | ~n828 | (n4460 & n7220));
  assign n7220 = (x1 | x2 | x6 | ~x7) & (~x1 | ~x2 | ~x6 | x7);
  assign n7221 = (x1 & x2) | (~x1 & ~x2 & ~x3 & ~x4 & ~x5);
  assign z414 = n7224 | ~n7225 | ~n7226 | (~x4 & ~n7223);
  assign n7223 = (~x0 | x1 | x2 | ~x3 | x5) & (x0 | x3 | ~x5 | (~x1 ^ ~x2));
  assign n7224 = ~x0 & (x1 ? (x2 & x3) : (x2 ^ x3));
  assign n7225 = x3 | ((x0 | ~x1 | ~x2 | ~x4) & (x1 | x2 | (~x0 & ~x4)));
  assign n7226 = (~n681 | ~n626 | n3234) & (n4282 | ~n7227);
  assign n7227 = x7 & ~x5 & ~x4 & ~x0 & ~x3;
  assign z415 = n7232 | ~n7234 | (~x4 & (~n7229 | ~n7231));
  assign n7229 = x0 ? (~n804 | ~n3848) : n7230;
  assign n7230 = (~x1 | x2 | x3 | ~x5 | x6) & (x1 | x5 | (x2 ? (~x3 | ~x6) : (~x3 ^ x6)));
  assign n7231 = (x0 | ~x1 | x3 | (~x2 ^ ~x5)) & (x1 | ((x3 | ~x5 | x0 | x2) & (~x3 | (x0 ? (~x2 ^ x5) : (~x2 | ~x5)))));
  assign n7232 = n828 & ((n560 & n942) | (~x0 & ~n7233));
  assign n7233 = (x1 | x2 | x5 | x6 | ~x7) & (~x1 | ~x6 | (x2 ? (x5 | ~x7) : (~x5 | x7)));
  assign n7234 = (x0 | ~x2 | ((~x3 | ~x4) & (~x1 | (~x3 & ~x4)))) & (x1 | ((x3 | ~x4 | x0 | x2) & (~x0 | (x2 ? x3 : (~x3 | ~x4)))));
  assign z416 = ~n7239 | (~x2 & ~n7236) | (x4 & ~n7238);
  assign n7236 = (~n830 | ~n866) & (x3 | (~n528 & ~n7237));
  assign n7237 = ~x1 & ((n951 & n1167) | (x0 & ~n990));
  assign n7238 = (x0 | ~x1 | x3) & (x1 | ((~x0 | ((~x3 | ~x5) & (x2 | x3 | x5))) & (~x3 | (x5 ? x2 : (x0 & ~x2)))));
  assign n7239 = ~n7241 & n7242 & (x5 | ~n1167 | n7240);
  assign n7240 = (x1 | ~x3 | ~x6) & (x6 | (x1 ^ (~x2 | x3)));
  assign n7241 = n1145 & ((~x3 & ~x5 & n995) | (x5 & (x3 | n600)));
  assign n7242 = (n2528 | n2267) & (~n543 | ~n1156 | ~n3709);
  assign z417 = n7244 | ~n7248 | (n1723 & ~n7247);
  assign n7244 = ~x2 & (n7245 | (n699 & n830));
  assign n7245 = x0 & ((~x5 & ~n7246) | (x1 & n1311));
  assign n7246 = x1 ? (x3 | ~x4) : (~x6 | ~x7 | (~x3 ^ ~x4));
  assign n7247 = (~x0 | x1 | x2 | ~x4 | x7) & (x0 | ~x1 | (~x4 ^ x7));
  assign n7248 = n7249 & (n710 | (~n2332 & ~n926));
  assign n7249 = ~n1723 | (x4 ? ~n1209 : ~n626);
  assign z418 = n7251 | n7254 | ~n7255 | (n608 & ~n7253);
  assign n7251 = ~x2 & (x0 ? ~n7252 : (n978 & n927));
  assign n7252 = x1 ? (x3 | ~x5) : (~x6 | ~x7 | (~x3 ^ ~x5));
  assign n7253 = (~x0 | x1 | ~x4 | ~x5 | ~x7) & (x0 | ~x1 | x7 | (~x4 ^ ~x5));
  assign n7254 = ~x0 & ((x5 & ~x6) | (~x1 & ~x5 & x6));
  assign n7255 = ~n2955 & ~n7256 & (~x6 | ~n1966 | n3134);
  assign n7256 = x6 & ((~x0 & x1 & ~x5 & x7) | (x0 & ~x1 & x5 & ~x7));
  assign z419 = n7258 | n7260 | ~n7261 | (~n640 & ~n2877);
  assign n7258 = n743 & ((n943 & n944) | (~x5 & ~n7259));
  assign n7259 = (x1 | x3 | ~x4 | ~x6 | ~x7) & (x4 | x6 | ~x1 | ~x3);
  assign n7260 = ~x1 & (x0 ? (~x6 & (x2 | x3)) : x6);
  assign n7261 = ~n1923 & (~n744 | ~n733) & (~n560 | ~n1525);
  assign z429 = ~x2 & (n7264 | ~n7265 | (~x1 & ~n7263));
  assign n7263 = (~x0 & (x3 | (x4 & x5 & x6))) | (x4 & ((x3 & x5) | (x0 & ~x5 & x6))) | (~x3 & ((~x4 & ~x5 & ~x6) | (x0 & (~x4 | ~x6))));
  assign n7264 = ~x1 & ((n5168 & n951) | (n525 & ~n2780));
  assign n7265 = ~n533 & (~n543 | ~n7266);
  assign n7266 = ~x4 & x5 & (x3 ? (~x6 & ~x7) : (x6 & x7));
  assign z430 = n7271 | ~n7268 | n7270;
  assign n7268 = ~n540 & n7269 & (~n543 | n544);
  assign n7269 = (~n931 | ~n5198) & (~n1364 | ~n774 | ~n733);
  assign n7270 = ~x1 & ((~n538 & n539) | (n549 & n728));
  assign n7271 = x3 & (n7272 | (n543 & n1835 & ~n2504));
  assign n7272 = n5260 & ((n757 & n1518) | (n750 & n1156));
  assign z431 = ~n7280 | (x0 ? (n7277 | n7279) : ~n7274);
  assign n7274 = ~n7275 & (~n979 | ~n1725);
  assign n7275 = x2 & ((n978 & n1288) | (~x5 & ~n7276));
  assign n7276 = x1 ? (x4 | (x3 ? (x6 | ~x7) : (~x6 | x7))) : (~x4 | (x3 ? (x6 | x7) : (~x6 | ~x7)));
  assign n7277 = ~x1 & ((n1562 & n1070) | (x2 & ~n7278));
  assign n7278 = (x3 | ~x4 | x5 | x6 | x7) & (~x3 | x4 | ~x5 | ~x6 | ~x7);
  assign n7279 = n576 & n993;
  assign n7280 = (~x1 | n7283) & (x1 | n554) & (x0 | n7281);
  assign n7281 = (~x5 | n7282) & (x4 | x5 | ~n1133 | n1026);
  assign n7282 = (x1 | x2 | x3 | ~x4 | ~x6) & (~x1 | ~x3 | (x2 ? (~x4 | x6) : (x4 | ~x6)));
  assign n7283 = (x2 | ((x4 | x5 | ~x0 | x3) & (x0 | ~x3 | ~x4))) & (x0 | ~x3 | ((~x4 | x5) & (~x2 | x4 | ~x5)));
  assign z432 = ~n7293 | ~n7290 | n7285 | n7288;
  assign n7285 = ~x0 & (n7287 | (~n627 & ~n7286));
  assign n7286 = (x1 | ~x2 | ~x4 | x5 | ~x7) & (x4 | ((x1 | x2 | ~x5 | x7) & (~x1 | ~x7 | (~x2 ^ x5))));
  assign n7287 = x7 & ((n559 & n2135) | (n558 & n696));
  assign n7288 = n3637 & ((n576 & n728) | (~x1 & ~n7289));
  assign n7289 = x2 ? ((~x3 | x4 | ~x5 | ~x6) & (x3 | ~x4 | x5 | x6)) : (~x4 | (x3 ? (x5 | ~x6) : (~x5 | x6)));
  assign n7290 = ~n7291 & (~n1268 | ~n837) & (x1 | n7292);
  assign n7291 = ~x5 & n626 & (n5787 | (x2 & n5072));
  assign n7292 = x2 ? ((x4 | x5 | x0 | x3) & (~x0 | ~x4 | (~x3 ^ x5))) : (~x3 | ((~x4 | ~x5) & (x0 | x4 | x5)));
  assign n7293 = n5806 & ~n7294 & (n968 | n7295);
  assign n7294 = x5 & ((n762 & n3828) | (x0 & ~n5809));
  assign n7295 = (x0 | ~x1 | ~x3 | x4 | ~x6) & (x3 | ((x0 | ~x1 | ~x4 | x6) & (~x0 | x1 | (~x4 ^ ~x6))));
  assign z433 = n7297 | n7301 | ~n7307 | (n543 & ~n7306);
  assign n7297 = ~x4 & (n7298 | (n742 & ~n627 & ~n2864));
  assign n7298 = ~x2 & ((x6 & ~n7299) | (n3074 & ~n7300));
  assign n7299 = (x0 | ~x1 | x3 | ~x5 | ~x7) & (x7 | ((x3 | x5 | x0 | ~x1) & (~x0 | x1 | (~x3 ^ ~x5))));
  assign n7300 = (x1 | x3 | x5 | ~x7) & (~x1 | ~x3 | (~x5 ^ ~x7));
  assign n7301 = x4 & (x2 ? ~n7303 : (n7302 | n7305));
  assign n7302 = n978 & n866;
  assign n7303 = (x1 | n7304) & (x0 | ~x1 | ~x5 | n3427);
  assign n7304 = (x0 | ~x3 | x5 | x6 | ~x7) & (x3 | ((~x6 | ~x7 | x0 | x5) & (~x0 | x6 | (~x5 ^ x7))));
  assign n7305 = n841 & ((n1769 & n3151) | (x3 & n881));
  assign n7306 = x4 ? ((x5 | ~x6 | ~x2 | x3) & (x2 | ~x3 | ~x5 | x6)) : (x2 ? (x3 ? (x5 | ~x6) : (~x5 | x6)) : (x3 ? (~x5 | ~x6) : (x5 | x6)));
  assign n7307 = ~n7308 & ~n7312 & n7313 & (x1 | n7310);
  assign n7308 = ~n1097 & ~n7309;
  assign n7309 = (~x0 | ((x1 | ~x2 | ~x3 | ~x4) & (x2 | x3 | x4))) & (x2 | ((x1 | x3 | ~x4) & (x0 | ((x3 | ~x4) & (x1 | ~x3 | x4)))));
  assign n7310 = (~n828 | n7311) & (x0 | ~n629) & (~x0 | n7087);
  assign n7311 = (x0 | x2 | x5 | ~x6) & (~x0 | ~x2 | ~x5 | x6);
  assign n7312 = ~n1014 & (n1675 | (~x2 & n626 & ~n627));
  assign n7313 = (n7314 | ~n2446) & (~x0 | n7315);
  assign n7314 = x1 ? (~x2 | x5) : (x2 | ~x5);
  assign n7315 = (x1 | ~x2 | ~x3 | x4 | x5) & (~x1 | x2 | x3 | ~x4 | ~x5);
  assign z434 = n7321 | ~n7323 | ~n7328 | (~x0 & ~n7317);
  assign n7317 = x1 ? n7319 : (~n7318 & (x2 | ~n5835));
  assign n7318 = ~x5 & (x2 ? (x3 & ~n1850) : (~x3 & n1395));
  assign n7319 = (~n658 | ~n1780) & (x2 | n7320);
  assign n7320 = (x3 | ~x6 | (x4 ? (~x5 | x7) : (x5 | ~x7))) & (~x3 | x4 | ~x5 | x6 | ~x7);
  assign n7321 = ~x5 & ((~n627 & ~n1961) | (~x4 & ~n7322));
  assign n7322 = (x0 | ~x1 | x2 | x3 | x6) & (x1 | ((x0 | (x2 ? (x3 | x6) : (~x3 | ~x6))) & (~x0 | x2 | ~x3 | x6)));
  assign n7323 = (~n841 | n7326) & (~x5 | (~n7324 & n7325));
  assign n7324 = ~n627 & ((~x2 & ~x4 & x0 & ~x1) | (~x0 & (x1 ? (x2 & ~x4) : x4)));
  assign n7325 = (~n3575 | ~n816) & (~n525 | n1009);
  assign n7326 = (~x6 | n7327) & (~x2 | ~x4 | ~n719);
  assign n7327 = (~x2 | x3 | x4 | ~x5 | x7) & (x2 | ((~x3 | x4 | ~x5 | ~x7) & (x3 | ~x4 | x5 | x7)));
  assign n7328 = ~n7329 & (n640 | (n7333 & (x0 | n7332)));
  assign n7329 = ~n643 & (x2 ? ~n7331 : ~n7330);
  assign n7330 = (x0 | ~x1 | ~x3 | x4 | x5) & (~x0 | x1 | x3 | ~x4 | ~x5) & ((x0 ? (~x1 | x3) : (x1 | ~x3)) | (~x4 ^ x5));
  assign n7331 = (~x0 | x1 | x3 | ~x4 | x5) & (x0 | ((~x1 | (x3 ? (x4 | x5) : (~x4 | ~x5))) & (x1 | ~x3 | x4 | ~x5)));
  assign n7332 = (x1 | x3 | ~x4 | x5) & (~x5 | ((x3 | x4 | x1 | ~x2) & (~x1 | x2 | (~x3 ^ ~x4))));
  assign n7333 = (n1920 | n1957) & (~n1365 | n7334);
  assign n7334 = (~x4 | x5) & (~x2 | x4 | ~x5);
  assign z435 = n7336 | ~n7339 | n7344 | (~x0 & ~n7346);
  assign n7336 = ~x5 & (x2 ? ~n7338 : ~n7337);
  assign n7337 = (x0 | x3 | ~x4 | (x1 ^ ~x7)) & (~x3 | ((x0 | ~x1 | x4 | ~x7) & (~x0 | ((x4 | x7) & (x1 | ~x4 | ~x7)))));
  assign n7338 = (x0 | ~x1 | x3 | x4 | ~x7) & (~x0 | x1 | ((~x4 | ~x7) & (x3 | x4 | x7)));
  assign n7339 = n7342 & (n765 | n7340) & (n1408 | n7341);
  assign n7340 = (~x0 | x2 | x3 | (x1 ^ ~x4)) & (x1 | ~x2 | ~x3 | x4) & (x0 | (~x2 & ~x3) | (~x1 ^ ~x4));
  assign n7341 = (~n1269 | ~n2476) & (~x5 | n2227 | n3134);
  assign n7342 = x5 ? (x7 | (n7343 & (x1 | n5194))) : (~x7 | n7343);
  assign n7343 = (~x0 | ~x1 | x2 | x3 | ~x4) & (x0 | ~x3 | (x1 ? (~x2 | x4) : (x2 | ~x4)));
  assign n7344 = ~n1353 & (x3 ? (n750 & n1209) : ~n7345);
  assign n7345 = (x0 | ~x1 | x2 | ~x5 | ~x7) & (x1 | ((~x0 | (x2 ? (~x5 | x7) : (x5 | ~x7))) & (x0 | x2 | ~x5 | x7)));
  assign n7346 = x1 ? (x2 | n7348) : (~n7347 & (x2 | ~n7266));
  assign n7347 = ~x5 & ((n1044 & n550) | (n859 & ~n871));
  assign n7348 = (x3 | x4 | x5 | ~x6 | ~x7) & (x6 | ((~x3 | x4 | ~x5 | ~x7) & (x3 | x7 | (~x4 ^ ~x5))));
  assign z436 = n7350 | n7353 | ~n7356 | (x5 & ~n7355);
  assign n7350 = ~x2 & (n7351 | (n828 & n7256));
  assign n7351 = ~x6 & ((n607 & n1922) | (~x3 & ~n7352));
  assign n7352 = (x4 | (x0 ? (x1 ? (x5 | x7) : (~x5 | ~x7)) : (x1 ? ~x5 : (x5 | ~x7)))) & (x0 | ~x4 | ((x1 | ~x5 | ~x7) & (x5 | (~x1 & x7))));
  assign n7353 = ~x1 & (n7354 | (x6 & n742 & ~n1558));
  assign n7354 = ~x2 & (x0 ? (~x3 & ~n1701) : (x3 & n943));
  assign n7355 = x0 ? (x1 ? (x2 | x3) : (~x2 | ~x6)) : ((~x2 | ~x3 | x6) & (x1 | (~x2 ^ x6)));
  assign n7356 = n7362 & ~n7361 & ~n7360 & ~n7357 & ~n7359;
  assign n7357 = ~n7358 & x6 & n742;
  assign n7358 = (~x1 | ~x3 | x4 | ~x5 | ~x7) & (x1 | ((x3 | ~x4 | x5 | ~x7) & (~x3 | x7 | (~x4 ^ x5))));
  assign n7359 = ~n3315 & (n5552 | (x2 & n681 & n841));
  assign n7360 = ~n1682 & ~n765 & ~n815;
  assign n7361 = ~n2227 & ((n1364 & n543) | (n904 & n841));
  assign n7362 = (~n3269 | ~n733) & (~n569 | ~n1301 | ~n746);
  assign z437 = ~n7373 | n7371 | n7364 | ~n7367;
  assign n7364 = ~n640 & ((n1145 & ~n7366) | (x4 & ~n7365));
  assign n7365 = (x0 | ~x1 | (x2 ? (~x3 | ~x5) : (x3 | x5))) & (x1 | (x0 ? (x2 | (~x3 & x5)) : (~x2 | x3)));
  assign n7366 = x0 ? (x5 ? x2 : x3) : (~x2 | ~x3);
  assign n7367 = (~n1621 | ~n3796) & (x2 | (~n7368 & n7369));
  assign n7368 = x1 & ((~n714 & ~n4925) | (~x0 & n744));
  assign n7369 = x0 ? (x6 | n647) : (x1 ? (~x6 | n647) : n7370);
  assign n7370 = (x3 | x4 | x5 | ~x6) & (~x3 | ~x4 | x6);
  assign n7371 = n1145 & ((n1693 & n943) | (x6 & ~n7372));
  assign n7372 = x0 ? (~x3 | x5 | (x2 ^ ~x7)) : (x3 | ~x5 | (~x2 ^ ~x7));
  assign n7373 = (n643 | n7377) & (~x2 | (~n7374 & n7375));
  assign n7374 = ~x0 & ((~x4 & ~x6 & x1 & x3) | (~x1 & (x3 ? (x4 & x6) : (~x4 & ~x6))));
  assign n7375 = ~n7376 & (~n577 | ~n661) & (~n926 | ~n866);
  assign n7376 = x6 & x4 & ~x3 & x0 & ~x1;
  assign n7377 = n7379 & (x4 ? (~n543 | n1916) : n7378);
  assign n7378 = (~x0 | ((x1 | ~x2 | ~x3 | ~x5) & (~x1 | x2 | x3 | x5))) & (x0 | x1 | x2 | ~x3 | x5);
  assign n7379 = (~x0 | x1 | ~x2 | ~x3 | ~x4) & (x0 | x3 | (x1 ? (~x2 | x4) : (x2 | ~x4)));
  assign z438 = ~n7387 | (x0 ? ~n7384 : ~n7381);
  assign n7381 = ~n1995 & (~x5 | (~n7382 & (x4 | n7383)));
  assign n7382 = ~n627 & ((n1133 & n1379) | (~x1 & n4089));
  assign n7383 = (~x1 | x2 | x3 | ~x6 | ~x7) & (x1 | x7 | ((x3 | x6) & (x2 | ~x3 | ~x6)));
  assign n7384 = ~n7386 & (x1 | (~n7385 & (~n978 | ~n2385)));
  assign n7385 = n681 & ((n902 & n1857) | (x7 & ~n5714));
  assign n7386 = n576 & n845;
  assign n7387 = ~n7389 & n7391 & (x1 | n7388);
  assign n7388 = (~x0 | x2 | x3 | x4 | ~x7) & (~x4 | (x0 ? ((~x3 | ~x7) & (~x2 | x3 | x7)) : (~x3 ^ x7)));
  assign n7389 = ~x7 & ((~n905 & n6127) | (~n1566 & ~n7390));
  assign n7390 = (x0 | ~x1 | x2 | ~x4) & (~x0 | x4 | (x1 ^ ~x2));
  assign n7391 = (~x1 | n7393) & (~x7 | (~n7392 & (x1 | n7394)));
  assign n7392 = ~x0 & x1 & x4 & (x3 ^ ~x5);
  assign n7393 = (x0 | ~x2 | x3 | x4 | ~x7) & (x7 | ((x3 | ~x4 | ~x0 | x2) & (x0 | x4 | (x2 & ~x3))));
  assign n7394 = (x4 | x5 | x0 | ~x3) & (~x0 | ((~x3 | x4 | ~x5) & (x2 | x3 | ~x4 | x5)));
  assign z439 = ~n5961 | n5970 | (x6 & n5966);
  assign z440 = n7403 | n7401 | n5981 | n7397;
  assign n7397 = ~x0 & (n7398 | (n2999 & n4248));
  assign n7398 = ~x7 & (x4 ? ~n7399 : (n1317 & ~n7400));
  assign n7399 = (x3 | ~x5 | ~x1 | x2) & (x1 | x5 | (x2 ? (~x3 | ~x6) : (x3 | x6)));
  assign n7400 = x2 ? (~x5 | x6) : x5;
  assign n7401 = ~x1 & (~n5979 | (~x7 & ~n7402));
  assign n7402 = x0 ? (x2 | (x3 ? (~x5 ^ x6) : (x5 | x6))) : ((~x2 | x3 | ~x5 | ~x6) & (x2 | ~x3 | x5 | x6));
  assign n7403 = x6 & n841 & n691 & (n828 | n3090);
  assign z441 = n7405 | n7408 | ~n7412 | (~n835 & ~n7411);
  assign n7405 = ~x5 & (n7406 | (n1392 & n1769 & n560));
  assign n7406 = ~x7 & ((n1331 & n746) | (x3 & ~n7407));
  assign n7407 = (x0 | x1 | ~x2 | x4 | ~x6) & (~x0 | x2 | (x1 ? (x4 | x6) : (~x4 | ~x6)));
  assign n7408 = ~x0 & (x4 ? ~n7409 : ~n7410);
  assign n7409 = (~x6 | ((~x2 | x3 | x7) & (x1 | ((x3 | ~x7) & (x2 | ~x3 | x7))))) & (~x1 | x6 | (x2 ? (~x3 | ~x7) : (~x3 ^ x7)));
  assign n7410 = (~x1 | x2 | ~x3 | x6) & (x1 | ~x6 | ((x3 | ~x7) & (x2 | ~x3 | x7)));
  assign n7411 = (x1 | x2 | ~x6) & (x0 | (x1 ? (x6 | (~x2 ^ x4)) : (x4 | ~x6)));
  assign n7412 = n7413 & (n640 | (~n4828 & ~n2875 & ~n3377));
  assign n7413 = (~n1586 | n5318) & (n871 | (~n746 & ~n7414));
  assign n7414 = ~x4 & ~x2 & x0 & ~x1;
  assign z442 = ~n7428 | ~n7424 | n7416 | n7420;
  assign n7416 = x7 & (n7417 | (n543 & ~n7419));
  assign n7417 = x0 & ((~x2 & ~n7418) | (~x1 & x2 & ~n1026));
  assign n7418 = (~x1 | x3 | x4 | x5 | x6) & (x1 | ~x3 | ~x4 | ~x5 | ~x6);
  assign n7419 = (x2 | x3 | x4 | ~x5 | x6) & (~x2 | ~x4 | (~x3 ^ ~x6));
  assign n7420 = n1986 & (n7421 | n7422 | ~n7423);
  assign n7421 = ~x2 & (x3 ? (x6 & (~x1 | x4)) : (x4 & ~x6));
  assign n7422 = n1145 & ((n706 & n1044) | (n1723 & n885));
  assign n7423 = (~n926 | ~n1498) & (~n570 | ~n3575);
  assign n7424 = ~n5968 & (n627 | n7425) & (~x4 | n7427);
  assign n7425 = ~n7426 & (~n543 | ~n1539) & (~n743 | n1944);
  assign n7426 = ~x1 & (x0 ? (x2 & x7) : (~x7 & (~x2 | ~x4)));
  assign n7427 = (~x0 | ~x1 | x2 | x3 | ~x7) & (x0 | x1 | ~x2 | (~x3 ^ ~x7));
  assign n7428 = ~n7429 & (~x7 | (~n7431 & (~n639 | ~n1269)));
  assign n7429 = ~x4 & ~n7430;
  assign n7430 = (x0 | ~x1 | ~x2 | (~x3 ^ ~x7)) & (x2 | ((x0 | ~x1 | ~x3 | x7) & (~x0 | x1 | (~x3 ^ x7))));
  assign n7431 = n1044 & ((n681 & n543) | (x0 & ~n1148));
  assign z443 = ~n4638 | n7433 | n7435 | (n873 & n6244);
  assign n7433 = x3 & ((n696 & n837) | (n772 & ~n7434));
  assign n7434 = (~x0 | (x2 ? (x5 | ~x6) : (~x5 | x6))) & (x0 | x2 | x5 | ~x6);
  assign n7435 = x3 & ((n1269 & n993) | (n2061 & ~n4642));
  assign z444 = ~n7441 | (x1 ? (n3926 | n7440) : ~n7437);
  assign n7437 = ~n5270 & ~n7438;
  assign n7438 = ~x6 & ((n547 & n717) | (x3 & ~n7439));
  assign n7439 = (x0 | ~x2 | x4 | ~x5 | x7) & (~x0 | x5 | (x2 ? (~x4 | x7) : (x4 | ~x7)));
  assign n7440 = ~x0 & (x2 ? ~n7278 : (n1392 & n978));
  assign n7441 = x2 ? n4647 : (n4651 & n7442);
  assign n7442 = x0 ? (x3 | (x1 ? ~x4 : (x4 | x5))) : (~x3 | (x1 ? (~x4 | ~x5) : x4));
  assign z445 = n7452 | ~n7454 | (x0 ? ~n7449 : ~n7444);
  assign n7444 = x1 ? n7445 : (~n7448 & (x4 | n7447));
  assign n7445 = (x5 | n2803 | ~x2 | x3) & (~x5 | n7446);
  assign n7446 = (~x2 | ~x3 | x4 | ~x6 | x7) & (x2 | ((x3 | ~x4 | ~x6 | x7) & (~x3 | x4 | x6 | ~x7)));
  assign n7447 = (x2 | ~x3 | x5 | ~x6 | ~x7) & (~x2 | x6 | (x3 ? (~x5 | x7) : (x5 | ~x7)));
  assign n7448 = n658 & n2385;
  assign n7449 = x1 ? (x2 | n985) : (x2 ? n7451 : n7450);
  assign n7450 = (x3 | ~x4 | x5 | ~x6 | ~x7) & (~x3 | x4 | (x5 ? (~x6 | ~x7) : (x6 | x7)));
  assign n7451 = (x3 | x4 | ~x5 | x6 | ~x7) & (~x4 | ((~x3 | (x5 ? (~x6 | ~x7) : (x6 | x7))) & (x3 | x5 | ~x6 | x7)));
  assign n7452 = ~x2 & (n5958 | (~x6 & ~n7453));
  assign n7453 = (x0 | ~x1 | x3 | ~x4) & (~x3 | ((x0 | x1 | ~x4 | x5) & (~x0 | (x1 ? (x4 | x5) : (~x4 | ~x5)))));
  assign n7454 = ~n7456 & ~n7457 & n7458 & (n1353 | n7455);
  assign n7455 = (~x0 | ~x1 | x2 | x3 | ~x5) & (x0 | ((x1 | ~x2 | x3 | ~x5) & (~x1 | (x2 ? (~x3 | ~x5) : (x3 | x5)))));
  assign n7456 = ~n1566 & ~n2276;
  assign n7457 = n2343 & (x0 ? (~x4 & x5) : (x4 ^ ~x5));
  assign n7458 = (x2 | n7459) & (x1 | ~x2 | n7460);
  assign n7459 = (x4 | x5 | ~x0 | x3) & (x0 | ((~x1 | ~x3 | ~x4 | x5) & (x1 | (x3 ? (x4 | ~x5) : (~x4 | x5)))));
  assign n7460 = (x3 | x4 | ~x6 | (x0 & ~x5)) & (~x0 | x5 | (x3 ? (x4 | ~x6) : (~x4 | x6)));
  assign z446 = ~n7475 | ~n7472 | ~n7468 | n7462 | n7466;
  assign n7462 = ~x0 & (x1 ? (n7463 | n7464) : ~n7465);
  assign n7463 = ~x7 & (x2 ? (~x3 & n2826) : (x3 & n728));
  assign n7464 = n4972 & (x2 ? (~x3 & n706) : (x3 & ~n1097));
  assign n7465 = x2 ? (n877 | n3098) : (~n530 | ~n774);
  assign n7466 = n841 & ((n1392 & ~n737) | (x3 & ~n7467));
  assign n7467 = x2 ? (x6 | (x4 ? (x5 | x7) : (~x5 | ~x7))) : (~x6 | (x4 ? (x5 | ~x7) : (~x5 | x7)));
  assign n7468 = ~n7469 & ~n7471 & (n1100 | (~n880 & ~n2535));
  assign n7469 = ~n1408 & ~n7470;
  assign n7470 = (x0 | ~x1 | x2 | x3 | ~x5) & (x1 | (x0 ? (x2 ? (~x3 | ~x5) : (x3 | x5)) : (~x2 | (~x3 ^ x5))));
  assign n7471 = ~n627 & (x0 ? (~x1 & ~n1122) : (x1 & n5525));
  assign n7472 = (~n1686 | n7473) & (n1205 | n7474);
  assign n7473 = x1 ? ((~x2 | x3 | x4 | ~x5) & (x2 | ~x3 | x5)) : (~x3 | ~x4 | (x2 ^ ~x5));
  assign n7474 = (x0 | x1 | x2 | ~n704) & (~x0 | (x1 ? (x2 | ~n704) : n7135));
  assign n7475 = ~n7476 & ~n7478;
  assign n7476 = ~x6 & (x5 ? (n1145 & ~n3486) : ~n7477);
  assign n7477 = x0 ? ((~x1 | x2 | ~x3 | x4) & (x1 | ~x2 | x3 | ~x4)) : (x1 ? (x3 | x4) : (x2 | ~x3));
  assign n7478 = ~n1008 & ((n1141 & n746) | (~x3 & ~n7479));
  assign n7479 = (x0 | ~x1 | x2 | ~x4 | ~x6) & (x6 | ((~x0 | (x1 ? (x2 | ~x4) : (~x2 | x4))) & (x0 | x1 | x2 | ~x4)));
  assign z447 = ~n7485 | ~n7490 | (x7 ? ~n7483 : ~n7481);
  assign n7481 = (~n597 | n1036) & (~x3 | (n7482 & (~n1835 | n1036)));
  assign n7482 = (x4 | ~x6 | x1 | x2) & (x0 | ((x1 | ~x4 | (~x2 ^ ~x6)) & (x4 | ~x6 | ~x1 | ~x2)));
  assign n7483 = ~n7484 & (~x5 | (~n2502 & (x0 | n5809)));
  assign n7484 = ~n615 & (x0 ? (~x1 & ~n605) : (x1 & n691));
  assign n7485 = (x6 | x7 | n7486) & (~x7 | (n7487 & (~x6 | n7486)));
  assign n7486 = (x0 | x1 | ~x2 | ~x3 | x4) & (x3 | (x0 ? (x1 ? (x2 | ~x4) : (~x2 | x4)) : (~x4 | (~x1 ^ ~x2))));
  assign n7487 = (x3 | n7489) & (x6 | n7488 | ~x3 | ~x4);
  assign n7488 = (x1 | x2) & (x0 | ~x1 | ~x2);
  assign n7489 = (x0 | x1 | ~x2 | ~x4 | x6) & (x4 | ((x6 | ((~x1 | x2) & (x0 | (~x1 & x2)))) & (x1 | ~x6 | (x0 ^ ~x2))));
  assign n7490 = ~n7491 & (x7 | (x0 & n7494) | (~x0 & n7496));
  assign n7491 = ~n1353 & (x1 ? ~n7493 : ~n7492);
  assign n7492 = (x0 | x2 | ~x5 | (~x3 ^ ~x7)) & (x5 | ((~x0 | x2 | x7) & (~x2 | ((~x3 | ~x7) & (x0 | x3 | x7)))));
  assign n7493 = (~x0 | x2 | x3 | ~x5 | x7) & (x0 | ((x2 | ~x3 | x5 | ~x7) & (~x2 | ~x5 | (~x3 ^ ~x7))));
  assign n7494 = (x2 | n7495) & (x1 | ~x2 | n4302);
  assign n7495 = (x5 | ~x6 | ~x1 | x4) & (x1 | ~x5 | (x3 ? (~x4 | x6) : (x4 | ~x6)));
  assign n7496 = (n605 | n4687) & (x4 | ~n1317 | n2291);
  assign z448 = n7512 | n7510 | n7506 | n7498 | n7503;
  assign n7498 = x5 & (n7501 | (x3 & (n7499 | ~n7500)));
  assign n7499 = n570 & (x0 ? ~n1850 : n569);
  assign n7500 = (~n548 | ~n733) & (n643 | (~n7414 & ~n5895));
  assign n7501 = ~x3 & ((n733 & n1585) | (n570 & ~n7502));
  assign n7502 = (x0 | ~x4 | x6 | ~x7) & (~x0 | (x4 ? (~x6 | x7) : (x6 | ~x7)));
  assign n7503 = ~n640 & (x4 ? ~n7504 : ~n7505);
  assign n7504 = (x0 | ((x3 | ~x5) & (~x1 | ~x3 | x5))) & (~x1 | x2 | x3 | ~x5) & (x1 | ((~x2 | x3 | ~x5) & (~x0 | ~x3 | x5)));
  assign n7505 = (x0 | ~x1 | x2 | x3 | x5) & (x1 | (x0 ? (x2 ? (x3 | ~x5) : x5) : (~x2 | (~x3 ^ ~x5))));
  assign n7506 = ~x1 & (~n7508 | (~x2 & ~n7507));
  assign n7507 = (x0 | ~x3 | (x4 ? (x5 | ~x7) : (~x5 | x7))) & (x3 | ((x4 | ~x5 | ~x7) & (x5 | x7 | ~x0 | ~x4)));
  assign n7508 = (~n867 | ~n1783) & (n835 | n7509);
  assign n7509 = (x0 | ~x2 | ~x4 | x5) & (~x0 | (x2 ? (x4 | x5) : (~x4 | ~x5)));
  assign n7510 = n1445 & ~n7511;
  assign n7511 = (x0 | (x3 ? ((~x5 | x7) & (x2 | x5 | ~x7)) : ((~x5 | ~x7) & (~x2 | x5 | x7)))) & (x2 | x3 | ((~x5 | ~x7) & (~x0 | x5 | x7)));
  assign n7512 = ~x5 & (n7515 | n7516 | n7513 | n7514);
  assign n7513 = n895 & (n3684 | (x3 & ~n3319));
  assign n7514 = ~n643 & (n2030 | (~x0 & ~n1062));
  assign n7515 = ~n3762 & ((n774 & n1769) | (n1392 & n569));
  assign n7516 = ~x0 & ((n550 & n689) | (n548 & n2135));
  assign z449 = n7527 | ~n7531 | (x0 ? ~n7518 : ~n7521);
  assign n7518 = ~n4428 & (x1 | (~x6 & n7519) | (x6 & n7520));
  assign n7519 = x2 ? (x4 ? (x5 | ~x7) : (~x5 | x7)) : (x3 ? (x4 ? (x5 | x7) : (~x5 | ~x7)) : (x7 | (~x4 ^ ~x5)));
  assign n7520 = (~x2 | x3 | x4 | x5 | ~x7) & (x2 | ((x3 | ~x4 | ~x5 | x7) & (~x7 | (x3 ? (~x4 ^ ~x5) : (x4 | ~x5)))));
  assign n7521 = x5 ? (~n7526 & (~x3 | n7525)) : n7522;
  assign n7522 = x4 ? n7523 : (x6 | n7524);
  assign n7523 = (~x7 | ((x1 | x2 | ~x3 | ~x6) & (~x1 | (x2 ? (~x3 | ~x6) : x6)))) & (x1 | ~x2 | ~x6 | (x3 & x7));
  assign n7524 = (x3 | ~x7 | ~x1 | x2) & (x1 | ~x2 | (~x3 & x7));
  assign n7525 = x1 ? (~x2 | (x4 ? (x6 | ~x7) : (~x6 | x7))) : ((~x4 | x6 | x7) & (x2 | (x4 ? x6 : (~x6 | x7))));
  assign n7526 = n689 & ((n569 & n1084) | (x2 & ~n2803));
  assign n7527 = ~n643 & (n7529 | n7530 | n3694 | n7528);
  assign n7528 = x0 & ((~x1 & x2 & x4 & x5) | (x1 & ~x2 & ~x4 & ~x5));
  assign n7529 = n828 & (x0 ? (~x1 & ~x2) : (x1 ? (~x2 & x5) : (x2 & ~x5)));
  assign n7530 = ~x0 & (x1 ? (x2 ? (~x4 & ~x5) : (x4 & x5)) : (~x4 & (x2 ^ ~x5)));
  assign n7531 = ~n7533 & ~n7534 & ~n7536 & (n615 | n7532);
  assign n7532 = (~x2 | x5 | x7 | ~x0 | x1) & (x0 | ((~x5 | ~x7 | x1 | x2) & (~x1 | (x2 ? (~x5 | ~x7) : (x5 | x7)))));
  assign n7533 = ~n2803 & (x0 ? (x1 ? (~x2 & ~x3) : (x2 & x3)) : (x1 ? (x2 ^ x3) : (~x2 & ~x3)));
  assign n7534 = ~x1 & ((n2435 & n1668) | (n743 & ~n7535));
  assign n7535 = (x6 | x7 | ~x3 | x4) & (~x6 | ~x7 | x3 | ~x4);
  assign n7536 = ~n2075 & n543 & n1857;
  assign z450 = ~n7548 | (~x1 & ~n7538) | (~x0 & ~n7545);
  assign n7538 = x6 ? n7542 : (n7540 & (x3 | n7539));
  assign n7539 = x0 ? ((~x4 | x5 | ~x7) & (x2 | x4 | ~x5 | x7)) : (x4 | ~x5 | (x2 ^ ~x7));
  assign n7540 = n7541 & (n1794 | n5108) & (~n549 | ~n670);
  assign n7541 = (x0 | ~x2 | x3 | x5 | ~x7) & (~x0 | x2 | ~x3 | ~x5 | x7);
  assign n7542 = n7544 & (n697 | n732) & (x3 | n7543);
  assign n7543 = (~x0 | x5 | x7 | (x2 & x4)) & (~x7 | ((x4 | ~x5 | ~x0 | x2) & (x0 | ~x4 | (~x2 ^ ~x5))));
  assign n7544 = (x2 | ~x3 | ~x4 | x5 | x7) & (~x2 | x3 | x4 | ~x5 | ~x7);
  assign n7545 = (~x1 | n7546) & (x1 | ~x3 | ~x4 | n7547);
  assign n7546 = (x2 | x3 | (x4 ? (~x5 | x7) : (x5 | ~x7))) & (~x3 | ((x5 | ~x7 | x2 | ~x4) & (~x2 | ((~x5 | ~x7) & (~x4 | x5 | x7)))));
  assign n7547 = x2 ? (x5 ^ ~x7) : (~x5 | ~x7);
  assign n7548 = n7553 & (~x1 | (~n7549 & ~n7551 & n7552));
  assign n7549 = ~x7 & ((~n5570 & n7550) | (n2446 & n3895));
  assign n7550 = ~x3 & ~x4 & (x5 ^ ~x6);
  assign n7551 = ~n1998 & n1465 & ~n1198;
  assign n7552 = (~n547 | ~n601) & (~n1693 | ~n978);
  assign n7553 = (n1548 | n7554) & (~n841 | n7555);
  assign n7554 = (((x1 | ~x5) & (x0 | ~x1 | x5)) | (~x2 ^ x7)) & (x2 | x5 | x7 | (~x0 ^ ~x1));
  assign n7555 = (x2 | ~x3 | x4 | x5 | x7) & (~x2 | ((x3 | x4 | ~x5 | x7) & (~x3 | x5 | ~x7)));
  assign z451 = n7562 | ~n7564 | ~n7568 | (~x1 & ~n7557);
  assign n7557 = x0 ? (~n7561 & (x4 | n7560)) : n7558;
  assign n7558 = x2 ? (~n2836 & (~x3 | ~n728)) : n7559;
  assign n7559 = (~x5 | x6 | x7 | ~x3 | x4) & (x3 | x5 | (x4 ? (~x6 ^ ~x7) : (~x6 | x7)));
  assign n7560 = (x2 | x3 | x5 | x6 | ~x7) & (x7 | ((x5 | x6 | x2 | ~x3) & (~x2 | (x3 ? (~x5 | x6) : (x5 | ~x6)))));
  assign n7561 = ~n3309 & n1392 & ~x5 & x6;
  assign n7562 = n543 & (n7563 | (x5 & n902 & ~n4773));
  assign n7563 = ~x3 & ((n813 & n859) | (~x2 & ~n1282));
  assign n7564 = ~n7566 & (~n5479 | n7565);
  assign n7565 = (x4 | x7 | x2 | x3) & (x1 | ((x2 | ~x3 | ~x4 | ~x7) & (~x2 | (x3 ? (~x4 | x7) : (x4 | ~x7)))));
  assign n7566 = ~n714 & ((n560 & n1403) | (~x6 & ~n7567));
  assign n7567 = (x0 | ~x1 | ~x2 | ~x3 | x7) & (~x0 | x1 | (x2 ? (x3 | x7) : (~x3 | ~x7)));
  assign n7568 = ~n7569 & n7573 & (n647 | n7572);
  assign n7569 = ~x0 & (x1 ? (~n1744 & ~n7570) : ~n7571);
  assign n7570 = (~x6 | x7) & (x2 | x6 | ~x7);
  assign n7571 = (~x2 | (x3 ? (~x4 | x6) : (x4 | ~x6))) & (~x6 | ((x2 | ~x3 | ~x4 | x7) & (x3 | x4 | ~x7)));
  assign n7572 = (x0 | x1 | ~x2 | ~x6 | ~x7) & (x6 | ((x0 | (x7 & (~x1 | x2))) & (~x1 | x2 | x7) & (x1 | ((~x2 | x7) & (~x0 | x2 | ~x7)))));
  assign n7573 = (~n560 | ~n3057) & (~x7 | n7574);
  assign n7574 = x0 ? ((x1 | ~x2 | ~x3 | x6) & (~x1 | x2 | x3 | ~x6)) : ((x1 | x2 | ~x3 | x6) & (~x1 | ~x2 | (~x3 ^ x6)));
  assign z452 = ~n7583 | (x4 ? ~n7580 : ~n7576);
  assign n7576 = x0 ? (~n7579 & (~n530 | ~n1439)) : n7577;
  assign n7577 = (~n558 | ~n658) & (~x6 | n7578);
  assign n7578 = (x5 | x7 | x1 | x3) & (~x1 | ~x2 | (x3 ? (x5 | x7) : (~x5 | ~x7)));
  assign n7579 = n934 & ((n1857 & n1188) | (x1 & ~n3315));
  assign n7580 = x5 ? n7582 : n7581;
  assign n7581 = x6 ? (~x7 | n4075) : ((x7 | n4075) & (x2 | ~x7 | n1682));
  assign n7582 = (~n1269 | ~n3352) & (n643 | n4066);
  assign n7583 = ~n7584 & n7587 & (n671 | n7586);
  assign n7584 = ~x2 & ((n4569 & ~n6098) | (~x4 & ~n7585));
  assign n7585 = (x0 | ~x1 | ~x7 | (~x3 ^ ~x5)) & (x1 | ((~x5 | ~x7 | x0 | x3) & (~x0 | (x3 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n7586 = (x0 | ~x1 | x2 | x3 | ~x5) & (x1 | ((~x3 | x5 | x0 | ~x2) & (~x0 | x2 | (~x3 ^ ~x5))));
  assign n7587 = (n1218 | n7588) & (~n526 | ~n828 | ~n1209);
  assign n7588 = (~x0 | ((~x1 | x2 | x3 | ~x5) & (x1 | ~x2 | x5))) & (~x3 | ((x1 | ~x2 | ~x5) & (x0 | (x5 ? x1 : x2)))) & (x0 | ~x2 | (~x5 & (~x1 | x3)));
  assign z453 = n7598 | ~n7600 | (x1 ? ~n7590 : ~n7593);
  assign n7590 = ~n7591 & (~n742 | (~x3 & ~n4900) | (x3 & n3409));
  assign n7591 = ~x2 & (x5 ? (n622 & n6470) : ~n7592);
  assign n7592 = (x0 | ~x3 | ~x4 | x6 | ~x7) & (x7 | ((x0 | x3 | ~x4 | ~x6) & (~x0 | x4 | (~x3 ^ ~x6))));
  assign n7593 = x2 ? (x0 ? n7594 : n7595) : n7596;
  assign n7594 = (x3 | ~x4 | x5 | x6 | ~x7) & (~x3 | x4 | ~x5 | ~x6 | x7);
  assign n7595 = (x3 | x4 | x5 | x6 | x7) & (~x4 | ((~x6 | ~x7 | x3 | ~x5) & (~x3 | x6 | (~x5 ^ x7))));
  assign n7596 = x5 ? (~n1857 | ~n5168) : n7597;
  assign n7597 = (x0 | x3 | x6 | ~x7) & (~x3 | ((~x6 | ~x7 | x0 | x4) & (~x0 | x7 | (~x4 ^ ~x6))));
  assign n7598 = ~n1198 & ~n7599;
  assign n7599 = (x0 | ~x1 | x2 | (~x3 ^ ~x4)) & (x1 | ((x3 | ~x4 | x0 | x2) & (~x0 | ~x2 | (~x3 ^ x4))));
  assign n7600 = n7601 & ~n7603 & ~n7605 & (n2259 | n4099);
  assign n7601 = x0 | (n7602 & (~n561 | ~n570));
  assign n7602 = x1 ? ((~x2 | x3 | ~x4 | ~x5) & (x2 | ~x3 | x4 | x5)) : (~x3 | (x2 ? (x4 | x5) : ~x5));
  assign n7603 = n841 & ((x2 & ~n1920) | (n1044 & ~n7604));
  assign n7604 = ~x4 & x5;
  assign n7605 = ~x4 & ((n3269 & n837) | (n653 & ~n7606));
  assign n7606 = (x1 | x2 | x5 | ~x6) & (~x1 | ~x2 | ~x5 | x6);
  assign z454 = ~n7619 | ~n7615 | ~n7613 | n7608 | n7612;
  assign n7608 = ~n643 & ((~n1480 & n1167) | n7609 | ~n7611);
  assign n7609 = n1044 & (x0 ? ~n7610 : n2074);
  assign n7610 = x1 ? (~x4 | ~x5) : (x4 | x5);
  assign n7611 = ~n3694 & (n753 | n1433) & (~n731 | ~n746);
  assign n7612 = n1365 & ((~x2 & ~x4 & x5 & ~x6) | (x2 & (x4 ? x6 : (~x5 & ~x6))));
  assign n7613 = (n5411 | n1939) & (n2022 | n7614);
  assign n7614 = (~x0 | x2 | x3) & (x0 | ~x2 | ~x3 | x5);
  assign n7615 = ~n7616 & (n1408 | (n7618 & (~n626 | ~n6084)));
  assign n7616 = ~x1 & (x5 ? (n1181 & ~n3427) : ~n7617);
  assign n7617 = (x0 | ~x2 | x3 | x6 | x7) & (~x0 | ((~x2 | x3 | ~x6 | ~x7) & (x2 | ~x3 | x6 | x7)));
  assign n7618 = (n2373 | n2864) & (n765 | n4066);
  assign n7619 = x0 | (n7620 & ~n7621 & (~n601 | ~n1439));
  assign n7620 = x1 ? (~n3425 & (~n1044 | ~n696)) : n3424;
  assign n7621 = ~x2 & ((~n7610 & ~n5269) | (n658 & n2871));
  assign z455 = ~n7631 | (x0 ? ~n7628 : ~n7623);
  assign n7623 = x6 ? n7624 : (~n7627 & (~x4 | n7626));
  assign n7624 = x2 ? (~n1821 & (~n1317 | ~n2209)) : n7625;
  assign n7625 = x7 ? (x1 ? (x3 ? (~x4 | x5) : ~x5) : (x3 ? (x4 | ~x5) : (~x4 | x5))) : (x1 ? (x4 | ~x5) : (~x3 | (~x4 ^ ~x5)));
  assign n7626 = (x1 | ~x3 | ~x5 | (x2 ^ ~x7)) & (x3 | (~x2 ^ ~x7) | (x1 ^ x5));
  assign n7627 = n1156 & ((n1429 & n1188) | (x1 & ~n2830));
  assign n7628 = (x2 | n7629) & (x1 | ~x2 | n7630);
  assign n7629 = (n1042 | (~n2723 & ~n1585)) & (~n530 | ~n3194);
  assign n7630 = (x3 | x4 | ~x5 | ~x6 | x7) & (x6 | ((x3 | x4 | ~x5 | ~x7) & (~x3 | x5 | (x4 ^ ~x7))));
  assign n7631 = n7632 & n7634 & ~n7637 & (n671 | n7636);
  assign n7632 = (~n4413 | ~n837) & (n1218 | n7633);
  assign n7633 = x0 ? ((x1 | ~x2 | ~x3 | ~x5) & (~x1 | x2 | x3 | x5)) : ((~x1 | ~x2 | ~x3 | x5) & (x3 | ~x5 | x1 | x2));
  assign n7634 = (n765 | (~n1265 & ~n2030)) & (n1744 | n7635);
  assign n7635 = (~x0 | x1 | ~x2 | x5 | ~x7) & (x0 | ((~x1 | ~x2 | ~x5 | x7) & (x5 | ~x7 | x1 | x2)));
  assign n7636 = (~x0 | x1 | x2 | ~x5) & (x0 | x5 | (x1 ? (x2 | x3) : (~x2 | ~x3)));
  assign n7637 = ~x0 & ((~n2099 & ~n2864) | (n885 & n867));
  assign z456 = n7648 | ~n7651 | (x2 ? ~n7644 : ~n7639);
  assign n7639 = x3 ? n7642 : (x0 ? n7640 : n7641);
  assign n7640 = (~x1 | x4 | x5 | ~x6 | x7) & (~x4 | ((~x5 | x6 | ~x7) & (x1 | ((x6 | ~x7) & (~x5 | ~x6 | x7)))));
  assign n7641 = (~x1 | x4 | ~x5 | x6 | ~x7) & (x7 | ((~x1 | x5 | (~x4 ^ ~x6)) & (~x5 | ((x4 | ~x6) & (x1 | ~x4 | x6)))));
  assign n7642 = (~n657 | ~n978) & (~x7 | n7643);
  assign n7643 = (x0 | ~x1 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (x1 | (~x5 ^ ~x6) | (x0 ^ x4));
  assign n7644 = ~n7645 & (~n2758 | ~n1244) & (n835 | n7647);
  assign n7645 = x4 & (x0 ? (n658 & n1188) : ~n7646);
  assign n7646 = (~x1 | ~x3 | x5 | x6 | x7) & (~x6 | (x3 ^ ~x7) | (x1 ^ x5));
  assign n7647 = (x0 | ~x1 | x4 | ~x5 | x6) & (x1 | x5 | (x0 ? (~x4 ^ x6) : (x4 | x6)));
  assign n7648 = ~x3 & (x4 ? ~n7649 : ~n7650);
  assign n7649 = (x0 | ~x1 | ~x2 | x5) & (x1 | (x2 ? (~x5 | (~x0 & x6)) : (x5 | ~x6)));
  assign n7650 = (x0 | ~x1 | ~x2 | x5 | ~x6) & (~x0 | x1 | x2 | (~x5 ^ x6));
  assign n7651 = n7654 & (n1097 | n7652) & (x1 | n7653);
  assign n7652 = (x0 | ~x3 | (x1 ^ ~x4)) & (x3 | ((~x1 | x2 | ~x4) & (~x0 | (x1 ? x2 : (~x2 | x4)))));
  assign n7653 = (x0 | x3 | x4 | ~x5 | x6) & (~x3 | ((x5 | ~x6 | x0 | x4) & (~x0 | (x4 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n7654 = (~n1358 | ~n866) & (~n774 | ~n1723 | ~n560);
  assign z457 = ~n7667 | n7665 | n7663 | n7656 | n7660;
  assign n7656 = ~x1 & (n7657 | (~x5 & n622 & ~n7659));
  assign n7657 = ~x0 & ((n902 & n3476) | (~x3 & ~n7658));
  assign n7658 = (~x2 | ~x6 | ~x7 | (x4 ^ ~x5)) & (x2 | x4 | ~x5 | x6 | x7);
  assign n7659 = (x2 | ~x4 | x6 | ~x7) & (~x2 | x4 | (~x6 ^ ~x7));
  assign n7660 = ~n643 & (n7661 | (~x2 & ~n7662));
  assign n7661 = x2 & ((~x0 & ~x4 & (x1 ^ ~x5)) | (x0 & ~x1 & x4 & ~x5));
  assign n7662 = (x0 | ~x1 | x3 | x4 | x5) & (~x4 | ((x0 | x1 | x3 | ~x5) & (~x0 | (x1 ? (x3 | ~x5) : (~x3 | x5)))));
  assign n7663 = n4894 & (x0 ? (n1044 & n942) : ~n7664);
  assign n7664 = (x2 | x3 | x5 | x6 | x7) & (~x2 | ~x3 | ~x7 | (~x5 ^ ~x6));
  assign n7665 = x6 & ((~n807 & ~n7666) | (n731 & n1269));
  assign n7666 = (x3 | ~x5 | ~x1 | x2) & (x1 | (x2 ? (x3 | ~x5) : x5));
  assign n7667 = n7675 & ~n7673 & ~n7671 & ~n7668 & ~n7669;
  assign n7668 = n895 & (n662 | (~x4 & n2862));
  assign n7669 = ~n3266 & ~n7670;
  assign n7670 = (~x0 | x1 | ~x2 | ~x3 | x6) & (x0 | ~x1 | ~x6 | (~x2 ^ x3));
  assign n7671 = ~x0 & ((~n1538 & n7672) | (n530 & n3084));
  assign n7672 = ~x6 & (x1 ^ ~x5);
  assign n7673 = ~x6 & ((n560 & n959) | (~x4 & ~n7674));
  assign n7674 = (~x0 | ~x1 | x2 | x5) & (x0 | x1 | ~x5 | (~x2 & ~x3));
  assign n7675 = (n3394 | n7676) & (n1701 | n7677);
  assign n7676 = (~x2 | (x3 ? (x4 | ~x6) : (~x4 | x6))) & (x2 | ~x3 | ~x4 | x6);
  assign n7677 = x0 ? (x4 | (x1 ? (x2 | x3) : (~x2 | ~x3))) : (~x4 | (x1 ? x2 : (~x2 | ~x3)));
  assign z458 = n7690 | n7688 | ~n7685 | n7679 | n7681;
  assign n7679 = x0 & (x1 ? n6321 : ~n7680);
  assign n7680 = (~x3 | n3656) & (x7 | n1198 | x2 | x3);
  assign n7681 = ~n1097 & (n7683 | ~n7684 | (~x2 & ~n7682));
  assign n7682 = (~x0 | ~x1 | x3 | x4 | x7) & (x0 | ~x3 | (x1 ? (x4 | x7) : (~x4 | ~x7)));
  assign n7683 = x0 & ~x1 & (x2 ? (x3 & ~x7) : x7);
  assign n7684 = x0 | (x1 ? (x2 | ~n683) : (~x2 | ~n2647));
  assign n7685 = (x2 | n7687) & (~n5802 | ~n746) & (~x2 | n7686);
  assign n7686 = (x0 | ~x1 | (x3 ? (~x5 | ~x7) : (x5 | x7))) & (x1 | ((x3 | ~x5 | x7) & (x5 | ~x7 | (~x0 & ~x3))));
  assign n7687 = (~x0 | x1 | ~x3 | ~x5 | x7) & (x0 | x3 | ~x7 | (~x1 ^ x5));
  assign n7688 = ~x7 & ((n639 & n1269) | (~x5 & ~n7689));
  assign n7689 = (x0 | x1 | x2 | x3 | ~x4) & (~x1 | ((~x3 | x4 | x0 | ~x2) & (~x0 | x2 | (~x3 ^ x4))));
  assign n7690 = ~x0 & (n7691 | n7694 | (~n1198 & ~n7693));
  assign n7691 = ~x7 & (x3 ? ~n7692 : (n804 & ~n1040));
  assign n7692 = (x1 | ~x2 | ~x4 | ~x5 | ~x6) & (~x1 | x6 | (x2 ? (x4 | ~x5) : (~x4 | x5)));
  assign n7693 = (x1 | x2 | ~x3 | x7) & (~x1 | (x2 ? (x3 ? (~x4 | x7) : (x4 | ~x7)) : (~x3 | ~x7)));
  assign n7694 = n619 & (n7695 | (n596 & n926));
  assign n7695 = x6 & x5 & ~x4 & ~x2 & x3;
  assign z459 = ~n7707 | n7704 | n7697 | n7700;
  assign n7697 = x7 & ((n733 & n1202) | (~x1 & ~n7698));
  assign n7698 = (~x2 | n7699) & (x0 | x2 | ~x3 | ~n5163);
  assign n7699 = (x0 | x3 | ~x4 | x5 | ~x6) & (~x0 | x6 | (x3 ? (~x4 | x5) : (x4 | ~x5)));
  assign n7700 = ~x7 & (n7701 | (n927 & ~n7703));
  assign n7701 = ~x1 & ((n5479 & ~n3538) | (n3074 & ~n7702));
  assign n7702 = (~x2 | ~x3 | ~x4 | x5) & (x3 | ((x4 | ~x5) & (x2 | ~x4 | x5)));
  assign n7703 = (~x0 | x2 | x4 | x5 | x6) & (x0 | (x2 ? (x4 | (~x5 ^ ~x6)) : (~x4 | (~x5 ^ x6))));
  assign n7704 = ~x1 & ((x2 & ~n7705) | (n1181 & ~n7706));
  assign n7705 = (x0 | ~x3 | ~x4 | (~x6 ^ x7)) & (x4 | ((x0 | x3 | ~x6 | ~x7) & (~x0 | x6 | (~x3 ^ ~x7))));
  assign n7706 = (~x3 | x4 | ~x6 | x7) & (x3 | (x4 ? (~x6 | x7) : (x6 | ~x7)));
  assign n7707 = ~n7709 & n7711 & (x0 ? n7708 : n7710);
  assign n7708 = (x4 | ~x6 | x2 | x3) & (x1 | (x2 ? (~x4 | (~x3 ^ ~x6)) : (x3 | ~x6)));
  assign n7709 = ~n640 & (n4058 | (n743 & n4416));
  assign n7710 = x1 ? ((~x2 | x3 | ~x4 | x6) & (x2 | ~x3 | x4 | ~x6)) : (~x3 | (x2 ? (x4 | x6) : (~x4 | ~x6)));
  assign n7711 = (n697 | n7712) & (~n543 | n7713);
  assign n7712 = (x0 | ~x4 | (x1 ? (~x3 | ~x6) : (x3 | x6))) & (~x0 | x1 | ~x3 | x4 | ~x6);
  assign n7713 = (x2 | x3 | (~x6 ^ x7)) & (~x2 | ~x3 | x6 | ~x7);
  assign z460 = n7715 | ~n7722 | ~n7725 | (~x2 & ~n7721);
  assign n7715 = ~x1 & (n7719 | (~x4 & (n7716 | ~n7717)));
  assign n7716 = n569 & (n2177 | (~x3 & ~x5 & ~n6891));
  assign n7717 = (~n3434 | ~n951) & (n640 | n7718);
  assign n7718 = (~x3 | ~x5 | ~x0 | x2) & (x3 | x5 | x0 | ~x2);
  assign n7719 = x4 & ((n547 & n813) | (x2 & ~n7720));
  assign n7720 = (~x5 | x6 | x7 | ~x0 | x3) & (x0 | ~x7 | (x3 ? (x5 | ~x6) : (~x5 | x6)));
  assign n7721 = (~x0 | ~x4 | ~x7 | (x1 ^ ~x3)) & ((~x1 ^ x4) | (x0 ? (x3 | x7) : (~x3 ^ x7)));
  assign n7722 = ~n7724 & (~n1621 | ~n3791) & (n981 | n7723);
  assign n7723 = (x0 | x1 | ~x2 | ~x4 | x7) & (~x0 | ~x7 | (x1 ? (x2 | x4) : (~x2 | ~x4)));
  assign n7724 = n543 & ((n1044 & n635) | (~n765 & n1619));
  assign n7725 = (~x2 | n7726) & (x1 | n7727);
  assign n7726 = (x0 | ~x1 | x3 | (~x4 ^ x7)) & (~x3 | ((x0 | (x1 ? (~x4 | ~x7) : (x4 | x7))) & (x4 | ~x7 | ~x0 | x1)));
  assign n7727 = (x4 | n7729) & (n877 | n7728 | ~x2 | ~x4);
  assign n7728 = x0 ^ ~x7;
  assign n7729 = (x0 | ~x7 | (x2 ? (x3 | ~x5) : (~x3 | x5))) & (x7 | ((x2 | x3 | ~x5) & (~x0 | ((x3 | ~x5) & (x2 | ~x3 | x5)))));
  assign z461 = n7735 | ~n7743 | (x0 ? ~n7731 : ~n7739);
  assign n7731 = ~n7733 & (x1 | (~n7732 & (~n885 | n5658)));
  assign n7732 = n1044 & (n588 | (x5 & ~n6633));
  assign n7733 = n632 & ~n7734;
  assign n7734 = (~x3 | x4 | x5 | ~x6 | x7) & (x3 | ((x6 | ~x7 | ~x4 | ~x5) & (x4 | (x5 ? (~x6 | x7) : (x6 | ~x7)))));
  assign n7735 = ~x5 & (n7737 | ~n7738 | (~x2 & ~n7736));
  assign n7736 = (~x0 | ((~x3 | x4 | x6) & (x1 | x3 | ~x4))) & (x1 | ~x3 | x4) & (~x1 | ((x3 | x4 | ~x6) & (~x4 | x6 | x0 | ~x3)));
  assign n7737 = ~x0 & ((~x1 & x2 & x4 & ~x6) | (x1 & x6 & (x2 ^ x4)));
  assign n7738 = ~x2 | (x0 ? (x1 | ~n1479) : (~x1 | ~n761));
  assign n7739 = ~n7740 & (~n804 | n7742);
  assign n7740 = x1 & ((n1044 & n978) | (x7 & ~n7741));
  assign n7741 = (~x2 | ~x3 | ~x4 | x5 | ~x6) & (x2 | x6 | (x3 ? (x4 | ~x5) : x5));
  assign n7742 = (~x5 | x6 | x7 | ~x3 | x4) & (x3 | ((~x6 | ~x7 | x4 | x5) & (~x4 | (x5 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n7743 = ~n7744 & (~x5 | (n7747 & (x0 | n7746)));
  assign n7744 = ~n1353 & ~n7745;
  assign n7745 = (x1 | ~x2 | x3 | x5) & (~x5 | ((x0 | ~x1 | ~x2 | x3) & (~x0 | x2 | (~x1 ^ x3))));
  assign n7746 = x2 ? ((x4 | x6 | x1 | ~x3) & (~x1 | (x3 ? ~x4 : (x4 | ~x6)))) : ((x3 | x4 | x6) & (x1 | (~x3 ^ ~x4)));
  assign n7747 = (x2 | n615 | x0 | ~x1) & (x1 | ((~x2 | n615) & (~x0 | x2 | ~n745)));
  assign z462 = ~n7757 | (x2 ? (n7749 | n7750) : ~n7752);
  assign n7749 = ~n1100 & ((~x0 & ~x3 & x7) | (~x1 & ((~x3 & x7) | (x0 & x3 & ~x7))));
  assign n7750 = x3 & (x0 ? (n1145 & n951) : ~n7751);
  assign n7751 = (~x1 | ~x4 | x5 | ~x6 | x7) & (x4 | ~x7 | ((x5 | x6) & (x1 | ~x5 | ~x6)));
  assign n7752 = ~n7756 & (n1097 | n7753) & (x7 | n7754);
  assign n7753 = x0 ? ((x1 | ~x3 | ~x4 | ~x7) & (x3 | x4 | x7)) : (~x4 | ((x3 | x7) & (~x1 | ~x3 | ~x7)));
  assign n7754 = (~n774 | n7755) & (x3 | n573 | n682);
  assign n7755 = (~x0 | ~x1 | x5 | ~x6) & (x0 | ~x5 | x6);
  assign n7756 = n619 & ((n704 & n536) | (~x0 & ~n928));
  assign n7757 = x2 ? n7760 : (x0 ? n7758 : n7759);
  assign n7758 = ((x1 & x3) | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (x6 | ((x4 | x5 | ~x1 | ~x3) & (x1 | x3 | ~x5)));
  assign n7759 = (x5 & (x3 | (x4 & x6))) | (~x1 & ~x4 & ~x6) | (~x5 & (~x3 | (x1 & ~x6)));
  assign n7760 = n710 | (n2077 & (n1744 | n1097));
  assign z463 = n7762 | n7766 | ~n7773 | (~n823 & ~n7770);
  assign n7762 = ~x1 & (n7763 | (n825 & ~n7765));
  assign n7763 = ~x3 & ((n951 & n2058) | (~x7 & ~n7764));
  assign n7764 = x0 ? (x6 | (x2 ? (x4 | x5) : (~x4 | ~x5))) : (~x6 | (x2 ? (~x4 ^ x5) : (~x4 ^ ~x5)));
  assign n7765 = (~x2 | x4 | ~x5 | ~x6 | x7) & (x2 | ~x7 | (x4 ? (~x5 ^ x6) : (x5 | x6)));
  assign n7766 = ~n640 & (n7768 | ~n7769 | (~x0 & ~n7767));
  assign n7767 = (x2 | ((~x3 | x4 | ~x5) & (x1 | x3 | ~x4 | x5))) & (x1 | ~x5 | ((x3 | x4) & (~x2 | ~x3 | ~x4))) & (~x2 | x4 | x5 | (~x1 & x3));
  assign n7768 = n564 & (n1195 | (~x1 & x3 & ~n968));
  assign n7769 = (n1062 | n2585) & (n1744 | n605 | n823);
  assign n7770 = (~x4 | n7772) & (x3 | x4 | x6 | ~n7771);
  assign n7771 = x7 & (x2 ^ x5);
  assign n7772 = (x2 | ~x5 | (x3 ? (x6 | ~x7) : (~x6 | x7))) & (~x2 | x5 | ~x6 | x7);
  assign n7773 = ~n7776 & ~n7779 & (x3 ? n7778 : n7774);
  assign n7774 = (~n548 | ~n1269) & (~n1084 | n7775);
  assign n7775 = (x0 | x1 | x6 | ~x7) & (~x6 | x7 | (~x0 & ~x1));
  assign n7776 = ~n7777 & ((x0 & ~x1 & ~n605) | (x1 & ~n2267));
  assign n7777 = (~x3 | x4 | ~x6 | x7) & (x3 | ~x4 | x6 | ~x7);
  assign n7778 = x4 ? (n710 | n785) : (~n1769 | ~n560);
  assign n7779 = n3047 & x7 & ~n1447;
  assign z464 = ~n7794 | n7792 | n7789 | n7781 | n7784;
  assign n7781 = ~x2 & ((n1511 & n7002) | (x3 & ~n7782));
  assign n7782 = x0 ? (~n3573 & (~n772 | ~n978)) : n7783;
  assign n7783 = (x1 | ~x4 | x5 | ~x6 | ~x7) & (~x1 | ~x5 | x7 | (~x4 ^ x6));
  assign n7784 = ~n640 & (~n7786 | (~x1 & ~n7785));
  assign n7785 = (x0 | x2 | x3 | ~x4 | x5) & (~x3 | ((~x2 | (x0 ? (x4 | ~x5) : (~x4 | x5))) & (x0 | x2 | (~x4 ^ ~x5))));
  assign n7786 = ~n7787 & ~n7788 & (~n746 | ~n1641);
  assign n7787 = ~x3 & ((x0 & x1 & ~x2 & ~x5) | (~x0 & ~x1 & x2 & x5));
  assign n7788 = (x0 ^ x1) & (x2 ? (~x3 & x5) : ~x5);
  assign n7789 = ~n643 & ((n742 & n7790) | (x5 & ~n7791));
  assign n7790 = ~x3 & ~x5 & (~x1 ^ x4);
  assign n7791 = (~x3 | ~x4 | x0 | ~x2) & (x2 | ((x0 | x1 | x3 | ~x4) & (~x0 | x4 | (~x1 ^ x3))));
  assign n7792 = ~n1647 & ~n7793;
  assign n7793 = (x3 | (x0 ? (x1 ? (x2 | ~x4) : (~x2 | x4)) : (~x1 | x4))) & (x0 | x2 | ~x3 | (x1 & ~x4));
  assign n7794 = n7796 & ~n7798 & ~n7799 & (n1116 | n7795);
  assign n7795 = (~x0 | x1 | ~x2 | ~x3 | ~x4) & (x0 | x4 | ((~x2 | ~x3) & (x1 | x2 | x3)));
  assign n7796 = (n1014 | n7797) & (~n699 | ~n1621);
  assign n7797 = (~x0 | x1 | ~x2 | ~x3 | x6) & (x0 | ~x1 | ~x6 | (~x2 ^ ~x3));
  assign n7798 = n1467 & ((n653 & n1585) | (x0 & ~n7777));
  assign n7799 = n570 & ((n3074 & ~n4213) | (n1070 & n1908));
  assign z465 = ~n7814 | (x2 ? ~n7801 : (n7806 | n7810));
  assign n7801 = ~n7802 & (n643 | n7804) & (n640 | n7805);
  assign n7802 = ~x0 & ((n530 & n3194) | (~x6 & ~n7803));
  assign n7803 = (x1 | x3 | (x4 ? (~x5 | x7) : (x5 | ~x7))) & (~x3 | ((~x1 | (x4 ? (~x5 | ~x7) : (x5 | x7))) & (x5 | ~x7 | x1 | ~x4)));
  assign n7804 = x0 ? (x1 | (x3 ? (~x4 | ~x5) : (~x4 ^ x5))) : ((x1 | ~x3 | x4 | ~x5) & (~x1 | (x3 ? (~x4 | x5) : x4)));
  assign n7805 = (~x0 | x1 | ~x3 | x4) & (x0 | x3 | ~x4 | (~x1 ^ ~x5));
  assign n7806 = ~x5 & (n7807 | n7808 | (x0 & ~n7809));
  assign n7807 = ~n640 & ((x0 & x1 & ~x3 & x4) | (~x0 & (x1 ? (x3 ^ ~x4) : (x3 & ~x4))));
  assign n7808 = ~n1433 & ((x6 & ~x7) | (~x1 & ~x6 & x7));
  assign n7809 = (~x1 | x3 | x4 | x6 | ~x7) & (x1 | ~x4 | (x3 ? (~x6 | ~x7) : (x6 | x7)));
  assign n7810 = x5 & (n7812 | n7813 | (~x3 & ~n7811));
  assign n7811 = (x0 | ~x1 | ~x4 | x6 | ~x7) & (x7 | ((~x4 | ~x6 | x0 | ~x1) & ((~x1 ^ x6) | (x0 ^ x4))));
  assign n7812 = ~n640 & (x0 ? (~x1 & ~n1744) : n774);
  assign n7813 = n2724 & x3 & ~x0 & ~x1;
  assign n7814 = ~n7817 & (x3 | (~n7815 & n7816));
  assign n7815 = ~n1353 & ((~x0 & ~x1 & x2 & x5) | (x0 & ~x2 & (x1 ^ ~x5)));
  assign n7816 = (~x0 | x1 | ~x2 | n1040) & (x0 | (x1 ? n2760 : (x2 | n1040)));
  assign n7817 = x3 & ((~x1 & ~n7818) | (n543 & ~n7819));
  assign n7818 = x4 ? ((x0 | ~x2 | ~x5 | x6) & (x5 | (x0 ? (~x2 ^ ~x6) : (x2 | ~x6)))) : ((~x0 | x2 | ~x5 | x6) & (x0 | ~x2 | x5 | ~x6));
  assign n7819 = x2 ? (x4 | ~x6) : (x4 ? (~x5 | ~x6) : (x5 | x6));
  assign z466 = n7836 | n7834 | ~n7827 | n7821 | n7825;
  assign n7821 = ~x2 & ((~x5 & ~n7822) | (n551 & ~n7824));
  assign n7822 = (~x1 | n7823) & (~x3 | ~n2724 | ~x0 | x1);
  assign n7823 = (x0 | x3 | ~x4 | ~x6 | x7) & (~x0 | ~x3 | x4 | x6 | ~x7);
  assign n7824 = (~x0 | x3 | ~x4 | ~x6 | x7) & (x0 | ((~x3 | ~x4 | ~x6 | x7) & (x6 | ~x7 | x3 | x4)));
  assign n7825 = ~n640 & (n4126 | n7826 | (~n1134 & ~n4075));
  assign n7826 = n543 & (n2775 | (n2332 & n596));
  assign n7827 = ~n7828 & ~n7830 & n7833 & (n1014 | n4075);
  assign n7828 = ~n1134 & ~n7829;
  assign n7829 = (x0 | ~x1 | x2 | (~x3 ^ ~x7)) & (x1 | ((x3 | ~x7 | x0 | x2) & (~x0 | (x2 ? (x3 | ~x7) : (~x3 | x7)))));
  assign n7830 = ~x1 & ((x0 & ~n7831) | (n825 & ~n7832));
  assign n7831 = (x2 | x3 | ~x4 | x6 | ~x7) & (~x2 | ~x3 | x4 | ~x6 | x7);
  assign n7832 = (x2 | x4 | ~x6 | x7) & (~x2 | ~x4 | x6 | ~x7);
  assign n7833 = (~n1241 | ~n3796) & (~n746 | (~n3684 & ~n2992));
  assign n7834 = ~x1 & (n7835 | (x7 & n902 & ~n1679));
  assign n7835 = ~n1008 & (n2329 | (x0 & ~n2075));
  assign n7836 = ~n714 & ((n1209 & n1135) | (n1181 & ~n7837));
  assign n7837 = (x1 | x3 | ~x6 | x7) & (~x1 | (x3 ? (~x6 | x7) : (x6 | ~x7)));
  assign z467 = ~n7853 | n7850 | n7846 | n7839 | n7844;
  assign n7839 = ~x0 & (n7840 | (n1300 & ~n7843));
  assign n7840 = ~x6 & ((~x2 & ~n7841) | (n3517 & ~n7842));
  assign n7841 = (~x1 | x3 | ~x4 | x5 | ~x7) & (x1 | ((~x5 | ~x7 | x3 | x4) & (~x3 | x7 | (x4 & ~x5))));
  assign n7842 = x1 ? (x3 | (x4 & ~x5)) : (~x3 | ~x4);
  assign n7843 = (~x5 | ((x1 | x2 | ~x3 | ~x4) & (~x1 | x3 | (x2 & ~x4)))) & (x4 | ((~x1 | x2 | ~x3 | x5) & (x1 | (x2 ? ~x3 : (x3 | x5)))));
  assign n7844 = ~n714 & ((~n5540 & n2797) | (~x3 & ~n7845));
  assign n7845 = x0 ? ((~x1 | x2 | ~x6 | ~x7) & (x1 | ~x2 | x6 | x7)) : ((x1 | ~x2 | ~x6 | ~x7) & (x2 | x6 | x7));
  assign n7846 = ~n643 & (n7847 | n7848 | (~x4 & ~n7849));
  assign n7847 = n772 & (x0 ? ~n1916 : ~n1515);
  assign n7848 = ~n1566 & ((~x2 & ~x4 & x0 & x1) | (~x0 & (x1 ? (~x2 & x4) : (x2 & ~x4))));
  assign n7849 = (x0 | ~x1 | ~x2 | ~x5) & (x1 | ((~x3 | ~x5 | x0 | x2) & (~x0 | (x2 ? (~x3 | ~x5) : x5))));
  assign n7850 = ~x3 & (x6 ? ~n7852 : ~n7851);
  assign n7851 = x0 ? (x2 | ((~x4 | ~x5) & (~x1 | x4 | x5))) : (x1 | ~x2 | (~x4 ^ ~x5));
  assign n7852 = (x0 | x1 | x2 | ~x4 | ~x5) & ((~x2 ^ ~x4) | (x0 ? (x1 | ~x5) : (~x1 | x5)));
  assign n7853 = ~n7854 & (~n841 | (~x2 & n7856) | (x2 & n7857));
  assign n7854 = x3 & ((n696 & n746) | (x4 & ~n7855));
  assign n7855 = (x0 | ~x1 | ~x5 | (~x2 ^ x6)) & (x1 | x5 | (x0 ? (~x2 ^ ~x6) : (x2 | ~x6)));
  assign n7856 = (~x6 | ~x7 | ~x3 | ~x5) & (x5 | ((x4 | ~x6 | ~x7) & (x3 | ~x4 | x6 | x7)));
  assign n7857 = (x3 | x4 | x5 | ~x6 | ~x7) & (~x3 | ((x4 | x6 | x7) & (~x6 | ~x7 | ~x4 | ~x5)));
  assign z468 = ~n7859 | n7866 | n7872 | (~n1014 & ~n7871);
  assign n7859 = n7863 & (~n828 | n7860) & (~x4 | n7861);
  assign n7860 = (x0 | ~x1 | ~x2 | x5 | x7) & (x2 | ((x5 | x7 | ~x0 | x1) & (x0 | (x1 ? (~x5 ^ x7) : (~x5 | ~x7)))));
  assign n7861 = (~x5 | x7 | n7862) & (~x7 | ((~n885 | n814) & (x5 | n7862)));
  assign n7862 = (x1 | x2 | ~x3) & (x0 | ~x1 | x3);
  assign n7863 = (n4213 | n7864) & (x7 | ~n570 | n7865);
  assign n7864 = (~x0 | ~x1 | x2) & (x1 | ~x2);
  assign n7865 = (x0 | x3 | ~x4 | ~x5 | x6) & (~x0 | ~x6 | (x3 ? (~x4 | ~x5) : (x4 | x5)));
  assign n7866 = ~x2 & (n7869 | (~x0 & (n7867 | ~n7868)));
  assign n7867 = ~n752 & ~x7 & n1467;
  assign n7868 = (n3345 | n2085) & (~n530 | ~n3408);
  assign n7869 = n841 & ~n7870;
  assign n7870 = x3 ? ((x5 | x6 | x7) & (~x6 | ~x7 | ~x4 | ~x5)) : (~x7 | ((x5 | ~x6) & (~x4 | ~x5 | x6)));
  assign n7871 = ((~x1 ^ ~x6) | (x0 ? (x2 | x3) : ~x3)) & (~x2 | ((x0 | ~x1 | x3 | x6) & (x1 | (~x3 ^ x6))));
  assign n7872 = ~n1008 & (x0 ? ~n7874 : ~n7873);
  assign n7873 = (x4 | (x1 ? ((~x3 | x6) & (~x2 | x3 | ~x6)) : (~x3 ^ ~x6))) & (~x2 | ~x3 | (~x1 ^ x6));
  assign n7874 = (x3 | x6 | ~x1 | x2) & (x1 | x4 | ((~x3 | ~x6) & (~x2 | x3 | x6)));
  assign z469 = ~n7888 | (x4 ? ~n7876 : (n7883 | ~n7885));
  assign n7876 = ~n7877 & ~n7881 & (n643 | n7880);
  assign n7877 = ~x0 & (x1 ? ~n7878 : ~n7879);
  assign n7878 = (~x3 | ((x6 | ~x7 | x2 | x5) & (~x2 | (x5 ? (x6 | ~x7) : (~x6 | x7))))) & (x2 | ~x5 | ((~x6 | ~x7) & (x3 | x6 | x7)));
  assign n7879 = x2 ? ((~x3 | x5 | ~x6 | x7) & (x3 | ~x5 | x6 | ~x7)) : (x3 | ~x7 | (~x5 ^ ~x6));
  assign n7880 = x0 ? ((~x1 | x2 | x3 | ~x5) & (x1 | ~x2 | x5)) : ((~x2 | x3 | x5) & (x1 | ~x3 | (~x2 ^ ~x5)));
  assign n7881 = x0 & ((n943 & n1439) | (~x2 & ~n7882));
  assign n7882 = (~x1 | x3 | x5 | ~x6 | x7) & (x1 | ~x7 | ((~x5 | ~x6) & (~x3 | x5 | x6)));
  assign n7883 = x7 & ((n746 & n2026) | (~x1 & ~n7884));
  assign n7884 = (~x0 | x2 | x3 | ~x5 | ~x6) & ((x2 ? (x5 | ~x6) : (~x5 | x6)) | (x0 ^ x3));
  assign n7885 = (n1701 | n2373) & (x7 | (~n7886 & n7887));
  assign n7886 = n3488 & (x2 ? (~x3 & ~x5) : (~x3 ^ ~x5));
  assign n7887 = (n2466 | ~n6748) & (n538 | (~n712 & ~n7101));
  assign n7888 = ~n7889 & ~n7892 & n7893 & (n823 | n7891);
  assign n7889 = ~x3 & ((n841 & n1417) | (x1 & ~n7890));
  assign n7890 = (~x0 | x2 | x4 | ~x5 | ~x6) & (x0 | ((~x2 | x4 | ~x5 | ~x6) & (x2 | ~x4 | x5 | x6)));
  assign n7891 = (x2 | x4 | x5 | (~x3 ^ ~x6)) & (~x5 | ((x2 | ~x3 | ~x4 | x6) & (~x2 | (x3 ? (x4 | ~x6) : (~x4 | x6)))));
  assign n7892 = n626 & ((n1364 & n1156) | (~x2 & ~n1040));
  assign n7893 = (~n1269 | ~n1203) & (~n696 | ~n837);
  assign z470 = ~n7909 | ~n7904 | n7900 | n7895 | n7898;
  assign n7895 = ~n1097 & (x2 ? ~n7896 : ~n7897);
  assign n7896 = (x0 | ~x3 | x7 | (~x1 & x4)) & (x1 | ((~x0 | (x3 ? (~x4 | x7) : (x4 | ~x7))) & (x0 | x3 | ~x4 | x7)));
  assign n7897 = (~x0 | ~x1 | x3 | x4 | x7) & (x0 | ~x3 | ~x7 | (~x1 ^ ~x4));
  assign n7898 = n543 & (x2 ? (n828 & n951) : ~n7899);
  assign n7899 = (x3 | ~x4 | ~x5 | x6 | x7) & (~x3 | ~x6 | (x4 ? (x5 | x7) : (~x5 | ~x7)));
  assign n7900 = ~n1198 & (n7901 | n7902 | ~n7903);
  assign n7901 = ~x2 & ((n543 & n2047) | (n841 & ~n2017));
  assign n7902 = ~x0 & ~x1 & (x2 ? (x3 & x7) : (~x3 & ~x7));
  assign n7903 = (~n2492 | ~n746) & (~n922 | ~n5758);
  assign n7904 = n7907 & (x1 | n7905) & (n1548 | n7906);
  assign n7905 = (~x0 | ~x2 | ~x3 | x5 | ~x7) & (x0 | ((x2 | ~x3 | ~x5 | x7) & (~x2 | x3 | x5 | ~x7)));
  assign n7906 = (x0 | ~x1 | ~x2 | x5 | ~x7) & (~x0 | ((x2 | x5 | x7) & (x1 | ~x5 | (~x2 ^ x7))));
  assign n7907 = (~n733 | ~n923) & (~n873 | n7908);
  assign n7908 = x2 ? (~x5 | x7) : (~x5 ^ ~x7);
  assign n7909 = x1 | (~n7910 & n7911 & (~n670 | ~n2435));
  assign n7910 = n828 & (x2 ? (x5 & ~x7) : (x0 ? (~x5 & ~x7) : (x5 & x7)));
  assign n7911 = (x5 | n2466 | n1850) & (x2 | ~x5 | n7912);
  assign n7912 = (x0 | x3 | ~x4 | ~x6 | ~x7) & (~x0 | ~x3 | (x4 ? (~x6 | ~x7) : (x6 | x7)));
  assign z471 = n7914 | ~n7922 | (x1 ? ~n7932 : ~n7930);
  assign n7914 = ~x0 & (n7920 | (x6 & (n7915 | ~n7917)));
  assign n7915 = ~x1 & ~n7916;
  assign n7916 = (x2 | ~x3 | ~x4 | x5 | ~x7) & (~x2 | x3 | x7 | (~x4 ^ x5));
  assign n7917 = ~n7919 & (x1 ? (~n902 | ~n670) : n7918);
  assign n7918 = (x2 | x3 | ~x4 | x5) & (~x2 | ~x3 | x4 | ~x5);
  assign n7919 = x5 & ~x4 & x3 & x1 & ~x2;
  assign n7920 = ~x6 & ((n867 & n2135) | (~x2 & ~n7921));
  assign n7921 = (x1 | ~x3 | x4 | ~x5 | x7) & (x3 | ~x4 | x5 | (~x1 & ~x7));
  assign n7922 = ~n7923 & ~n7926 & n7928 & (n647 | n7925);
  assign n7923 = n841 & (x2 ? (n7033 | n7034) : ~n7924);
  assign n7924 = (~x3 | ~x5 | ~x6 | (~x4 ^ ~x7)) & (x6 | (~x3 ^ ~x7) | (x4 ^ ~x5));
  assign n7925 = x0 ? (x6 | ((x2 | x7) & (x1 | (x2 & x7)))) : ((~x1 | x6 | ~x7) & (~x6 | (x1 & (x2 | x7))));
  assign n7926 = ~n1408 & ((n1209 & n4531) | (n3483 & ~n7927));
  assign n7927 = (x1 | x2 | ~x3 | ~x5) & (x3 | x5 | ~x1 | ~x2);
  assign n7928 = x7 ? n7929 : (n1026 | ~n2940);
  assign n7929 = (~x0 | ((x1 | ~x2 | ~x3 | x6) & (~x1 | x2 | x3 | ~x6))) & (x0 | x1 | ~x2 | x3 | x6);
  assign n7930 = (~n5479 | n2017) & (x0 | (n7931 & (~n878 | n2017)));
  assign n7931 = (x2 | x3 | x4 | ~x6 | x7) & (~x2 | ((x6 | x7 | x3 | x4) & (~x3 | ~x4 | (~x6 ^ ~x7))));
  assign n7932 = (~n550 | ~n600) & (x0 | n7933);
  assign n7933 = (~x6 | ~x7 | ~x3 | ~x4) & (x4 | x6 | x2 | x3);
  assign z472 = n7935 | ~n7940 | ~n7942 | (~n1218 & ~n7939);
  assign n7935 = ~x2 & (n7936 | (n681 & ~n7938));
  assign n7936 = x4 & (x7 ? (n1451 & ~n1312) : ~n7937);
  assign n7937 = (~x0 | x3 | x5 | (x1 ^ ~x6)) & (~x3 | ~x5 | ((x1 | ~x6) & (x0 | ~x1 | x6)));
  assign n7938 = (~x0 | x6 | (x1 ? (~x3 | ~x7) : (x3 | x7))) & (x3 | ~x6 | ((~x1 | x7) & (x0 | x1 | ~x7)));
  assign n7939 = x1 ? (x2 | ~x5 | (x0 & x3)) : ((~x3 | x5) & (~x2 | (~x3 & x5)));
  assign n7940 = n7941 & (~x2 | ~n543 | (~n2648 & ~n5212));
  assign n7941 = (~n746 | ~n1598) & (~n560 | ~n2647);
  assign n7942 = (x2 | n7943) & (~n686 | n7945);
  assign n7943 = (~n551 | n3972) & (x0 | (n7944 & (~n1093 | n3972)));
  assign n7944 = (~x1 | ~x3 | ~x4 | x5 | x7) & (x1 | x3 | x4 | ~x5 | ~x7);
  assign n7945 = ((~x4 ^ ~x7) | ((x1 | x6) & (x0 | ~x1 | ~x6))) & (x4 | ~x7 | ((x1 | ~x6) & (x0 | ~x1 | x6)));
  assign z473 = ~n7955 | (x5 ? (n7947 | n7950) : ~n7951);
  assign n7947 = x4 & (n7948 | n7949 | (n1269 & n1135));
  assign n7948 = ~x2 & ((n922 & n1403) | (n626 & ~n5269));
  assign n7949 = ~n823 & ((n902 & n1857) | (x2 & ~n3315));
  assign n7950 = n733 & n828 & n1769;
  assign n7951 = ~n7953 & (~n1585 | ~n1250) & (n823 | n7952);
  assign n7952 = (~x2 | x3 | ~x4 | ~x6 | ~x7) & (x2 | x6 | (x3 ? (~x4 | ~x7) : (x4 | x7)));
  assign n7953 = ~x4 & ((~n1026 & ~n7954) | (n2155 & n816));
  assign n7954 = (x0 | x1 | ~x2 | ~x7) & (x2 | x7 | ~x0 | ~x1);
  assign n7955 = x2 ? (~n7958 & n7959) : (~n7956 & n7957);
  assign n7956 = ~x5 & n1188 & (x0 ? x6 : (x4 & ~x6));
  assign n7957 = (~x5 | ~x6 | x3 | x4) & (x5 | (x3 ? (x6 ? x0 : x4) : (~x4 | x6)));
  assign n7958 = x5 & ((~x0 & ~x1 & ~x6) | ((~x0 | ~x1) & (x3 ^ ~x6)));
  assign n7959 = (x0 & (x1 | x4)) | (x1 & x4) | (~n2026 & (~n624 | (~x0 & ~x1)));
  assign z474 = ~n7971 | (x0 ? ~n7967 : (n7961 | ~n7963));
  assign n7961 = ~x4 & ((n1070 & n2135) | (~x2 & ~n7962));
  assign n7962 = (x1 | ~x3 | x5 | ~x6 | ~x7) & (x3 | ((x6 | ~x7 | x1 | x5) & (~x1 | (x5 ? (x6 | x7) : (~x6 | ~x7)))));
  assign n7963 = ~n7964 & (~x4 | (x3 & n7965) | (~x3 & n7966));
  assign n7964 = ~n1954 & ((n530 & n1029) | (n828 & n813));
  assign n7965 = (~x1 & (x2 | ~x5)) | (x2 & ~x5) | (x6 & ~x7) | (x7 & (~x6 | (x1 & ~x2 & x5)));
  assign n7966 = (~x1 | ((x2 | ~x5 | ~x6 | ~x7) & (~x2 | x5 | x6 | x7))) & (x1 | x2 | x5 | x6 | x7);
  assign n7967 = ~n1505 & (x1 | (~n7448 & ~n7968 & ~n7970));
  assign n7968 = x3 & ~n7969;
  assign n7969 = (x2 | ~x5 | (x4 ? (x6 | x7) : (~x6 | ~x7))) & (~x2 | ~x4 | x5 | ~x6 | ~x7);
  assign n7970 = ~n640 & ((n1121 & n885) | (~n1744 & n934));
  assign n7971 = ~n7972 & n7976 & (n643 | (~n7974 & ~n7975));
  assign n7972 = ~x1 & ((n704 & n549) | (x5 & ~n7973));
  assign n7973 = (x0 | x2 | x3 | x4 | x6) & (~x0 | ((~x4 | ~x6 | x2 | x3) & (~x2 | x4 | (~x3 ^ ~x6))));
  assign n7974 = ~n647 & (~x0 ^ (x1 & ~x2));
  assign n7975 = n1392 & (~n1036 | (~x0 & ~x5 & ~n3802));
  assign n7976 = (n714 | n7977) & (n1011 | n7978);
  assign n7977 = (x3 | x6 | ~x0 | x2) & (~x3 | ~x6 | x0 | ~x2);
  assign n7978 = (x0 | x4 | (~x1 & ~x5)) & (x1 | x5 | (x0 ^ ~x4));
  assign z475 = n7988 | ~n7990 | (x1 ? ~n7985 : ~n7980);
  assign n7980 = x0 ? (~n7984 & (~x2 | n7983)) : n7981;
  assign n7981 = x5 ? (~n885 | (~n1786 & ~n2724)) : n7982;
  assign n7982 = (x2 | ~x3 | x6 | (~x4 ^ ~x7)) & (~x6 | ((~x2 | x3 | x4 | ~x7) & (x2 | (x3 ? (x4 | ~x7) : (~x4 | x7)))));
  assign n7983 = (x3 | x4 | ~x5 | x6 | ~x7) & (~x3 | ~x4 | x5 | ~x6 | x7);
  assign n7984 = x5 & n902 & (x4 ? (x6 ^ ~x7) : (x6 ^ x7));
  assign n7985 = (~n547 | ~n662) & (x5 | (~n7986 & ~n7987));
  assign n7986 = x7 & ((~n1408 & ~n2373) | (n742 & n1331));
  assign n7987 = n683 & (x0 ? (~x2 & n1835) : (x2 & ~n1353));
  assign n7988 = x5 & (x3 ? (n4089 & n1269) : ~n7989);
  assign n7989 = (x0 | ~x1 | x2 | x7) & (~x0 | x1 | (x2 ? (~x4 | x7) : ~x7));
  assign n7990 = ~n7991 & (x5 | (n7994 & (x1 | n7993)));
  assign n7991 = ~n671 & ~n7992;
  assign n7992 = ((~x2 ^ x3) | (x0 ? (x1 | x5) : ~x5)) & (x0 | ~x1 | x2 | ~x3) & (~x5 | (x0 ? (x1 ? (x2 | x3) : (~x2 | ~x3)) : (~x1 ^ ~x3)));
  assign n7993 = (x0 | ~x2 | ((x4 | x7) & (~x3 | ~x4 | ~x7))) & (x2 | x3 | (x0 ? (~x4 ^ ~x7) : (x4 | ~x7)));
  assign n7994 = (~n5388 | n7995) & (n1433 | n3823);
  assign n7995 = x2 ? (x3 ^ ~x7) : (x3 | x7);
  assign z476 = n7997 | ~n8001 | ~n8007 | (x3 & ~n7999);
  assign n7997 = x0 & ((n576 & n1358) | (~x1 & ~n7998));
  assign n7998 = (x5 | ((~x2 | (x3 ? (~x4 | ~x6) : (x4 | x6))) & (x2 | ~x3 | ~x4 | x6))) & (x2 | ~x5 | ~x6 | (~x3 & ~x4));
  assign n7999 = (~n746 | ~n817) & (x6 | ~n1145 | n8000);
  assign n8000 = (~x5 | ~x7 | x0 | ~x2) & (x7 | (x0 ? (~x2 ^ ~x5) : (~x2 | x5)));
  assign n8001 = n8006 & (x1 | n8002) & (x0 | n8003);
  assign n8002 = (x0 | ~x2 | x3 | ~x5) & (~x0 | ((x4 | ~x5 | x2 | x3) & (~x2 | x5 | (~x3 ^ x4))));
  assign n8003 = n8005 & (~n1467 | n8004) & (n1932 | n5950);
  assign n8004 = (x2 | x3 | x4 | ~x6) & (~x2 | ~x3 | ~x4 | x6);
  assign n8005 = (~x1 | x2 | x3 | x5 | x6) & (x1 | ~x2 | ~x3 | ~x5 | ~x6);
  assign n8006 = (n1198 | n5235) & (~n2797 | (~n934 & ~n5525));
  assign n8007 = ~n8008 & (x3 | n8010);
  assign n8008 = ~n1008 & ((n543 & n5244) | (x4 & ~n8009));
  assign n8009 = x0 ? ((x1 | ~x2 | ~x3 | x6) & (~x1 | x2 | x3 | ~x6)) : (x1 | x2 | (~x3 ^ ~x6));
  assign n8010 = (x5 | x7 | n8011) & (~x7 | ((~x5 | n8011) & (~n1167 | n8012)));
  assign n8011 = (x0 | ~x1 | x2 | ~x4 | ~x6) & (~x0 | x1 | (x2 ? (x4 | ~x6) : (~x4 | x6)));
  assign n8012 = (~x5 | ~x6 | ~x1 | x2) & (x1 | x5 | (~x2 ^ ~x6));
  assign z477 = n8018 | n8021 | ~n8023 | (~x1 & ~n8014);
  assign n8014 = x0 ? (~n8017 & (n1555 | ~n859)) : n8015;
  assign n8015 = ~n7695 & (n3770 | n1932) & (x3 | n8016);
  assign n8016 = (~x2 | x6 | ~x7 | (x4 ^ ~x5)) & (x2 | x4 | ~x5 | x7);
  assign n8017 = n1364 & n1084 & (x3 | ~x7);
  assign n8018 = x2 & (~n8020 | (~x7 & ~n8019));
  assign n8019 = (x0 | ~x1 | x3 | ~x4 | ~x6) & (x1 | ((x0 | (x3 ? (x4 | ~x6) : x6)) & (x3 | x4 | x6) & (~x4 | ~x6 | ~x0 | ~x3)));
  assign n8020 = (n3134 | n2527) & (~n699 | ~n1395);
  assign n8021 = n543 & ((n942 & n1556) | ~n7658 | n8022);
  assign n8022 = n1301 & ((n1769 & n859) | (~x2 & ~n3319));
  assign n8023 = ~n8024 & ~n8027 & n8028 & (~n572 | n8026);
  assign n8024 = ~n647 & ~n8025;
  assign n8025 = x1 ? ((x2 | x6 | x7) & (~x6 | ~x7 | x0 | ~x2)) : ((x6 | ((~x2 | ~x7) & (~x0 | (~x2 & ~x7)))) & (x2 | ~x6 | (x0 & x7)));
  assign n8026 = (x0 | x1 | ~x3 | ~x4 | ~x6) & (x3 | ((~x1 | ~x4 | ~x6) & (x0 | (~x1 ^ ~x6))));
  assign n8027 = ~n7918 & (x0 ? (~x1 & ~n643) : (x1 & n1857));
  assign n8028 = (~x3 | ~x4 | n8029) & (x3 | x4 | ~n743 | n1312);
  assign n8029 = (x2 | ~x6 | ~x0 | x1) & (x0 | (x1 ? (x2 | x6) : (~x2 | ~x6)));
  assign z478 = n8039 | ~n8042 | (x0 ? ~n8035 : ~n8031);
  assign n8031 = ~n8032 & (x2 | n8033);
  assign n8032 = ~n3924 & ((~x4 & ~x6 & x1 & x2) | (~x1 & x4 & (x2 ^ ~x6)));
  assign n8033 = (n1198 | n1246 | x3 | x4) & (~x3 | n8034);
  assign n8034 = (~x4 | ((~x6 | ~x7 | x1 | x5) & (x6 | x7 | ~x1 | ~x5))) & (~x1 | x4 | x5 | (~x6 ^ x7));
  assign n8035 = (x2 | n8036) & (x1 | ~x2 | ~x4 | n8038);
  assign n8036 = x6 ? (~n551 | (~n2647 & ~n6035)) : n8037;
  assign n8037 = (~x1 | x5 | (x3 ? (x4 | ~x7) : (~x4 | x7))) & (x1 | x3 | x4 | ~x5 | x7);
  assign n8038 = (x3 | x5 | (~x6 ^ x7)) & (~x3 | ~x5 | x6 | ~x7);
  assign n8039 = ~x1 & (x4 ? ~n8041 : ~n8040);
  assign n8040 = x2 ? (x0 ? (~x3 | (~x5 ^ ~x7)) : (x3 | (~x5 ^ x7))) : ((~x5 | ~x7 | x0 | x3) & (~x0 | x5 | (~x3 ^ ~x7)));
  assign n8041 = (x0 | x2 | ~x7 | (~x3 ^ ~x5)) & (~x2 | ((~x5 | x7 | x0 | ~x3) & (~x0 | (x3 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n8042 = n8045 & (x2 | n8043) & (~n543 | n8044);
  assign n8043 = (x0 | ~x1 | x3 | ~x4 | ~x7) & (x7 | ((x0 | x1 | ~x3 | x4) & (~x0 | (x1 ? (x3 | x4) : (~x3 | ~x4)))));
  assign n8044 = (x5 | (~x2 ^ ~x7) | (~x3 ^ ~x4)) & (~x3 | ~x5 | (x2 ? (~x4 | x7) : (~x4 ^ ~x7)));
  assign n8045 = ~n8046 & (~n743 | ~n3468) & (~n1209 | ~n2647);
  assign n8046 = ~x0 & x2 & (x3 ? (~x4 & x7) : (x4 & ~x7));
  assign z479 = n8053 | ~n8059 | (x2 ? ~n8056 : ~n8048);
  assign n8048 = x5 ? (~n8050 & (x1 | n8049)) : n8051;
  assign n8049 = (x0 | ~x3 | ~x4 | ~x6 | ~x7) & (x7 | ((~x0 | x3 | ~x4 | x6) & ((~x4 ^ ~x6) | (~x0 ^ ~x3))));
  assign n8050 = n543 & (n1526 | (~x3 & n3251));
  assign n8051 = (~n550 | ~n1234) & (x3 | n8052);
  assign n8052 = (~x0 | ~x4 | (x1 ? (x6 | x7) : (~x6 | ~x7))) & (x4 | ((x1 | x6 | ~x7) & (x0 | ~x1 | ~x6 | x7)));
  assign n8053 = ~x1 & ((~x4 & ~n8054) | (n1479 & ~n8055));
  assign n8054 = x3 ? (x0 ? (x5 | x6) : (~x5 | (x2 & x6))) : ((~x2 | (x0 ? (~x5 | ~x6) : (x5 | x6))) & (~x0 | x2 | (~x5 ^ x6)));
  assign n8055 = x0 ? ((~x3 | ~x5) & (~x2 | x3 | x5)) : ((x3 | ~x5) & (x2 | ~x3 | x5));
  assign n8056 = ~n8057 & (~n841 | n6710);
  assign n8057 = ~x0 & (x7 ? ~n8058 : (~n981 & ~n2208));
  assign n8058 = (x1 | x3 | ~x4 | x5 | x6) & (~x1 | ~x3 | x4 | ~x5 | ~x6);
  assign n8059 = n8062 & (~x1 | (~n8060 & ~n8061));
  assign n8060 = ~n1566 & ((n743 & n1835) | (~x0 & n597));
  assign n8061 = n1310 & ((n1044 & n1835) | (x2 & ~n2527));
  assign n8062 = x0 ? (~x6 | n8064) : n8063;
  assign n8063 = x1 ? (x6 | (x2 ? (x3 | ~x5) : (~x3 | x5))) : (~x6 | ((x3 | x5) & (~x2 | ~x3 | ~x5)));
  assign n8064 = (x3 | ~x5 | ~x1 | x2) & (x1 | ~x3 | x5);
  assign z480 = n8066 | n8071 | ~n8075 | (~n1850 & ~n8074);
  assign n8066 = ~x7 & (n8067 | (n1012 & ~n8070));
  assign n8067 = ~x4 & (x6 ? ~n8068 : ~n8069);
  assign n8068 = (x0 | ~x1 | x2 | x3 | ~x5) & (~x0 | x1 | ~x2 | ~x3 | x5);
  assign n8069 = (x0 | ~x1 | (~x2 & (~x3 | x5))) & (x1 | ((x2 | x3 | ~x5) & (~x0 | ((x3 | ~x5) & (x2 | (x3 & ~x5))))));
  assign n8070 = (x2 | ((x5 | ~x6) & (~x3 | ~x5 | x6))) & (~x6 | ((x3 | x5) & (~x2 | ~x3 | ~x5)));
  assign n8071 = x7 & ((~n1353 & ~n8072) | (n1686 & ~n8073));
  assign n8072 = (~x0 | x1 | x2 | x3 | ~x5) & (x0 | ~x1 | x5 | (~x2 ^ x3));
  assign n8073 = (x1 | x2 | x3 | x4 | ~x5) & (~x1 | ~x4 | ((~x2 | (~x3 & ~x5)) & (~x3 | ~x5) & (x2 | x3 | x5)));
  assign n8074 = (~x0 | x3 | (x1 ? (x2 | ~x5) : (~x2 | x5))) & (x1 | ((x2 | ~x3 | x5) & (x0 | (x2 ? (~x3 | ~x5) : x5))));
  assign n8075 = (n2803 | n8079) & (n643 | (~n8076 & n8077));
  assign n8076 = ~x3 & ((n841 & n3509) | (~x0 & ~n5769));
  assign n8077 = ~n8078 & (n6891 | ~n3711) & (n1934 | ~n2797);
  assign n8078 = ~x4 & ((x0 & x1 & ~x2 & ~x5) | (~x0 & x2 & (x1 ^ ~x5)));
  assign n8079 = (~x2 & ((~x1 & ~x3 & x5) | (x0 & (x3 ? x5 : ~x1)))) | (x1 & (x2 | x3 | (~x0 & ~x5)));
  assign z481 = n8086 | ~n8094 | (~x1 & (~n8081 | ~n8089));
  assign n8081 = x3 ? n8084 : (~n8083 & (~x5 | n8082));
  assign n8082 = (x0 | ~x2 | x6 | ~x7) & (~x0 | ((~x4 | ~x6 | x7) & (x2 | (x4 ? ~x6 : (x6 | ~x7)))));
  assign n8083 = n757 & ((~x4 & x6 & x0 & ~x2) | (~x0 & (x2 ? x6 : (~x4 & ~x6))));
  assign n8084 = (x0 | ~n978 | ~n1084) & (~n6842 | n8085);
  assign n8085 = (~x6 & (~x5 | (~x0 & x4))) | (x5 & x6) | (x0 & ~x4);
  assign n8086 = ~n1097 & ((~n697 & ~n8087) | (~x7 & ~n8088));
  assign n8087 = (~x0 | x1 | ~x3 | x4) & (x0 | ~x1 | x3 | ~x4);
  assign n8088 = (x0 | ~x1 | ~x2 | x4) & (x1 | ((~x3 | ~x4 | ~x0 | ~x2) & (x0 | (x2 ? x3 : (~x3 | ~x4)))));
  assign n8089 = n8091 & (x5 | n8090);
  assign n8090 = (~x0 | ~x2 | ~x3 | x4 | ~x7) & (x2 | ((x4 | ~x7 | x0 | ~x3) & (~x4 | (x0 ? (~x3 ^ ~x7) : (x3 | ~x7)))));
  assign n8091 = ~n8093 & (~n1986 | n4336) & (n605 | n8092);
  assign n8092 = (x4 | x7 | ~x0 | x3) & (~x4 | ~x7 | x0 | ~x3);
  assign n8093 = x0 & ((~x2 & x3 & x5 & ~x7) | (x2 & ~x3 & ~x5 & x7));
  assign n8094 = ~x1 | (n8095 & ~n8097 & (~n588 | ~n600));
  assign n8095 = (x2 | n8096) & (~n6127 | (~n1465 & ~n3090));
  assign n8096 = (x7 | ((x0 | ~x5 | (~x3 & ~x4)) & (x5 | (x0 ? (x3 ^ ~x4) : (x3 | x4))))) & (x0 | ~x7 | (x3 ? x5 : (x4 | ~x5)));
  assign n8097 = x7 & ((~n1198 & ~n2373) | (n1358 & n1783));
  assign z482 = n8106 | ~n8109 | (~x2 & (~n8099 | ~n8103));
  assign n8099 = x4 ? (~n8100 & (~n1301 | n4587)) : n8101;
  assign n8100 = ~x6 & ~x5 & ~x3 & x0 & ~x1;
  assign n8101 = (x7 | n8102) & (x3 | ~x7 | ~n626 | n1198);
  assign n8102 = (x0 | x1 | ~x5 | (~x3 ^ ~x6)) & (x5 | ((x0 | x1 | ~x3 | x6) & (~x1 | (x0 ? (~x3 ^ x6) : (x3 | x6)))));
  assign n8103 = x0 ? n8104 : n8105;
  assign n8104 = (x1 | ~x3 | ~x4 | x6 | x7) & (~x1 | x3 | x4 | ~x6 | ~x7);
  assign n8105 = (x1 | ~x3 | ~x4 | ~x6 | x7) & (x6 | ((~x1 | (~x3 & (x4 | ~x7))) & (x1 | x3 | ~x4) & (~x3 | ~x7)));
  assign n8106 = x2 & (n8107 | (n543 & n4972 & ~n8108));
  assign n8107 = ~x1 & ((n825 & n1358) | (x0 & ~n7278));
  assign n8108 = x3 ? (x5 | ~x6) : (~x5 ^ ~x6);
  assign n8109 = ~n8110 & (~x2 | (~n8113 & n8114));
  assign n8110 = ~n640 & ((n743 & ~n8112) | (~x0 & ~n8111));
  assign n8111 = (~x2 | ~x3 | (x1 ^ (x4 & x5))) & (~x1 | x2 | x3 | (~x4 & ~x5));
  assign n8112 = x4 ? (x3 | (~x1 & ~x5)) : x1;
  assign n8113 = ~n643 & (x0 ? (~x1 & ~n1548) : (x1 & n828));
  assign n8114 = ~n8115 & (~n699 | ~n1585) & (~n543 | ~n1141);
  assign n8115 = ~x1 & (x0 ? (x3 ? (x4 & x6) : (~x4 & ~x6)) : (~x3 & x6));
  assign z483 = n8117 | ~n8120 | (x1 ? ~n8130 : ~n8129);
  assign n8117 = x2 & (n8118 | (n5257 & n2797));
  assign n8118 = ~x1 & ((~x0 & n8119) | (n2337 & ~n5085));
  assign n8119 = x6 & ((x3 & x4 & x5 & ~x7) | (~x3 & (x4 ? (x5 & x7) : (~x5 & ~x7))));
  assign n8120 = (~x2 & n8121 & ~n8124 & n8125) | (x2 & n8127);
  assign n8121 = (n1558 | n8122) & (~n1411 | n8123);
  assign n8122 = (x0 | x1 | x4 | ~x6) & (~x0 | x6 | (x1 ^ ~x4));
  assign n8123 = (x3 | x4 | ~x6 | ~x7) & (~x3 | ~x4 | (~x6 ^ ~x7));
  assign n8124 = ~n765 & ((~x0 & ~x1 & x3 & ~x4) | (x0 & ~x3 & (x1 ^ x4)));
  assign n8125 = (~n674 | ~n712) & (~n1310 | n8126);
  assign n8126 = (x1 | x3 | x4 | ~x7) & (~x1 | ~x3 | ~x4 | x7);
  assign n8127 = (x1 | n8128) & (~n1012 | (~n2575 & ~n4042));
  assign n8128 = (x0 | ((x3 | x4 | ~x5 | x7) & (x5 | ~x7 | ~x3 | ~x4))) & (~x0 | ~x3 | x4 | x5 | ~x7);
  assign n8129 = x7 ? (x0 ? (x2 ? (x3 | ~x4) : x4) : (~x3 | (~x2 ^ x4))) : (x0 ? (~x2 | (~x3 ^ ~x4)) : (x3 | ~x4));
  assign n8130 = (x0 | x4 | ((~x3 | x7) & (~x2 | x3 | ~x7))) & (x2 | ((x3 | ~x4 | ~x7) & (x0 | x4 | x7)));
  assign z484 = ~n8132 | n8138 | ~n8140 | (~x0 & ~n8136);
  assign n8132 = (n1011 | n8135) & (~x2 | n8133) & (x2 | n8134);
  assign n8133 = (x1 | (x0 ? (x4 | (~x3 ^ x5)) : (~x4 | x5))) & (x0 | ((x3 | ~x4 | x5) & (x4 | ~x5 | ~x1 | ~x3)));
  assign n8134 = (~x0 | x4 | (x1 ? (x3 | x5) : ~x5)) & (~x4 | ((~x1 | x3 | ~x5) & (x0 | (x1 ? (~x3 | x5) : ~x5))));
  assign n8135 = (~x4 | x5 | x7 | ~x0 | x1) & (x0 | x4 | (x1 ? (~x5 | ~x7) : (x5 | x7)));
  assign n8136 = ~n8137 & (~x2 | (~n3403 & (~n1294 | ~n3711)));
  assign n8137 = n1044 & (x1 ? ~n2128 : (~x4 & n962));
  assign n8138 = n564 & ((n978 & n1439) | (~x2 & ~n8139));
  assign n8139 = (x1 | x3 | x5 | x6 | ~x7) & (~x1 | x7 | (x3 ? (x5 | ~x6) : (~x5 | x6)));
  assign n8140 = x1 ? n8143 : (x4 ? n8142 : n8141);
  assign n8141 = (~x0 | ((x3 | x5 | ~x6) & (~x2 | ~x3 | ~x5 | x6))) & (x5 | ~x6 | x2 | x3) & (x0 | ~x3 | (x2 ? (~x5 | ~x6) : (x5 | x6)));
  assign n8142 = (x0 | ~x2 | x3 | ~x5 | x6) & (~x3 | ((~x0 | (x2 ? (~x5 | ~x6) : (x5 | x6))) & (x0 | x2 | x5 | ~x6)));
  assign n8143 = (~n696 | ~n594) & (x0 | n8144);
  assign n8144 = x2 ? ((~x5 | ~x6 | x3 | x4) & (x5 | x6 | ~x3 | ~x4)) : ((~x3 | ~x4 | ~x5 | x6) & (x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))));
  assign z485 = ~n8149 | ~n8156 | ~n8160 | (~x4 & ~n8146);
  assign n8146 = ~n8148 & (~x1 | (~n8147 & (~n742 | ~n4976)));
  assign n8147 = ~x2 & (x0 ? n2660 : (~x3 & n992));
  assign n8148 = n841 & n1051 & ((x5 & x7) | (~x2 & ~x5 & ~x7));
  assign n8149 = ~n8150 & ~n8153 & ~n8154 & (x2 | n8152);
  assign n8150 = ~n1134 & ~n8151;
  assign n8151 = (x0 | ~x1 | x2 | x3 | ~x6) & (~x0 | x1 | (x2 ? (x3 | x6) : (~x3 | ~x6)));
  assign n8152 = x0 ? (x5 | (x1 ? (x3 | ~x6) : (~x3 | x6))) : (~x3 | ~x5 | (x1 ^ ~x6));
  assign n8153 = ~n627 & ((x2 & x5 & x0 & ~x1) | (~x0 & ~x5 & (x1 ^ ~x2)));
  assign n8154 = ~n8155 & n1479 & n622;
  assign n8155 = (x5 | ~x7 | ~x1 | x2) & (x1 | x7 | (x2 ^ ~x5));
  assign n8156 = x2 ? (x0 | n8159) : (~n8157 & ~n8158);
  assign n8157 = n564 & ((n1364 & n689) | (n904 & n927));
  assign n8158 = n566 & ((n904 & n689) | (x1 & ~n975));
  assign n8159 = (x1 | (x3 ? (x4 ? (x5 | ~x6) : (~x5 | x6)) : (~x5 | (~x4 ^ x6)))) & (~x1 | ~x3 | ~x4 | ~x5 | ~x6);
  assign n8160 = ~n8162 & (n3309 | (~n8161 & (~n592 | ~n712)));
  assign n8161 = ~x0 & (x1 ? ~n2693 : n5846);
  assign n8162 = ~n697 & (x0 ? (n577 & n1188) : ~n8163);
  assign n8163 = (~x3 | ((~x5 | x6 | x1 | ~x4) & (x5 | ~x6 | ~x1 | x4))) & (x1 | x3 | (x4 ? (~x5 | ~x6) : (x5 | x6)));
  assign z486 = ~n8173 | ~n8172 | n8170 | n8165 | n8167;
  assign n8165 = ~x2 & (n8166 | (n3687 & n1244));
  assign n8166 = x3 & ((n657 & n951) | (x0 & ~n7092));
  assign n8167 = ~n640 & (~n8169 | (~x3 & ~n8168));
  assign n8168 = (x4 | (~x1 ^ ~x5) | (x0 ^ ~x2)) & (~x0 | ~x4 | x5 | (x1 ^ ~x2));
  assign n8169 = (~x0 | x1 | x3 | x4 | ~x5) & (x0 | ((x1 | ~x3 | ~x4 | ~x5) & (~x1 | x3 | x4 | x5)));
  assign n8170 = x3 & (~n8171 | (~x6 & n859 & ~n3394));
  assign n8171 = (~x0 | x1 | x4 | x5 | ~x6) & (x0 | ~x4 | x6 | (~x1 ^ ~x5));
  assign n8172 = (~n1621 | ~n5198) & (n714 | n643 | ~n1365);
  assign n8173 = ~n8176 & (x3 | (~n8174 & (~x6 | n8175)));
  assign n8174 = ~n1954 & (x0 ? ~n2819 : (x6 & ~n714));
  assign n8175 = (x0 | x1 | x2 | x4 | ~x5) & (~x4 | ((x0 | ~x1 | (~x2 & ~x5)) & (x1 | x2 | (~x0 & x5))));
  assign n8176 = ~x0 & ((~x7 & ~n8177) | (x3 & n1395));
  assign n8177 = (~x1 | ((~x3 | x4 | ~x6) & (x3 | ~x4 | x5 | x6))) & (~x3 | x4 | x5 | ~x6) & (x1 | x3 | ~x5 | (~x4 ^ ~x6));
  assign z487 = n8184 | ~n8185 | ~n8190 | (~x7 & ~n8179);
  assign n8179 = n8182 & (x0 | (~n8181 & (x5 | n8180)));
  assign n8180 = (x1 | x2 | x3 | x4 | ~x6) & (~x1 | ((x2 | x3 | ~x4 | x6) & (x4 | ~x6 | ~x2 | ~x3)));
  assign n8181 = n551 & ((~n1353 & ~n5064) | (n885 & n1835));
  assign n8182 = (~n1209 | ~n1643) & (n1408 | n8183);
  assign n8183 = (~x0 | x1 | x2 | ~x3 | ~x5) & (x0 | ~x1 | x5 | (~x2 ^ x3));
  assign n8184 = ~n823 & (x2 ? (x3 & n809) : (~x3 & ~n3266));
  assign n8185 = ~n8187 & ~n8188 & n8189 & (n2227 | n8186);
  assign n8186 = (~x0 | x1 | x4 | x5 | ~x7) & (x0 | ~x1 | ~x5 | (~x4 ^ ~x7));
  assign n8187 = ~n765 & (n2369 | (~x1 & ~n1010 & ~n2737));
  assign n8188 = ~n2737 & n566 & ~x5 & x7;
  assign n8189 = (~n923 | ~n1269) & (~n600 | ~n809);
  assign n8190 = ~n8191 & (~n572 | (~n8193 & (~n696 | ~n1234)));
  assign n8191 = x7 & ((~n3275 & n5017) | (x4 & ~n8192));
  assign n8192 = (x0 | ~x1 | ~x2 | ~x3 | ~x5) & (x3 | x5 | x1 | x2);
  assign n8193 = n653 & (x1 ? ~n1100 : n2720);
  assign z488 = n8198 | ~n8203 | (~x6 & (~n8195 | ~n8202));
  assign n8195 = x2 ? (x7 | n8197) : n8196;
  assign n8196 = (x3 | x5 | ~x0 | ~x1) & (~x7 | ((x5 | (x1 ^ ~x3)) & (x0 | ~x5 | (~x1 ^ ~x3))));
  assign n8197 = (~x0 | x1 | ~x3 | x5) & (x0 | (x1 ? (~x3 ^ ~x5) : (x3 | ~x5)));
  assign n8198 = ~x2 & (n8200 | (~n643 & ~n8199));
  assign n8199 = (x0 | ~x1 | x3 | ~x4 | ~x5) & (~x0 | x4 | (x1 ? (~x3 | x5) : (x3 | ~x5)));
  assign n8200 = ~x4 & ((n543 & n2026) | (x0 & ~n8201));
  assign n8201 = (~x1 | ~x3 | x5 | x6 | x7) & (x1 | x3 | ~x5 | ~x6 | ~x7);
  assign n8202 = (x1 | (x2 ? (x5 | ~x7) : (~x5 | x7))) & (x0 | ~x1 | (x2 ? (~x5 | ~x7) : (x5 | x7)));
  assign n8203 = n8205 & (~n1156 | ~n1857 | n8204);
  assign n8204 = (x3 | ~x5 | ~x0 | x1) & (x0 | ~x3 | (~x1 ^ x5));
  assign n8205 = ~x6 | (n8206 & (x2 | n8207));
  assign n8206 = (x1 | ~x2 | x5) & (x0 | (x1 ? (~x5 | (~x2 & ~x7)) : x5));
  assign n8207 = (x0 | ~x1 | ~x3 | ~x5 | x7) & (~x0 | x5 | (x1 ^ ~x3));
  assign z489 = n8209 | n8213 | ~n8217 | (~x1 & ~n8216);
  assign n8209 = ~x7 & ((~x5 & ~n8210) | (n5223 & ~n8212));
  assign n8210 = (~x0 | x2 | ~x6 | n1820) & (~x2 | x6 | n8211);
  assign n8211 = (x3 | ~x4 | ~x0 | x1) & (x0 | ~x3 | (~x1 ^ x4));
  assign n8212 = (x4 | x6 | x0 | x2) & (~x4 | ~x6 | ~x0 | ~x2);
  assign n8213 = ~x7 & ((n543 & n8214) | (~x1 & ~n8215));
  assign n8214 = ~x2 & ~x3 & (x4 ^ x6);
  assign n8215 = (x0 | ~x2 | ~x3 | (~x4 ^ ~x6)) & (x3 | ((~x0 | x4 | (x2 ^ ~x6)) & (x0 | x2 | ~x4 | x6)));
  assign n8216 = (~x3 | ((~x2 | ~x6 | ~x7) & (~x0 | (x2 ? ~x6 : (x6 | x7))))) & (x2 | x3 | ~x7 | (x0 ^ x6));
  assign n8217 = n8218 & (~n1283 | ~n4033) & (n2227 | n6571);
  assign n8218 = (~n3236 | n2373) & (~n1300 | ~n1392 | ~n733);
  assign z490 = n8220 | ~n8224 | ~n8228 | (~x1 & ~n8223);
  assign n8220 = x4 & (n8221 | (n1269 & n2409));
  assign n8221 = ~x3 & ((n733 & n951) | (x6 & ~n8222));
  assign n8222 = (x0 | ~x1 | x2 | x5 | x7) & (~x0 | x1 | (x2 ? (x5 | ~x7) : (~x5 | x7)));
  assign n8223 = (x0 | ~x3 | ~x4 | (~x2 ^ ~x7)) & (x4 | ((x0 | ~x2 | ~x3 | x7) & (~x0 | x3 | (x2 ^ ~x7))));
  assign n8224 = ~n8225 & ~n8226 & ~n8227 & (~n543 | ~n3493);
  assign n8225 = x1 & ((~x3 & x7 & x0 & ~x2) | (~x0 & ~x7 & (x2 ^ x3)));
  assign n8226 = ~x1 & (x0 ? (x3 & (x2 ^ ~x7)) : (~x3 & (x2 ^ x7)));
  assign n8227 = ~n697 & n841 & ~x5 & n1392;
  assign n8228 = x5 ? n8229 : (~n774 | n8231);
  assign n8229 = x0 ? (~n570 | ~n3468) : n8230;
  assign n8230 = (x1 | x2 | ~x3 | x4 | x7) & (~x1 | ((x2 | x3 | ~x4 | x7) & (x4 | ~x7 | ~x2 | ~x3)));
  assign n8231 = (~x0 | ~x1 | x2 | x6 | ~x7) & (x0 | ((x1 | x2 | ~x6 | x7) & (~x1 | ~x2 | (~x6 ^ ~x7))));
  assign z491 = n8233 | n8236 | n8241 | (x0 & ~n8239);
  assign n8233 = ~x2 & (n8234 | (n610 & n661));
  assign n8234 = ~x4 & ((n653 & n4831) | (x3 & ~n8235));
  assign n8235 = (x0 | x1 | x5 | x6 | x7) & (~x0 | ~x6 | (x1 ? (x5 | x7) : (~x5 | ~x7)));
  assign n8236 = ~x0 & (x1 ? ~n8237 : ~n8238);
  assign n8237 = (~x2 | (x3 & (x4 | x5 | x6))) & (~x4 | ((x3 | x5 | x6) & (x2 | ~x3 | ~x5 | ~x6)));
  assign n8238 = x3 ? (~x2 | x4) : (~x4 & ((~x5 & ~x6) | (x2 & (~x5 | ~x6))));
  assign n8239 = ~n1917 & ~n4862 & n8240 & (~n828 | ~n570);
  assign n8240 = x1 ? (x2 | x3) : ((x3 | n2760) & (x2 | ~x3 | ~x4));
  assign n8241 = n570 & ((n943 & n5168) | (x4 & ~n8242));
  assign n8242 = (x0 | ~x3 | x5 | x6 | x7) & (~x0 | ~x6 | (x3 ? (~x5 | ~x7) : (x5 | x7)));
  assign z492 = n8244 | ~n8249 | ~n8253 | (~x2 & ~n8247);
  assign n8244 = n570 & (x3 ? ~n8246 : ~n8245);
  assign n8245 = x0 ? (x5 | (x4 ? (~x6 | x7) : (x6 | ~x7))) : (~x5 | (x4 ? (~x6 | ~x7) : (x6 | x7)));
  assign n8246 = (x0 | ~x4 | x5 | x6 | x7) & (~x0 | ~x5 | (x4 ? (~x6 | x7) : (x6 | ~x7)));
  assign n8247 = (x1 | ~x5 | n8248) & (x5 | ((n3098 | ~n1922) & (~x1 | n8248)));
  assign n8248 = (x0 | x3 | x4 | ~x6 | ~x7) & (~x0 | ((~x3 | x4 | ~x6 | x7) & (x3 | ~x4 | x6 | ~x7)));
  assign n8249 = ~n8250 & n8251 & (n1036 | n3133);
  assign n8250 = ~x0 & ((x4 & x5 & x1 & x2) | (~x1 & (x2 ? (~x4 & ~x5) : (x4 & x5))));
  assign n8251 = ~n8252 & (~n959 | ~n837) & (~n746 | ~n1203);
  assign n8252 = ~x5 & ~x4 & ~x2 & x0 & ~x1;
  assign n8253 = ~n8254 & (n877 | n8256) & (x0 | n8255);
  assign n8254 = n743 & ((~n752 & ~n2290) | (n689 & n728));
  assign n8255 = x1 ? ((~x2 | x3 | ~x4 | x5) & (x2 | ~x3 | x4 | ~x5)) : ((x2 | x3 | ~x4 | x5) & (x4 | ~x5 | ~x2 | ~x3));
  assign n8256 = (x0 | ~x1 | x2 | ~x4 | x6) & (~x0 | x1 | ~x2 | (~x4 ^ x6));
  assign z493 = ~n8261 | ~n8266 | (x1 & (n8258 | n8259));
  assign n8258 = ~n615 & ((n743 & n1429) | (n526 & n742));
  assign n8259 = ~x0 & (x2 ? (n828 & n1070) : ~n8260);
  assign n8260 = (~x3 | ~x4 | x5 | x6 | ~x7) & (x3 | ~x6 | ((~x5 | ~x7) & (x4 | x5 | x7)));
  assign n8261 = n8264 & (~x4 | (~n8263 & (x0 | n8262)));
  assign n8262 = (x1 | x3 | ~x5 | (x2 ^ ~x6)) & (~x3 | ((x1 | x2 | x5 | x6) & (~x1 | (x2 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n8263 = n841 & ((n1364 & n902) | (x2 & n4604));
  assign n8264 = x1 ? n8265 : (~n5326 & (~n742 | ~n3847));
  assign n8265 = (~x0 | x2 | x3 | ~x5 | ~x6) & (x0 | (x2 ? (x3 ? (x5 | x6) : (~x5 | ~x6)) : (x5 | (~x3 ^ ~x6))));
  assign n8266 = ~n8267 & (x1 | (~n8271 & (n1353 | n8270)));
  assign n8267 = ~x4 & (x2 ? ~n8269 : ~n8268);
  assign n8268 = (~x0 | ((x1 | x5 | ~x6) & (x3 | ~x5 | x6))) & (x5 | x6 | ~x1 | ~x3) & (x1 | ~x6 | ((x3 | x5) & (x0 | ~x3 | ~x5)));
  assign n8269 = (x0 | ~x1 | x3 | ~x5 | x6) & (x1 | (x0 ? (x3 ? (x5 | x6) : (~x5 | ~x6)) : (x6 | (~x3 ^ ~x5))));
  assign n8270 = (~x0 | x2 | x3 | x5 | ~x7) & (x7 | ((x0 | x2 | ~x3 | x5) & (~x2 | (x0 ? (~x3 ^ ~x5) : (x3 | ~x5)))));
  assign n8271 = ~x7 & ((n926 & n2435) | (n691 & ~n8272));
  assign n8272 = (~x0 | (x3 ? (x4 | ~x6) : (~x4 | x6))) & (x0 | x3 | x4 | ~x6);
  assign z494 = ~n8284 | ~n8281 | n8274 | n8278;
  assign n8274 = ~x0 & (n8275 | (n1857 & ~n8277));
  assign n8275 = x7 & ((n558 & n696) | (x6 & ~n8276));
  assign n8276 = (~x1 | ~x3 | (x2 ? (~x4 | ~x5) : (x4 | x5))) & (x3 | ((~x1 | ~x2 | ~x4 | x5) & (x1 | (x2 ? (x4 | x5) : ~x4))));
  assign n8277 = (~x4 | ~x5 | ~x1 | x3) & (x1 | x4 | ((x3 | ~x5) & (x2 | ~x3 | x5)));
  assign n8278 = ~n643 & (~n8280 | (~x2 & ~n8279));
  assign n8279 = (x4 | ((x0 | x1 | x3 | ~x5) & (~x0 | ~x3 | (x1 ^ ~x5)))) & (x0 | ~x4 | (x1 ? (x3 | ~x5) : x5));
  assign n8280 = (~n959 | ~n1269) & (n1580 | (~n934 & ~n1194));
  assign n8281 = ~n8282 & (n1040 | n1766) & (n1282 | n2953);
  assign n8282 = x6 & ((n746 & n1641) | (x5 & ~n8283));
  assign n8283 = (x0 | ((~x3 | ~x4 | x1 | x2) & (~x1 | x3 | x4))) & (~x0 | x1 | ~x2 | x3 | ~x4);
  assign n8284 = ~n8285 & (~n841 | (x3 & n8288) | (~x3 & n8289));
  assign n8285 = ~x6 & ((~x0 & ~n8286) | (n841 & ~n8287));
  assign n8286 = x1 ? ((x2 | ~x4 | (~x3 ^ ~x5)) & (x4 | x5 | ~x2 | ~x3)) : ((~x2 | x3 | ~x4 | x5) & (x2 | ~x3 | x4 | ~x5));
  assign n8287 = x3 ? (x5 | (x2 ^ x4)) : (x4 | ~x5);
  assign n8288 = (x2 | ~x4 | ~x6 | ~x7) & (x4 | ((~x5 | x6 | x7) & (~x6 | ~x7 | ~x2 | x5)));
  assign n8289 = (x2 | ~x4 | ~x5 | ~x6 | ~x7) & (x6 | x7 | x4 | x5);
  assign z495 = ~n8299 | (x5 ? ~n8295 : ~n8291);
  assign n8291 = x0 ? n8294 : (x1 ? n8292 : n8293);
  assign n8292 = (~x2 | x3 | ~x4 | (~x6 ^ x7)) & (~x3 | ((x6 | ~x7 | ~x2 | x4) & (x2 | ((~x6 | ~x7) & (x4 | x6 | x7)))));
  assign n8293 = (~x7 | (x2 ? (x3 ? (~x4 | ~x6) : (x4 | x6)) : (~x6 | (x3 ^ ~x4)))) & (~x4 | x6 | x7 | (~x2 ^ ~x3));
  assign n8294 = (~n1397 | n3042) & (~n2674 | ~n3818);
  assign n8295 = (x1 | n8296) & (x0 | ~x1 | n8298);
  assign n8296 = x2 ? (~n1861 & (~x0 | n1862)) : n8297;
  assign n8297 = (~x0 | ((~x4 | ~x6 | x7) & (x6 | ~x7 | x3 | x4))) & (~x4 | x7 | ((x3 | ~x6) & (x0 | ~x3 | x6)));
  assign n8298 = (~x6 | ((x2 | ~x3 | x4 | x7) & (~x4 | (x2 ? (x3 ^ ~x7) : (x3 | x7))))) & (x4 | x6 | (x2 ? (x3 | x7) : ~x7));
  assign n8299 = ~n8300 & n8304 & (~n543 | n8303);
  assign n8300 = ~x1 & (~n8302 | (~x5 & ~n8301));
  assign n8301 = (x0 | ~x2 | ~x3 | x4 | ~x7) & (x2 | ((~x4 | x7 | x0 | ~x3) & (~x0 | (x3 ? (x4 | ~x7) : (~x4 | x7)))));
  assign n8302 = (~x0 | ~x2 | x3 | x5 | x7) & (x0 | ~x5 | (x2 ? (x3 | x7) : (~x3 | ~x7)));
  assign n8303 = (x5 | x7 | x3 | x4) & (~x4 | ((x2 | ~x3 | ~x5 | ~x7) & (~x2 | (x3 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n8304 = (n1205 | n8305) & (n1850 | n8306);
  assign n8305 = x0 ? ((~x1 | x2 | x4 | x5) & (x1 | ~x2 | ~x5)) : ((x4 | x5 | x1 | x2) & (~x1 | (x2 ? (x4 | ~x5) : (~x4 | x5))));
  assign n8306 = (~x0 | ~x1 | x2 | x3 | ~x5) & (x1 | ((~x3 | ~x5 | x0 | ~x2) & ((~x2 ^ x5) | (x0 ^ x3))));
  assign z496 = n8320 | ~n8323 | (x5 ? ~n8314 : ~n8308);
  assign n8308 = ~n8309 & (~n560 | ~n1525) & (x0 | n8311);
  assign n8309 = ~n640 & ~n8310;
  assign n8310 = (x0 | ~x1 | x2 | ~x3 | ~x4) & (x1 | ((x0 | x2 | ~x3 | x4) & (~x2 | (x0 ? (~x3 ^ ~x4) : (x3 | ~x4)))));
  assign n8311 = (x4 | n8313) & (~x6 | ~n8312 | ~x3 | ~x4);
  assign n8312 = ~x7 & (x1 ^ ~x2);
  assign n8313 = x1 ? ((~x6 | ~x7 | ~x2 | ~x3) & (x6 | x7 | x2 | x3)) : ((~x2 | ~x3 | ~x6 | x7) & (x6 | ~x7 | x2 | x3));
  assign n8314 = x1 ? n8318 : (~n8315 & n8316);
  assign n8315 = ~n3309 & (n6063 | (x0 & ~n615));
  assign n8316 = (~x4 | n8317) & (x3 | x4 | ~n1181 | n643);
  assign n8317 = (x0 | x2 | ~x3 | x6 | ~x7) & (~x0 | ~x2 | x3 | ~x6 | x7);
  assign n8318 = (~n2435 | ~n1585) & (x3 | n8319);
  assign n8319 = (~x0 | x2 | ~x4 | ~x6 | ~x7) & ((x0 ? (x2 | x4) : (x2 ^ ~x4)) | (~x6 ^ x7));
  assign n8320 = x5 & (x6 ? ~n8322 : ~n8321);
  assign n8321 = ((~x3 ^ ~x4) | (x0 ? (x1 | ~x2) : (~x1 | x2))) & (x0 | ((~x1 | ~x2 | ~x3 | x4) & (x1 | (x2 ? (x3 | ~x4) : (~x3 | x4)))));
  assign n8322 = (x0 | ~x1 | x2 | ~x3 | x4) & (x1 | ((~x3 | ~x4 | ~x0 | x2) & (x0 | (x2 ? (~x3 | x4) : (x3 | ~x4)))));
  assign n8323 = ~n8328 & (x5 | (~n8324 & ~n8326 & n8327));
  assign n8324 = ~x0 & ~n8325;
  assign n8325 = (~x2 | ((~x1 | ~x3 | ~x4 | x6) & (x4 | ~x6 | x1 | x3))) & (x1 | x2 | ~x4 | (~x3 ^ x6));
  assign n8326 = ~n615 & ~n1036;
  assign n8327 = (~n560 | ~n744) & (n1353 | ~n3416);
  assign n8328 = ~n627 & ((~n4233 & n8329) | (n717 & n746));
  assign n8329 = ~x4 & (x0 ^ x2);
  assign z497 = n8337 | ~n8341 | (x3 ? ~n8334 : ~n8331);
  assign n8331 = ~n8333 & (~n733 | ~n809) & (~x7 | n8332);
  assign n8332 = (x0 | ~x1 | x2 | ~x4 | ~x5) & (x1 | ((x4 | ~x5 | x0 | x2) & (~x2 | (x0 ? (~x4 ^ ~x5) : (~x4 | x5)))));
  assign n8333 = ~n1998 & (x1 ? ~n1014 : n607);
  assign n8334 = ~n8335 & ~n8336 & (~n560 | ~n867);
  assign n8335 = n566 & ((~x5 & ~x7 & ~x1 & x2) | (x7 & (x1 ? (x2 ^ ~x5) : (~x2 & x5))));
  assign n8336 = ~n1008 & ((n841 & n859) | (~n3802 & n1167));
  assign n8337 = ~n640 & (n8338 | ~n8340 | (~n856 & ~n1036));
  assign n8338 = ~x0 & ~n8339;
  assign n8339 = (~x2 | ((~x1 | ~x3 | ~x4 | x5) & (x4 | ~x5 | x1 | x3))) & (x1 | x2 | ~x4 | (~x3 ^ x5));
  assign n8340 = (~n560 | ~n1311) & (n1134 | ~n3416);
  assign n8341 = ~n8345 & (x2 | (~n8342 & ~n8343 & n8344));
  assign n8342 = n1686 & (n5019 | (~x7 & n4894 & ~n877));
  assign n8343 = ~n2129 & (n3573 | (~x7 & n2315 & ~n7604));
  assign n8344 = (~n550 | ~n866) & (~n661 | (~n548 & ~n1725));
  assign n8345 = n570 & ((n3436 & n4422) | (n8346 & ~n6628));
  assign n8346 = ~x7 & x0 & x6;
  assign z498 = n8355 | (x3 ? ~n8359 : ~n8348);
  assign n8348 = n8351 & ~n8353 & ~n8354 & (x0 | n8349);
  assign n8349 = (~n1080 | n8350) & (~n1300 | ~n570 | n7604);
  assign n8350 = x1 ? ((x5 | x6) & (x4 | ~x5 | ~x6)) : (~x4 | x6);
  assign n8351 = (n714 | n8352) & (~n560 | (~n704 & ~n1621));
  assign n8352 = (x0 | ~x1 | ~x2 | ~x6 | ~x7) & (~x0 | ((x1 | x6 | x7) & (~x1 | x2 | ~x6 | ~x7)));
  assign n8353 = ~n1134 & ((n543 & n3431) | (x0 & ~n3703));
  assign n8354 = n1380 & ((~x1 & ~x4 & (x2 ^ x6)) | (x4 & x6 & x1 & ~x2));
  assign n8355 = ~n643 & (n8357 | n8358 | (~x1 & ~n8356));
  assign n8356 = x2 ? ((~x0 | ~x4 | x5) & (x4 | ~x5 | x0 | ~x3)) : ((x0 & ~x3) | (~x4 ^ ~x5));
  assign n8357 = ~n1998 & ((~x1 & ~x3 & x4 & ~x5) | (x1 & ~x4 & (x3 ^ x5)));
  assign n8358 = n543 & ((~x2 & ~x3 & ~x5) | (x3 & x5 & ~n1685));
  assign n8359 = n8364 & ~n8363 & ~n8362 & ~n5542 & ~n8360;
  assign n8360 = ~n1198 & ~n8361;
  assign n8361 = (~x0 | x1 | ~x2 | x4 | ~x7) & (x0 | ~x4 | x7 | (x1 ^ ~x2));
  assign n8362 = n1145 & ((n1857 & n995) | (~x0 & ~n3929));
  assign n8363 = n1300 & n566 & (x1 ? (x2 ^ ~x5) : (~x2 ^ ~x5));
  assign n8364 = (~n560 | ~n577) & (~n904 | ~n566 | n3802);
  assign z499 = n8366 | ~n8369 | ~n8373 | (n543 & ~n8368);
  assign n8366 = ~x3 & (n8367 | (n560 & n931));
  assign n8367 = ~x4 & ((n560 & n658) | (n992 & ~n1957));
  assign n8368 = (x3 | x4 | ~x5 | x6 | x7) & (~x4 | ((x3 | (x5 ? (x6 | ~x7) : (~x6 | x7))) & (~x6 | ~x7 | ~x3 | ~x5)));
  assign n8369 = ~n5710 & n8370 & (x7 | ~n1310 | n1820);
  assign n8370 = (n1008 | n8371) & (n8372 | (x1 & x2));
  assign n8371 = (x0 | ~x1 | ~x3 | ~x4) & (~x0 | x3 | x4 | (x1 ^ ~x2));
  assign n8372 = (~x0 | ((x3 | ~x4 | ~x5 | ~x7) & (~x3 | x4 | x5 | x7))) & (x0 | x3 | x4 | ~x5 | ~x7);
  assign n8373 = ~n8374 & (x1 | n8376);
  assign n8374 = ~n643 & (x3 ? (n2332 & n543) : ~n8375);
  assign n8375 = (x0 | x1 | ~x4 | ~x5) & (x5 | (x0 ? (~x4 | (x1 ^ ~x2)) : (x4 | (x1 & x2))));
  assign n8376 = x0 ? (~x3 | (~n5257 & ~n4050)) : n8377;
  assign n8377 = x3 ? ((x4 | ~x5 | ~x6 | x7) & (~x4 | x5 | x6 | ~x7) & ((~x6 ^ ~x7) | (~x4 ^ ~x5))) : ((~x4 | x5 | ~x6 | ~x7) & (x4 | ~x5 | x6 | x7));
  assign z500 = n8379 | n8384 | ~n8389 | (n743 & ~n8388);
  assign n8379 = ~x4 & (~n8382 | (~x0 & (n8380 | ~n8381)));
  assign n8380 = n632 & ((n569 & n1301) | (~x3 & ~n1116));
  assign n8381 = (~x1 | ~x2 | ~x5 | ~x6 | x7) & (x1 | (x5 ? (x6 | ~x7) : (~x6 | x7)));
  assign n8382 = x6 ? (x7 ? n8383 : (~n3151 | ~n560)) : (x7 | n8383);
  assign n8383 = (~x0 | x2 | x3 | (~x1 ^ ~x5)) & ((~x2 & ~x3) | (x0 ? (x1 | ~x5) : (~x1 | x5)));
  assign n8384 = x4 & (~n8386 | (~n643 & ~n8385));
  assign n8385 = (~x1 | ((x0 | x5) & (x3 | ~x5 | ~x0 | x2))) & (~x0 | x1 | ((x2 | x3 | x5) & (~x5 | (~x2 & ~x3))));
  assign n8386 = ~n8387 & (~n569 | ~n3151 | ~n560);
  assign n8387 = ~x0 & ((x6 & x7 & x1 & x5) | (~x1 & (x5 ? (~x6 & ~x7) : (x6 & x7))));
  assign n8388 = (~x1 | x3 | ~x4 | x5 | ~x6) & (x1 | ((x3 | ~x4 | ~x5 | x6) & (~x3 | x5 | (~x4 ^ ~x6))));
  assign n8389 = x6 ? (~n772 | n8390) : n8391;
  assign n8390 = x0 ? (~x2 | x5) : ~x5;
  assign n8391 = (x0 | ~x1 | ~x4 | ~x5) & (x5 | (x0 ? (x4 | (x1 ^ ~x2)) : (x1 | ~x4)));
  assign z501 = n8394 | n8396 | ~n8397 | (x7 & ~n8393);
  assign n8393 = x5 ? ((~x6 | n2877) & (x0 | x1 | x6)) : (x6 | n2877);
  assign n8394 = ~x2 & ((n1234 & n2209) | (n3151 & ~n8395));
  assign n8395 = x0 ? (x1 | (~x4 ^ ~x7)) : (~x1 | (~x4 ^ x7));
  assign n8396 = n6270 & ((n828 & n632) | (~x1 & ~n2861));
  assign n8397 = n8399 & (n1008 | (~n8398 & (~n560 | ~n1331)));
  assign n8398 = n1686 & (~x1 | (~x2 & n828));
  assign n8399 = (~x2 & ~x3) ? (n765 | ~n922) : n8400;
  assign n8400 = (x0 | ~x1 | ~x5 | x7) & (~x0 | x1 | (~x5 ^ ~x7));
  assign z138 = n611 | ~n614 | (x1 ? ~n602 : ~n590);
  assign z215 = n638 | ~n648 | n3163 | (~x3 & ~n3162);
  assign z254 = n1273 | n1277 | ~n1279 | (~x0 & ~n1276);
  assign z339 = ~n1245 | (~x2 & (n1242 | (n661 & n1241)));
  assign z340 = z033;
  assign z363 = n2495 | n2503 | ~n2506 | (~n1008 & ~n2498);
  assign z364 = n2517 | ~n2524 | ~n2532 | (~n643 & ~n2521);
  assign z420 = z033;
  assign z421 = z034;
  assign z422 = z034;
  assign z423 = z034;
  assign z424 = z034;
  assign z425 = z034;
  assign z426 = z034;
  assign z427 = z034;
  assign z428 = z034;
  assign z502 = z419;
  assign z503 = z033;
  assign z504 = z034;
  assign z505 = z034;
  assign z506 = z034;
  assign z507 = z034;
  assign z508 = z034;
  assign z509 = z034;
  assign z510 = z034;
  assign z511 = z034;
  assign z512 = z034;
endmodule


