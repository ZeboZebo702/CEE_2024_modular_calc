// Benchmark "mult_3x3_64_out" written by ABC on Fri May 27 23:37:13 2022

module mult_3x3_64 ( 
    a1, a2, a3, b1, b2, b3,
    r1,r2,r3,r4,r5,r6,r7,r8  );
  input  a1, a2, a3, b1, b2, b3;
  output r1,r2,r3,r4,r5,r6,r7,r8;
  assign r1 = (~a1 | ~b1 | ((~a2 | ~a3) & (~b2 | ~b3))) & (a1 | ((a2 | b2) & (~a2 | ~a3 | b1 | ~b2 | ~b3) & (a3 | b3))) & (a2 | (a3 & (b1 | b2))) & (b3 | (b2 & (a3 | b1)));
  assign r2 = (a3 & ((b3 & ((~a1 & (~b1 | ~b2)) | (~b1 & ~b2) | (~a2 & b2))) | (a1 & b1 & ~b2 & ~b3))) | (a1 & b1 & (b2 ? ~a2 : (a2 | (~a3 & b3))));
  assign r3 = (b1 & ((a2 & ((~a1 & (b2 ? ~b3 : a3)) | (~a3 & b3 & (a1 | b2)) | (a3 & ~b3))) | (a1 & ~b3 & ((a3 & b2) | (~a2 & ~a3 & ~b2))))) | (a1 & b2 & ((~a3 & b3) | (~b1 & (a2 ^ b3))));
  assign r4 = (b2 & ((a2 & ((~a1 & a3 & (b1 ^ b3)) | (~b1 & b3 & a1 & ~a3))) | (a1 & ~a2 & ~b3 & (~a3 | ~b1)))) | (b1 & ~b2 & (a1 ? ((~a3 & ~b3) | (~a2 & a3 & b3)) : (a2 & ~a3)));
  assign r5 = (~a1 | ~b1 | ((~a2 | (~b2 & (~a3 | ~b3))) & (~a3 | ~b2 | ~b3))) & (a1 | ((b1 | b2) & (a2 | (a3 & b1)))) & (b1 | b2 | b3);
  assign r6 = (~a3 & ((a2 & b2) | (a1 & ~a2 & b1 & ~b2 & ~b3))) | (b3 & ((a1 & ~b1 & (~a2 | ~b2)) | (a3 & b1 & (a2 ^ b2)))) | (~a1 & ((a2 & (b1 ^ b2)) | (a3 & b1 & (~b2 | ~b3)))) | (b2 & ~b3 & (a2 | (a1 & ~b1)));
  assign r7 = (a2 & ((~a1 & ((~b1 & b2) | (~a3 & b1 & ~b2))) | (a3 & b2 & b3) | (~b2 & ~b3 & ~a3 & b1))) | (a1 & ((~a2 & ((~b2 & b3) | (~b1 & b2 & ~b3))) | (~b2 & b3 & (a3 | ~b1)) | (b2 & ~b3 & ~a3 & b1))) | (a3 & b1 & ((b2 & b3) | (~a2 & (~a1 | ~b2))));
  assign r8 = (~b3 | (a1 ? ((~a2 | a3 | b1 | ~b2) & (~b1 | b2 | a2 | ~a3)) : (~a3 | b1))) & ((a2 & b2) | ((a3 | (a1 & b3)) & (b1 | b3))) & (a1 | ~a2 | ~a3 | ~b1 | ~b2 | b3);
endmodule


