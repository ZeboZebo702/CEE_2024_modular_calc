// Benchmark "mult_3_64" written by ABC on Fri Dec 09 22:21:04 2022

module mult_3_64 ( 
    x0, x1, x2,
    z0, z1, z2, z3, z4, z5, z6, z7, z8  );
  input  x0, x1, x2;
  output z0, z1, z2, z3, z4, z5, z6, z7, z8;
  assign z3 = 1'b0;
  assign z0 = x0;
  assign z1 = x1;
  assign z2 = x2;
  assign z4 = 1'b0;
  assign z5 = 1'b0;
  assign z6 = 1'b0;
  assign z7 = 1'b0;
  assign z8 = 1'b0;
endmodule


