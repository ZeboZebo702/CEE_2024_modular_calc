// Benchmark "64_64_mod" written by ABC on Thu Dec 01 02:01:36 2022

module const_64_64_mod ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z000, z001, z002, z003, z004, z005, z006, z007, z008, z009, z010, z011,
    z012, z013, z014, z015, z016, z017, z018, z019, z020, z021, z022, z023,
    z024, z025, z026, z027, z028, z029, z030, z031, z032, z033, z034, z035,
    z036, z037, z038, z039, z040, z041, z042, z043, z044, z045, z046, z047,
    z048, z049, z050, z051, z052, z053, z054, z055, z056, z057, z058, z059,
    z060, z061, z062, z063, z064, z065, z066, z067, z068, z069, z070, z071,
    z072, z073, z074, z075, z076, z077, z078, z079, z080, z081, z082, z083,
    z084, z085, z086, z087, z088, z089, z090, z091, z092, z093, z094, z095,
    z096, z097, z098, z099, z100, z101, z102, z103, z104, z105, z106, z107,
    z108, z109, z110, z111, z112, z113, z114, z115, z116, z117, z118, z119,
    z120, z121, z122, z123, z124, z125, z126, z127, z128  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z000, z001, z002, z003, z004, z005, z006, z007, z008, z009, z010,
    z011, z012, z013, z014, z015, z016, z017, z018, z019, z020, z021, z022,
    z023, z024, z025, z026, z027, z028, z029, z030, z031, z032, z033, z034,
    z035, z036, z037, z038, z039, z040, z041, z042, z043, z044, z045, z046,
    z047, z048, z049, z050, z051, z052, z053, z054, z055, z056, z057, z058,
    z059, z060, z061, z062, z063, z064, z065, z066, z067, z068, z069, z070,
    z071, z072, z073, z074, z075, z076, z077, z078, z079, z080, z081, z082,
    z083, z084, z085, z086, z087, z088, z089, z090, z091, z092, z093, z094,
    z095, z096, z097, z098, z099, z100, z101, z102, z103, z104, z105, z106,
    z107, z108, z109, z110, z111, z112, z113, z114, z115, z116, z117, z118,
    z119, z120, z121, z122, z123, z124, z125, z126, z127, z128;
  wire n139, n140, n141, n143, n144, n145, n146, n147, n148, n149, n150,
    n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n163,
    n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n233, n234, n235, n236, n237, n238,
    n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257, n258, n260, n261, n262, n263,
    n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
    n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
    n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
    n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n312, n313,
    n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
    n351, n352, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
    n376, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
    n401, n402, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n422, n423, n424, n425, n426,
    n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n444, n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
    n464, n465, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n487, n488, n489,
    n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
    n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
    n515, n516, n517, n518, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
    n553, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n597, n598, n599, n600, n601, n602, n603,
    n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n616,
    n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
    n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n647, n648, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n666, n667,
    n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n685, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
    n730, n731, n732, n733, n734, n735, n736, n737, n738, n740, n741, n742,
    n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
    n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
    n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n779, n780,
    n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n798, n799, n800, n801, n802, n803, n804, n805,
    n806, n807, n808, n809, n811, n812, n813, n814, n815, n816, n817, n818,
    n819, n820, n821, n822, n824, n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838, n839, n841, n842, n843, n844,
    n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
    n857, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n878, n879, n880, n881, n882,
    n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n900, n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n913, n914, n915, n916, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
    n933, n934, n935, n937, n938, n939, n940, n941, n942, n943, n944, n945,
    n946, n947, n948, n949, n950, n951, n952, n953, n954, n956, n957, n958,
    n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
    n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
    n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
    n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1006, n1007,
    n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
    n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
    n1103, n1104, n1105, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1186, n1187, n1188,
    n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
    n1199, n1200, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1227, n1228, n1229, n1230, n1231,
    n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1240, n1241, n1242,
    n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1253,
    n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1275,
    n1276, n1277, n1278, n1279, n1281, n1282, n1283, n1284, n1285, n1286,
    n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1320,
    n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1332, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
    n1363, n1364, n1365, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1384,
    n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
    n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1416, n1417,
    n1418, n1419, n1420, n1421, n1422, n1424, n1425, n1426, n1427, n1428,
    n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
    n1472, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
    n1483, n1484, n1485, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
    n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1503, n1504,
    n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
    n1515, n1516, n1517, n1518, n1519, n1520, n1522, n1523, n1524, n1525,
    n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
    n1536, n1537, n1538, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
    n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1562, n1563, n1564, n1565, n1566, n1567,
    n1568, n1569, n1570, n1571, n1573, n1574, n1575, n1576, n1577, n1578,
    n1579, n1580, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
    n1590, n1591, n1592, n1593, n1594, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
    n1622, n1623, n1624, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
    n1633, n1634, n1635, n1636, n1637, n1638, n1640, n1641, n1642, n1643,
    n1644, n1645, n1646, n1647, n1648, n1650, n1651, n1652, n1653, n1654,
    n1655, n1656, n1657, n1658, n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1671, n1672, n1673, n1674, n1675, n1676,
    n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1699,
    n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
    n1710, n1711, n1712, n1713, n1714, n1715, n1717, n1718, n1719, n1720,
    n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1736, n1737, n1738, n1739, n1740, n1741,
    n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1750, n1751, n1752,
    n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
    n1763, n1764, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1800, n1801, n1802, n1803, n1804, n1805,
    n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
    n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
    n1827, n1828, n1829, n1830, n1831, n1832, n1834, n1835, n1836, n1837,
    n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
    n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
    n1892, n1893, n1894, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
    n1903, n1904, n1905, n1906, n1908, n1909, n1910, n1911, n1912, n1913,
    n1914, n1915, n1916, n1917, n1919, n1920, n1921, n1922, n1923, n1924,
    n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
    n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
    n1946, n1947, n1948, n1949, n1950, n1952, n1953, n1954, n1955, n1956,
    n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
    n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
    n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
    n2011, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
    n2022, n2023, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
    n2033, n2035, n2036, n2037, n2038, n2039, n2040, n2041;
  assign z121 = 1'b0;
  assign z000 = n139 & n140 & n141;
  assign n139 = ~x6 & ~x4 & x5 & ~x7;
  assign n140 = ~x0 & ~x1;
  assign n141 = x2 & x3;
  assign z001 = ~n149 | (~x1 & (~n143 | ~n148));
  assign n143 = (x3 | (~n145 & (~x0 | n144))) & (x0 | ~x3 | n147);
  assign n144 = (~x2 | x4 | ~x5 | x6 | x7) & (x2 | ~x4 | x5 | ~x6 | ~x7);
  assign n145 = n146 & ((~x2 & ~x6 & (x4 ^ x7)) | (x2 & ~x4 & x6 & x7));
  assign n146 = ~x0 & ~x5;
  assign n147 = (~x2 | ~x5 | x6 | (x4 ^ ~x7)) & (x2 | ~x4 | x5 | ~x6 | x7);
  assign n148 = x5 ? (x0 ? (x2 | ~x4) : (x4 | (x2 & x3))) : (x0 ? (x4 | (~x2 ^ x3)) : (~x2 | ~x4));
  assign n149 = ~n150 & n156 & (~x4 | n154 | ~n155);
  assign n150 = ~x0 & (x6 ? ~n152 : (n151 & ~n153));
  assign n151 = ~x2 & x4;
  assign n152 = x1 ? ((x2 | x3 | x4 | ~x5) & (~x2 | ~x3 | ~x4 | x5)) : (x4 | (x2 ? (~x3 | ~x5) : x5));
  assign n153 = x1 ? (x3 | ~x5) : (~x3 | x5);
  assign n154 = x2 ? (x3 & ~x5) : (~x3 & x5);
  assign n155 = ~x0 & x1;
  assign n156 = (n160 | ~n161) & (~n157 | ~n158 | ~n159);
  assign n157 = ~x2 & x0 & ~x1;
  assign n158 = ~x3 & ~x4;
  assign n159 = ~x5 & ~x6;
  assign n160 = (~x2 | x5 | x6 | x7) & (x2 | ~x5 | ~x6 | ~x7);
  assign n161 = ~x4 & x3 & ~x0 & x1;
  assign z002 = ~n172 | (~x1 & (x6 ? ~n163 : ~n167));
  assign n163 = (x7 | n165) & (x4 | ~x7 | ~n164 | n166);
  assign n164 = x2 & ~x3;
  assign n165 = (x4 | ((~x0 | x3 | (~x2 ^ ~x5)) & (x0 | x2 | ~x3 | x5))) & (x0 | x2 | ~x3 | ~x4 | ~x5);
  assign n166 = x0 ^ x5;
  assign n167 = (n168 | ~n169) & (~n170 | ~n171);
  assign n168 = (~x2 | ~x3 | x5 | x7) & (x2 | x3 | ~x5 | ~x7);
  assign n169 = ~x0 & x4;
  assign n170 = x0 & x2 & ~x3;
  assign n171 = x7 & ~x4 & x5;
  assign n172 = ~n177 & (~n155 | (n173 & n180));
  assign n173 = (~x7 | n175) & (~x2 | ~n174 | ~n176);
  assign n174 = ~x7 & x5 & ~x6;
  assign n175 = (~x3 | ((~x2 | x6 | (x4 ^ x5)) & (~x5 | ~x6 | x2 | x4))) & (x2 | x3 | ~x4 | x5 | x6);
  assign n176 = ~x3 & x4;
  assign n177 = ~x1 & (x3 ? ~n179 : ~n178);
  assign n178 = x2 ? ((x0 | ~x5) & (~x0 | x5 | x6 | x7)) : (x5 ? ((x6 | x7) & (~x0 | (x6 & x7))) : ((~x6 | ~x7) & (x0 | (~x6 & ~x7))));
  assign n179 = (x0 | ((~x5 | (x6 ? ~x2 : ~x7)) & (~x6 | ~x7 | x2 | x5))) & (x2 | ~x5 | (~x0 & x6));
  assign n180 = (x2 | (x3 ? (x5 | x6) : (~x5 | ~x6))) & (x7 | (x3 ? ((x5 | ~x6) & (~x2 | ~x5 | x6)) : (x5 | x6))) & (~x2 | x5 | (x3 & ~x6));
  assign z003 = ~n194 | ~n190 | n182 | n186;
  assign n182 = ~n183 & ((n155 & ~n185) | (~x1 & ~n184));
  assign n183 = ~x6 ^ x7;
  assign n184 = x3 ? ((x0 | ~x2 | (~x4 & ~x5)) & (~x0 | x2 | ~x4 | ~x5)) : ((x4 & x5) | (x0 ^ x2));
  assign n185 = (~x2 | (~x3 ^ x4)) & (x2 | x3 | x4 | x5);
  assign n186 = ~x2 & ((n169 & ~n189) | (~n187 & ~n188));
  assign n187 = (x3 | x4 | ~x6 | x7) & (~x3 | ~x4 | x6 | ~x7);
  assign n188 = x0 ? (x1 | x5) : (~x1 | ~x5);
  assign n189 = (x1 | ~x5 | (x3 ? (x6 | x7) : ~x6)) & (~x1 | ~x3 | x5 | ~x6 | ~x7);
  assign n190 = (x2 | n192) & (x3 | ~n191 | ~n193);
  assign n191 = ~x6 & ~x7;
  assign n192 = (x0 | x1 | ~x3 | ~x6 | ~x7) & ((~x0 ^ x1) | (x3 ? (x6 | x7) : (~x6 | ~x7)));
  assign n193 = x2 & ~x0 & ~x1;
  assign n194 = ~n202 & (n195 | ~n196) & (x2 | n197);
  assign n195 = (~x1 | x3 | ~x4 | x6 | x7) & (x1 | x4 | (x3 ? x6 : (~x6 | ~x7)));
  assign n196 = ~x5 & ~x0 & x2;
  assign n197 = (n198 | n199) & (x0 | ~n200 | ~n201);
  assign n198 = x3 ? (x4 | ~x7) : (~x4 | x7);
  assign n199 = x0 ? (x1 | x6) : (~x1 | ~x6);
  assign n200 = ~x7 & ~x4 & x6;
  assign n201 = ~x1 & x3;
  assign n202 = n203 & ((x1 & ~n204) | (n205 & n206));
  assign n203 = ~x0 & x2;
  assign n204 = x3 ? (~x4 | ~x6) : (x4 | x6);
  assign n205 = ~x1 & ~x3;
  assign n206 = x7 & x4 & ~x6;
  assign z004 = ~n222 | (~x0 & (~n208 | n214 | ~n218));
  assign n208 = x3 ? (~n209 | ~n213) : n210;
  assign n209 = ~x1 & ~x2;
  assign n210 = (~x5 | n211) & (~x1 | x5 | x6 | n212);
  assign n211 = (x1 | ((~x2 | x4 | x6 | ~x7) & (~x6 | x7 | x2 | ~x4))) & (~x1 | x2 | ~x4 | ~x6 | ~x7);
  assign n212 = x2 ? (~x4 | x7) : (x4 | ~x7);
  assign n213 = x4 & ~x5 & (~x6 ^ x7);
  assign n214 = n215 & (n217 | (x3 & ~n216));
  assign n215 = x1 & ~x2;
  assign n216 = x4 ? (~x5 | x7) : (x5 | ~x7);
  assign n217 = ~x7 & x5 & ~x3 & x4;
  assign n218 = (n219 | n220) & (~x2 | n221);
  assign n219 = x3 ? (~x5 | x7) : (x5 | ~x7);
  assign n220 = x1 ? (~x2 | ~x4) : (x2 | x4);
  assign n221 = (x3 | ((x1 | (x4 ? x7 : (x5 | ~x7))) & (~x1 | x4 | ~x5 | x7))) & (~x1 | ~x3 | (x4 ? (x5 | x7) : ~x7));
  assign n222 = n227 & (n223 | n224) & (n225 | ~n226);
  assign n223 = ~x4 ^ x5;
  assign n224 = (x1 | ((~x0 | ((x2 | ~x3 | x7) & (x3 | ~x7))) & (~x7 | ((x2 | x3) & (x0 | ~x2 | ~x3))))) & (x0 | ~x1 | x2 | (~x3 ^ ~x7));
  assign n225 = (x3 | x4 | ~x5 | x6 | x7) & (~x3 | ((~x4 | ~x5 | (~x6 ^ ~x7)) & (~x6 | x7 | x4 | x5)));
  assign n226 = ~x2 & x0 & ~x1;
  assign n227 = (n229 | n230) & (~n158 | ~n228 | ~n231);
  assign n228 = ~x5 & x7;
  assign n229 = x4 ? (~x5 | ~x7) : (x5 | x7);
  assign n230 = (~x0 | x1 | x2 | x3) & (x0 | (x1 ? (~x2 | x3) : ~x3));
  assign n231 = x2 & x0 & ~x1;
  assign z005 = n233 | ~n246 | ~n255 | (~n244 & ~n245);
  assign n233 = ~x1 & (n234 | n239 | (n170 & n243));
  assign n234 = ~x2 & ((~n236 & n237) | (n235 & n238));
  assign n235 = x5 & ~x6 & (x4 ^ x7);
  assign n236 = (~x3 | x4 | x6 | x7) & (x3 | ~x4 | ~x6 | ~x7);
  assign n237 = x0 & ~x5;
  assign n238 = ~x0 & ~x3;
  assign n239 = ~n241 & (x0 ? n242 : n240);
  assign n240 = x2 & x6;
  assign n241 = (x3 | x4 | ~x5 | x7) & (~x3 | ~x4 | x5 | ~x7);
  assign n242 = ~x2 & ~x6;
  assign n243 = ~x7 & x4 & x5 & ~x6;
  assign n244 = ~x5 ^ x6;
  assign n245 = (x0 | (x1 ? (x2 ? (~x3 | x4) : (x3 | ~x4)) : (x4 | (~x2 ^ x3)))) & (~x0 | x1 | x2 | ~x3 | ~x4);
  assign n246 = ~n248 & ~n253 & (~n158 | ~n247 | ~n231);
  assign n247 = x5 & x6;
  assign n248 = n155 & ((~n250 & ~n251) | (n249 & n252));
  assign n249 = x4 & ~x2 & ~x3;
  assign n250 = x3 ? (~x5 | ~x7) : (x5 | x7);
  assign n251 = x2 ? (~x4 | x6) : (x4 | ~x6);
  assign n252 = x5 & x6 & ~x7;
  assign n253 = n254 & (x2 ? (x4 & ~x5) : (~x4 ^ x5));
  assign n254 = ~x3 & x0 & ~x1;
  assign n255 = x0 | (n256 & (x2 ? n258 : n257));
  assign n256 = x1 ? ((~x2 | x3 | x4 | ~x5) & (~x4 | x5 | x2 | ~x3)) : ((~x2 | ~x3 | (~x4 ^ ~x5)) & (~x4 | x5 | x2 | x3));
  assign n257 = (x1 | ((x4 | ~x5 | ~x6) & (~x3 | ~x4 | x5 | x6))) & (~x1 | x3 | x5 | x6);
  assign n258 = (x1 | x3 | ~x4 | ~x5 | ~x6) & (~x1 | ~x3 | ((~x5 | ~x6) & (x4 | x5 | x6)));
  assign z006 = n267 | n270 | (~x0 & ~n260) | ~n277;
  assign n260 = x5 ? n261 : (~n265 & (x2 | n264));
  assign n261 = (x7 | n262) & (x4 | ~x6 | ~x7 | ~n263);
  assign n262 = (x3 | ((~x1 | x2 | ~x4 | ~x6) & (x1 | (x2 ? (x4 | ~x6) : x6)))) & (~x1 | ~x3 | (x2 ? (~x4 | x6) : (x4 | ~x6)));
  assign n263 = x3 & ~x1 & x2;
  assign n264 = (~x7 | (~x3 ^ x4) | (~x1 ^ ~x6)) & (~x1 | x3 | x4 | ~x6 | x7);
  assign n265 = n164 & n266 & ~x1 & ~x4;
  assign n266 = x6 & x7;
  assign n267 = n268 & (x2 ? (n174 & n176) : ~n269);
  assign n268 = x0 & ~x1;
  assign n269 = (x3 | x4 | ~x5 | x6 | x7) & (x5 | ((x3 | ((x6 | ~x7) & (~x4 | ~x6 | x7))) & (~x3 | ~x4 | x6 | x7)));
  assign n270 = ~x3 & (~n272 | (~x5 & ~n271));
  assign n271 = (x0 | (x1 ? (x4 | x6) : (x2 | ~x6))) & (x1 | ~x2 | ~x6 | (~x0 & ~x4));
  assign n272 = (~n274 | ~n276) & (n273 | n275);
  assign n273 = x4 ^ x5;
  assign n274 = ~x1 & x2;
  assign n275 = (x0 | ~x2 | (x1 ^ x6)) & (~x0 | x1 | x2 | ~x6);
  assign n276 = ~x6 & ~x4 & x5;
  assign n277 = ~n278 & (n283 | n284) & (n281 | n282);
  assign n278 = n279 & ~n280;
  assign n279 = ~x0 & x3;
  assign n280 = (x2 | ((~x4 | x5 | x6) & (x1 | ~x5 | ~x6))) & (~x1 | (x4 ? (x5 | ~x6) : (~x5 | (~x2 & x6))));
  assign n281 = ~x4 ^ x6;
  assign n282 = (x0 | ((~x1 | x2 | x3 | ~x5) & (~x3 | x5 | x1 | ~x2))) & (~x0 | x1 | x2 | ~x3 | ~x5);
  assign n283 = x5 ^ x7;
  assign n284 = (n286 | ~n287) & (~x3 | ~n157 | ~n285);
  assign n285 = ~x4 & ~x6;
  assign n286 = x1 ? (x3 | x6) : (~x3 | ~x6);
  assign n287 = x4 & ~x0 & x2;
  assign z007 = ~n303 | (~x0 & ~n289) | (~n295 & ~n296);
  assign n289 = x5 ? (x3 ? n291 : n290) : n292;
  assign n290 = (~x4 | ((~x2 | x6 | x7) & (~x1 | (x2 ? x7 : (x6 | ~x7))))) & (~x6 | ((x2 | x4 | ~x7) & (x1 | (x2 ? (x4 | x7) : ~x7))));
  assign n291 = (~x6 | (x1 ? (x2 | ~x7) : (~x2 | x7))) & (x1 | x2 | x6 | (x4 ^ x7));
  assign n292 = (x1 | n294) & (~x1 | ~x4 | ~n266 | ~n293);
  assign n293 = ~x2 & x3;
  assign n294 = (~x4 | ((x2 | ~x7 | (~x3 ^ x6)) & (~x2 | ~x3 | ~x6 | x7))) & (~x2 | x6 | (x3 & x4) | x7);
  assign n295 = x3 ^ x5;
  assign n296 = ~n299 & (x0 ? (~n209 | ~n297) : n298);
  assign n297 = ~x7 & x4 & ~x6;
  assign n298 = (~x1 | ~x6 | (x2 ? x4 : x7)) & (x6 | ((x2 | x4 | ~x7) & (x1 | (x2 ? ~x7 : (~x4 | x7)))));
  assign n299 = ~n300 & (n302 | (n155 & n301));
  assign n300 = x6 ^ x7;
  assign n301 = x2 & x4;
  assign n302 = ~x4 & ~x2 & x0 & ~x1;
  assign n303 = ~n308 & ((~n304 & ~n305) | (~n306 & n307));
  assign n304 = ~x3 & x5;
  assign n305 = x3 & ~x5;
  assign n306 = ~x1 & ((~x2 & ((~x6 & ~x7) | (x0 & x6 & x7))) | (~x6 & x7 & ~x0 & x2));
  assign n307 = ~n155 | ((x2 | ((~x6 | x7) & (x4 | x6 | ~x7))) & (~x6 | (x7 ? ~x2 : x4)));
  assign n308 = ~n309 & n310;
  assign n309 = (~x2 | x3 | (x4 & x5 & x7)) & (~x5 | ~x7 | x2 | ~x4);
  assign n310 = ~x6 & x0 & ~x1;
  assign z008 = ~n319 | (n312 & ~n318) | (~x2 & ~n313);
  assign n312 = ~x0 & ~x4;
  assign n313 = ~n316 & (x3 | (~n315 & (~x4 | n314)));
  assign n314 = (x0 | ~x1 | x5 | ~x6 | x7) & (~x7 | ((~x0 | x1 | (~x5 ^ x6)) & (x0 | ~x1 | x5 | x6)));
  assign n315 = x5 & n312 & (x1 ? (~x6 ^ x7) : (x6 & ~x7));
  assign n316 = n317 & (x1 ? (x5 & n266) : (~x5 & ~n300));
  assign n317 = ~x4 & ~x0 & x3;
  assign n318 = (x1 | (x2 ? ((~x5 | x7) & (~x3 | x5 | ~x7)) : (~x7 | (x3 ^ x5)))) & (~x1 | x2 | x3 | x5 | x7);
  assign n319 = ~n320 & n328 & (~x4 | (~n323 & n325));
  assign n320 = n203 & ((~x3 & ~n321) | (x1 & x3 & n322));
  assign n321 = (x1 | x4 | ~x7 | (x5 ^ x6)) & (~x1 | ~x4 | ~x5 | x6 | x7);
  assign n322 = x4 & ~x5 & (x6 ^ x7);
  assign n323 = ~x3 & ~n324;
  assign n324 = (x0 | ~x1 | x2 | ~x5 | x7) & (~x0 | x1 | x5 | (x2 ^ x7));
  assign n325 = x5 ? ((~x7 | n326) & (~x3 | x7 | ~n327)) : (x7 | n326);
  assign n326 = (~x0 | x1 | x2 | ~x3) & (x0 | ~x1 | ~x2 | x3);
  assign n327 = x2 & ~x0 & x1;
  assign n328 = (x4 | n329) & (x0 | ~x4 | n330);
  assign n329 = x0 ? (x1 | (x2 ? (x3 | ~x7) : x7)) : (~x1 | (x2 ? ~x7 : (~x3 | x7)));
  assign n330 = (x2 | ~x3 | ~x7) & (x1 | (x2 ? (~x3 ^ x7) : (x3 | x7)));
  assign z009 = n342 | ~n346 | (~x1 & ~n332);
  assign n332 = (~n340 | ~n341) & (x3 | (~n333 & ~n337));
  assign n333 = n334 & (x0 ? (x4 & ~n335) : (~x4 & ~n336));
  assign n334 = x5 & ~x7;
  assign n335 = ~x2 ^ x6;
  assign n336 = x2 ^ x6;
  assign n337 = n339 & ~x0 & n338;
  assign n338 = ~x2 & ~x4;
  assign n339 = x7 & ~x5 & ~x6;
  assign n340 = x3 & ~x0 & x2;
  assign n341 = x7 & ~x6 & x4 & ~x5;
  assign n342 = ~x0 & ((x4 & ~n344) | (n343 & ~n345));
  assign n343 = ~x1 & ~x4;
  assign n344 = (~x1 | ((~x2 | ~x3 | ~x5 | ~x6) & (x5 | x6 | x2 | x3))) & (x1 | ~x2 | ~x3 | x5 | ~x6);
  assign n345 = (x2 | ~x6 | (x3 ^ x5)) & (~x2 | x3 | ~x5 | x6);
  assign n346 = n349 & (~x4 | (n347 & (~n155 | n348)));
  assign n347 = (~x0 | x1 | x3 | x5) & (x0 | ((~x1 | (x2 ? (x3 | x5) : (~x3 | ~x5))) & (~x3 | ~x5 | x1 | ~x2)));
  assign n348 = (~x2 | x3 | ~x5 | x6 | x7) & (x2 | ~x3 | x5 | ~x6 | ~x7);
  assign n349 = n350 & (~n193 | ~n351) & (~n157 | ~n352);
  assign n350 = (~x0 | x1 | x3 | x4) & (x0 | ((~x3 | ~x4 | x1 | x2) & (~x1 | x3 | x4)));
  assign n351 = ~x5 & ~x3 & ~x4;
  assign n352 = ~x6 & x5 & ~x3 & x4;
  assign z010 = n361 | ~n364 | (~x0 & ~n354) | ~n369;
  assign n354 = x2 ? (~n356 & (~x1 | n355)) : n358;
  assign n355 = (x3 | x4 | ~x5 | ~x6 | x7) & (~x3 | ~x4 | x5 | x6 | ~x7);
  assign n356 = n357 & ((n158 & n334) | (x3 & ~n229));
  assign n357 = ~x1 & x6;
  assign n358 = x4 ? n360 : (~n359 | ~n205);
  assign n359 = ~x6 & (~x5 ^ ~x7);
  assign n360 = (x1 | ~x7 | (x3 ? (~x5 | x6) : (x5 | ~x6))) & (~x1 | ~x3 | x5 | ~x6 | x7);
  assign n361 = ~x1 & (x5 ? ~n362 : (n312 & ~n363));
  assign n362 = (x0 | ((~x2 | x3 | (~x4 ^ ~x6)) & (x4 | x6 | x2 | ~x3))) & (x2 | ((~x3 | ~x4 | ~x6) & (~x0 | x3 | x4 | x6)));
  assign n363 = x2 ? (~x3 | x6) : (x3 | ~x6);
  assign n364 = (n366 | n367) & (~n365 | ~n368);
  assign n365 = ~x3 & ~x2 & x0 & ~x1;
  assign n366 = x4 ? (x6 | x7) : (~x6 | ~x7);
  assign n367 = x0 ? (x1 | ~x5 | (x2 & x3)) : ((~x2 | ~x3 | x5) & (~x1 | (~x2 & x5)));
  assign n368 = x4 & x5 & x6 & ~x7;
  assign n369 = ~n370 & ~n372 & ~n373 & (n375 | n376);
  assign n370 = ~x2 & ~n371;
  assign n371 = (x1 | (x0 ? (~x4 | x5) : (x3 ? (x4 | x5) : (~x4 | ~x5)))) & (x0 | ~x1 | x4 | ~x5);
  assign n372 = n274 & ((x0 & ~x3 & x4 & ~x5) | (~x0 & ~x4 & (~x3 ^ x5)));
  assign n373 = n155 & ((n159 & n338) | (x2 & ~n374));
  assign n374 = x4 ? (x5 | ~x6) : (~x5 | x6);
  assign n375 = x4 ? (x6 | ~x7) : (~x6 | x7);
  assign n376 = (x2 | (x0 ? (x1 | ~x5) : (~x1 | x5))) & (x0 | ~x1 | ((x3 | x5) & (~x2 | ~x3 | ~x5)));
  assign z011 = ~n395 | (~x1 & (n378 | ~n381 | ~n387));
  assign n378 = ~x0 & ((n301 & ~n380) | (~x2 & ~n379));
  assign n379 = (~x3 | ~x4 | ~x5 | x6 | x7) & (x3 | (x4 ? (~x6 | (x5 ^ x7)) : (x6 | (x5 ^ ~x7))));
  assign n380 = (x3 | x5 | ~x6 | ~x7) & (~x3 | x7 | (x5 ^ x6));
  assign n381 = (n384 | n385) & (~n382 | ~n383 | ~n386);
  assign n382 = ~x4 & ~x5;
  assign n383 = ~x6 & x7;
  assign n384 = x3 ? (x6 | ~x7) : (~x6 | x7);
  assign n385 = x0 ? (x2 | ~x4) : (~x2 | x4);
  assign n386 = ~x3 & x0 & ~x2;
  assign n387 = ~n389 & ~n390 & (x0 | n388) & n392;
  assign n388 = (x6 | (x2 ? (~x5 | (x3 ^ x4)) : (x5 | (~x3 ^ x4)))) & (x2 | x3 | x4 | x5 | ~x6);
  assign n389 = ~n374 & ((~x2 & x3) | (x0 & x2 & ~x3));
  assign n390 = ~n273 & (x3 ? (x6 & n391) : (~x6 & n203));
  assign n391 = x0 & ~x2;
  assign n392 = (~n386 | ~n393) & n394;
  assign n393 = x6 & ~x4 & ~x5;
  assign n394 = (~x0 | x2 | x3 | ~x4 | x6) & (x0 | ~x2 | ~x3 | x4 | ~x6);
  assign n395 = (n281 | n400) & (~n155 | (n396 & n399));
  assign n396 = (n223 | n397) & (~x2 | n398);
  assign n397 = (~x2 | x3 | x6 | ~x7) & (x2 | ~x3 | ~x6 | x7);
  assign n398 = (~x3 | x5 | ~x6 | (~x4 ^ ~x7)) & (x3 | ~x4 | ~x5 | x6 | x7);
  assign n399 = (x5 | (x2 ? ((x3 | ~x4 | ~x6) & (x4 | x6)) : ((~x4 | x6) & (x3 | x4 | ~x6)))) & (~x2 | ((x4 | ~x5 | ~x6) & (~x3 | ~x4 | x6))) & (x2 | ~x5 | (x4 ^ x6));
  assign n400 = (~n231 | ~n402) & (~x7 | n153 | ~n401);
  assign n401 = ~x0 & ~x2;
  assign n402 = ~x7 & ~x3 & x5;
  assign z012 = ~n412 | (~x1 & ~n404) | (~x0 & x1 & ~n410);
  assign n404 = x3 ? (n406 & (n385 | n405)) : n408;
  assign n405 = x5 ? (x6 | x7) : (~x6 | ~x7);
  assign n406 = n407 & (~n191 | ~n401 | n273);
  assign n407 = (~x0 | x2 | x4 | ~x5 | ~x7) & (x0 | ~x2 | ~x4 | x5 | x7);
  assign n408 = x0 ? (~n151 | ~n339) : n409;
  assign n409 = (~x5 | ((~x6 | (x2 ? (~x4 | ~x7) : (x4 ^ ~x7))) & (x2 | x4 | x6 | x7))) & (~x2 | x4 | x5 | (x6 ^ ~x7));
  assign n410 = (~x2 | x3 | ~x4 | ~n174) & (x4 | n411);
  assign n411 = (x2 | x3 | ~x5 | ~x6 | x7) & (~x7 | (x2 ? (x5 | (~x3 ^ x6)) : (~x5 | (x3 ^ x6))));
  assign n412 = ~n415 & (n413 | n414) & (n419 | n420);
  assign n413 = x5 ? (x6 | ~x7) : (~x6 | x7);
  assign n414 = (x2 | ((x1 | x3 | ~x4) & (x0 | ~x3 | x4))) & (~x0 | x1 | ~x2 | x3 | x4) & (x0 | (x1 ? ~x3 : (x3 | ~x4)));
  assign n415 = ~n416 & ((n155 & ~n418) | (~x1 & ~n417));
  assign n416 = ~x5 ^ x7;
  assign n417 = (x2 | ((~x3 | x4 | x6) & (~x0 | x3 | ~x6))) & (~x4 | ~x6 | x0 | ~x3) & (x3 | ((x4 | ~x6) & (~x2 | ~x4 | x6)));
  assign n418 = (~x2 | ~x4 | (~x3 ^ x6)) & (x3 | x4 | x6) & (x2 | (x3 ? (x4 | ~x6) : x6));
  assign n419 = x5 ? (~x6 | ~x7) : (x6 | x7);
  assign n420 = (x1 | ((x2 | ((~x3 | ~x4) & (~x0 | x3 | x4))) & (~x3 | x4 | x0 | ~x2))) & (x0 | ~x1 | ((x3 | ~x4) & (~x2 | (x3 & ~x4))));
  assign z013 = ~n436 | (x3 ? (n422 | n426) : ~n429);
  assign n422 = x4 & (x6 ? ~n425 : (~n423 & n424));
  assign n423 = x2 ^ x7;
  assign n424 = ~x0 & x5;
  assign n425 = (x1 | ((~x5 | x7 | x0 | ~x2) & (~x0 | x2 | x5))) & (x0 | ~x1 | ((x2 | ~x5 | ~x7) & (x5 | (~x2 & x7))));
  assign n426 = ~x4 & ((~n244 & ~n427) | (~x2 & ~n428));
  assign n427 = (~x0 | x1 | x2 | ~x7) & (x0 | ~x1 | ~x2 | x7);
  assign n428 = (~x0 | x1 | x5 | x6 | x7) & (x0 | ((~x1 | ~x5 | ~x6 | x7) & (x1 | x5 | (x6 ^ ~x7))));
  assign n429 = ~n430 & (x0 | (n433 & (~x6 | n432)));
  assign n430 = ~n416 & ~n431;
  assign n431 = (~x0 | x1 | x2 | ~x4 | ~x6) & (x0 | ~x1 | x4 | (x2 ^ ~x6));
  assign n432 = (~x7 | ((x1 | x2 | ~x4 | ~x5) & (~x1 | (x2 ? (x4 | ~x5) : (~x4 | x5))))) & (x1 | x5 | x7 | (~x2 ^ x4));
  assign n433 = (x5 | ~x6 | n434) & (x6 | ((~x5 | n434) & (n283 | ~n435)));
  assign n434 = (x1 | (x2 ? ~x7 : (x4 | x7))) & (~x1 | ~x2 | ~x4 | x7);
  assign n435 = ~x4 & x1 & ~x2;
  assign n436 = ~n438 & (n437 | n441) & (~n268 | n442);
  assign n437 = x4 ? (x5 | x6) : (~x5 | ~x6);
  assign n438 = ~x0 & (x2 ? ~n440 : ~n439);
  assign n439 = (~x5 | x7 | x3 | ~x4) & (~x3 | ((x1 | ((~x4 | x5 | x7) & (~x5 | ~x7))) & (~x1 | x4 | x5 | ~x7)));
  assign n440 = (~x1 | x3 | ~x4 | ~x5 | ~x7) & (x1 | x5 | (x3 ? (x4 ^ x7) : (~x4 | x7)));
  assign n441 = (x7 | ((x0 | ~x1 | ~x2 | x3) & (x1 | (x0 ? (~x2 ^ x3) : (~x2 | ~x3))))) & (x0 | ~x7 | (x3 ? ~x1 : x2));
  assign n442 = (x2 | ((~x3 | ~x4 | ~x5 | x7) & (x3 | ((x5 | x7) & (x4 | ~x5 | ~x7))))) & (~x2 | x3 | x5 | ~x7);
  assign z014 = n450 | ~n452 | (~x1 & ~n444);
  assign n444 = (~x7 | ~n445 | n446) & (x3 | n447);
  assign n445 = ~x5 & x3 & ~x0 & ~x2;
  assign n446 = x4 ^ x6;
  assign n447 = (x7 | n449) & (x0 | ~n448 | ~n338);
  assign n448 = x7 & ~x5 & x6;
  assign n449 = (x0 | ((~x2 | x4 | (~x5 ^ ~x6)) & (~x5 | ~x6 | x2 | ~x4))) & (~x5 | x6 | ~x0 | ~x4);
  assign n450 = x2 & (x0 ? (n205 & n393) : ~n451);
  assign n451 = x3 ? ((x6 | (x1 ? (~x4 ^ x5) : (~x4 | ~x5))) & (x5 | ~x6 | x1 | x4)) : ((x5 | ~x6 | ~x1 | ~x4) & (~x5 | x6 | x1 | x4));
  assign n452 = ~n453 & ~n459 & ~n463 & (~n155 | n456);
  assign n453 = ~x2 & (n455 | (~x1 & ~n454));
  assign n454 = (~x4 | ((x0 | x3 | x6) & (~x0 | ~x3 | ~x5 | ~x6))) & (x0 | (x3 ? (x4 | ~x6) : (~x5 | x6))) & (~x0 | (x3 ? (x4 | x6) : (~x6 | (x4 & x5))));
  assign n455 = ~x0 & x1 & (x3 ? (x4 & ~x6) : (x4 ^ ~x6));
  assign n456 = (~x2 | ~x3 | ~x4 | ~n457) & (x2 | x4 | n458);
  assign n457 = ~x7 & ~x5 & x6;
  assign n458 = (x3 | ~x5 | ~x6 | x7) & (~x3 | (x5 ? (x6 | x7) : (~x6 | ~x7)));
  assign n459 = ~n300 & ((n460 & n462) | (x2 & ~n461));
  assign n460 = x3 & x4 & x5;
  assign n461 = (x1 | (x0 ^ ~x3) | (x4 ^ ~x5)) & (x0 | ~x1 | (x3 ? (x4 | x5) : (~x4 | ~x5)));
  assign n462 = ~x2 & ~x0 & ~x1;
  assign n463 = ~n183 & ((n155 & n464) | (x4 & ~n465));
  assign n464 = ~x4 & x2 & ~x3;
  assign n465 = (~x0 | x1 | x2 | ~x3 | x5) & (x0 | ~x2 | (x1 ? (~x3 | ~x5) : x3));
  assign z015 = n474 | n479 | (x2 ? ~n481 : ~n467);
  assign n467 = x6 ? n470 : (~n469 & (x1 | n468));
  assign n468 = (x5 | (~x0 ^ x3) | (x4 ^ x7)) & (~x0 | ~x5 | (x3 ? (x4 | ~x7) : (~x4 | x7)));
  assign n469 = n155 & ((~x3 & x4 & ~x5 & ~x7) | (x7 & (x3 ? (~x4 ^ x5) : (~x4 & x5))));
  assign n470 = (~n471 | ~n472) & (x0 | n473);
  assign n471 = x4 & x5 & x7;
  assign n472 = ~x3 & x0 & ~x1;
  assign n473 = (x7 | ((x1 | x3 | x4 | x5) & ((~x3 ^ x5) | (x1 ^ ~x4)))) & (~x3 | x4 | ~x7 | (~x1 ^ ~x5));
  assign n474 = ~x1 & (n476 | n478 | (~x2 & ~n475));
  assign n475 = (~x7 | (x0 ? ((x4 | x5) & (~x3 | ~x4 | ~x5)) : (x3 | (~x4 ^ x5)))) & (~x3 | ~x4 | x7 | (~x0 ^ x5));
  assign n476 = ~n477 & (x0 ^ x3);
  assign n477 = (~x2 | ~x4 | x5 | x7) & (x4 | (x2 ? (~x5 ^ x7) : (~x5 | ~x7)));
  assign n478 = n203 & ((x3 & x4 & x5 & x7) | (~x3 & ~x7 & (x4 | ~x5)));
  assign n479 = n155 & ~n480;
  assign n480 = (~x5 | ((~x3 | x4 | (~x2 ^ ~x7)) & (~x2 | x7 | (x3 & ~x4)))) & (~x2 | x4 | x5 | x7) & (x2 | ~x7 | ((~x4 | x5) & (x3 | (~x4 & x5))));
  assign n481 = x0 ? (~n205 | ~n243) : (~n482 & n484);
  assign n482 = ~n483 & x1 & ~x6;
  assign n483 = (~x3 | x4 | ~x5 | x7) & (x3 | ~x4 | x5 | ~x7);
  assign n484 = (n183 | n485) & (x1 | ~n448 | ~n158);
  assign n485 = (~x1 | ~x3 | ~x4 | x5) & (x1 | x3 | x4 | ~x5);
  assign z016 = n487 | n490 | ~n496 | (~x1 & ~n495);
  assign n487 = ~x0 & (x1 ? ~n489 : ~n488);
  assign n488 = (x3 | ((~x5 | ~x6 | x2 | ~x4) & (~x2 | (x4 ? (x5 | x6) : (~x5 | ~x6))))) & (x2 | ~x3 | ~x4 | (x5 ^ ~x6));
  assign n489 = (~x2 | ~x3 | x4 | ~x5 | ~x6) & (x2 | ((~x5 | x6 | x3 | ~x4) & (x5 | (x3 ? (x4 ^ ~x6) : (~x4 | ~x6)))));
  assign n490 = ~x1 & (n491 | (~x2 & x7 & ~n494));
  assign n491 = ~x7 & (x0 ? ~n493 : ~n492);
  assign n492 = (x2 | ~x3 | x4 | ~x5 | x6) & (~x2 | x3 | ~x4 | x5 | ~x6);
  assign n493 = (~x2 | x3 | ~x4 | x5 | x6) & (x2 | ~x3 | ~x6 | (x4 ^ x5));
  assign n494 = (x0 | x3 | ~x4 | ~x5 | x6) & (~x0 | x4 | (x3 ? (~x5 | ~x6) : (x5 | x6)));
  assign n495 = x0 ? ((~x2 | x3 | x4 | ~x5) & (~x4 | x5 | x2 | ~x3)) : ((x2 | x3 | x4 | ~x5) & (~x3 | (x5 ? ~x2 : x4)));
  assign n496 = ~n501 & (~n155 | (n497 & n500));
  assign n497 = (x6 | n499) & (~x4 | ~x6 | ~x7 | n498);
  assign n498 = x2 ? (x3 | x5) : (~x3 | ~x5);
  assign n499 = x2 ? (~x3 | ~x5 | (x4 ^ ~x7)) : (x3 | x5 | (x4 ^ x7));
  assign n500 = (~x2 | x3 | (x4 ^ x5)) & (~x3 | (x2 ? (~x4 | x5) : (x4 | ~x5)));
  assign n501 = n226 & ((~x3 & ~x4 & x5 & ~x6) | ((x3 ^ x6) & (~x4 ^ x5)));
  assign z017 = ~n513 | (~x0 & (~n506 | (~x1 & ~n503)));
  assign n503 = (x2 | n504) & (~x2 | x3 | ~x5 | n505);
  assign n504 = (x3 | x4 | ~x5 | x6) & (~x4 | ((~x3 | ~x6 | (~x5 & ~x7)) & (x6 | x7 | x3 | x5)));
  assign n505 = x4 ? (x6 | x7) : ~x6;
  assign n506 = ~n509 & n512 & (~x1 | (n507 & n511));
  assign n507 = (~n249 | ~n252) & (n236 | n508);
  assign n508 = ~x2 ^ x5;
  assign n509 = n510 & ((x2 & ~x3 & (~x6 ^ x7)) | (x3 & (x2 ? (~x6 & x7) : (x6 & ~x7))));
  assign n510 = ~x1 & ~x5;
  assign n511 = (x2 | ~x3 | x5 | ~x6 | x7) & (~x2 | x3 | ~x5 | x6 | ~x7);
  assign n512 = (x1 | ~x2 | ~x3 | x6 | x7) & (~x1 | ((~x6 | ~x7 | x2 | ~x3) & (x6 | x7 | ~x2 | x3)));
  assign n513 = ~n516 & (n183 | (~n515 & (x1 | n514)));
  assign n514 = (x0 | x2 | x3 | ~x4) & ((x2 ^ x4) | (x0 ? (x3 | x5) : (~x3 | ~x5)));
  assign n515 = n155 & (x2 ? (x3 & (x5 | n382)) : (~x3 & ~x5));
  assign n516 = n268 & (~n518 | (~x2 & ~n517));
  assign n517 = (~x5 & (x4 ? x3 : ~x7)) | (~x3 & x5) | (x6 & ~x7) | (~x6 & x7);
  assign n518 = (~x2 | x3 | x4 | x6) & (x2 | ((x3 | ~x5 | ~x6) & (~x3 | ~x4 | x5 | x6)));
  assign z018 = n528 | ~n531 | (~x1 & ~n520);
  assign n520 = x6 ? (n522 & (~n279 | ~n521)) : n525;
  assign n521 = x7 & (x2 ? (x4 & x5) : (~x4 & ~x5));
  assign n522 = (n283 | n524) & (~n523 | ~n386);
  assign n523 = ~x7 & ~x4 & ~x5;
  assign n524 = (~x0 | ~x2 | x3 | x4) & (x0 | x2 | ~x3 | ~x4);
  assign n525 = x5 ? (~n203 | n527) : n526;
  assign n526 = (x4 | x7 | x2 | ~x3) & (x3 | (x0 ? (x2 | ~x7) : ((x4 | ~x7) & (x2 | ~x4 | x7))));
  assign n527 = x3 ? (~x4 ^ x7) : (~x4 | ~x7);
  assign n528 = x3 & ((n203 & ~n530) | (~x2 & ~n529));
  assign n529 = (x0 | ((~x5 | x7 | x1 | ~x4) & (~x1 | ((x5 | x7) & (~x4 | ~x5 | ~x7))))) & (x1 | ((~x7 | ((x4 | ~x5) & (~x0 | (x4 & ~x5)))) & (x5 | x7 | ~x0 | ~x4)));
  assign n530 = x1 ? (~x5 | ~x7) : (x5 | x7);
  assign n531 = ~n536 & (x3 | (n533 & (x2 | n532)));
  assign n532 = (x0 | ~x7 | (x1 ? (x4 | x5) : (~x4 | ~x5))) & (~x0 | x1 | ~x5 | x7);
  assign n533 = (x1 | ~x2 | n535) & (x0 | (n535 & (~x1 | ~x2 | ~n534)));
  assign n534 = x4 & x5 & ~x7;
  assign n535 = x4 ? (x5 | ~x7) : (~x5 | x7);
  assign n536 = n155 & ((n538 & ~n540) | (~n537 & ~n539));
  assign n537 = ~x4 ^ x7;
  assign n538 = x2 & ~x5;
  assign n539 = (~x2 | ~x3 | x5 | ~x6) & (x2 | ~x5 | (~x3 ^ x6));
  assign n540 = (x3 | x4 | x6 | ~x7) & (~x3 | (x4 ? (~x6 | ~x7) : (x6 | x7)));
  assign z019 = x0 ? (~x1 & ~n542) : (x1 ? ~n550 : ~n546);
  assign n542 = ~n544 & (x4 ? (~x5 | n545) : n543);
  assign n543 = (x2 & (x3 | x7)) | (~x5 & x6) | (~x6 & (x3 ? x7 : (x5 & ~x7)));
  assign n544 = ~n374 & (x2 ? ~x3 : (x3 & x7));
  assign n545 = (~x2 | x3 | x6 | x7) & (x2 | (~x6 & (~x3 | ~x7)));
  assign n546 = (x7 | n549) & (~x7 | n547) & (n537 | n548);
  assign n547 = (~x2 | x5 | ~x6 | (~x3 & ~x4)) & (~x4 | ~x5 | ((x2 | x3) & x6));
  assign n548 = (x2 | ((~x5 | ~x6) & (x3 | x5 | x6))) & (~x5 | (x6 ? x3 : ~x2));
  assign n549 = (x2 | ~x3 | ~x4 | x6) & (x4 | ((~x6 | (x3 & ~x5)) & (~x2 | (~x6 & (~x3 | ~x5)))));
  assign n550 = ~n551 & ~n552 & (x2 | n355) & ~n553;
  assign n551 = x4 & ((~x2 & (x5 ? (~x6 & ~x7) : x6)) | (x6 & ((x2 & x5 & x7) | (~x5 & ~x7))));
  assign n552 = n538 & ((x3 & x4 & ~x6 & ~x7) | (~x3 & (x4 ? x7 : (x6 & ~x7))));
  assign n553 = ~x4 & ((x2 & (~x5 ^ x6)) | (~x5 & (x6 ? ~x2 : x7)));
  assign z020 = ~n561 | (~x1 & ~n555);
  assign n555 = x2 ? n558 : (~n557 & (~x0 | n556));
  assign n556 = (x3 | (x4 ? (~x5 | x6) : (~x6 | ~x7))) & (x5 | x7 | (x4 ^ x6)) & (~x6 | ~x7 | ~x3 | ~x5);
  assign n557 = n238 & (x6 ? ~n229 : ~n537);
  assign n558 = x0 ? (~n158 | ~n559) : n560;
  assign n559 = x7 & x5 & ~x6;
  assign n560 = x6 ? ((~x4 | x5 | x7) & (x3 | (x4 ^ ~x7))) : ((~x4 | ~x5 | ~x7) & (~x3 | x4 | x5));
  assign n561 = ~n562 & n569 & (n416 | (~n565 & n566));
  assign n562 = n155 & (x4 ? ~n563 : ~n564);
  assign n563 = (~x3 | (x2 ? (~x5 | (x6 ^ ~x7)) : (x6 | x7))) & (x2 | (x5 ? (~x6 | ~x7) : (x6 | x7)));
  assign n564 = (x2 | ~x3 | ~x5 | x6 | ~x7) & (x3 | ((x6 | x7 | x2 | x5) & (~x2 | (x5 ? (x6 | ~x7) : (~x6 | x7)))));
  assign n565 = ~n281 & ((~x0 & x1 & ~x2 & ~x3) | (~x1 & (x0 ? (x2 ^ x3) : (x2 & x3))));
  assign n566 = x0 ? (~n209 | ~n567) : n568;
  assign n567 = ~x6 & ~x3 & ~x4;
  assign n568 = x2 ? ((~x1 | (x3 ? (x4 | x6) : (~x4 | ~x6))) & (x4 | x6 | x1 | x3)) : (x1 ? (~x3 | ~x6) : ((~x3 | x4 | x6) & (~x4 | ~x6)));
  assign n569 = (~n570 | n571) & (~n572 | (x1 ^ x2));
  assign n570 = ~x5 & ~x7;
  assign n571 = (~x0 | x1 | ~x2 | x3 | x4) & (x0 | ((~x3 | ~x4 | x1 | x2) & (~x1 | (x2 ? ~x4 : (~x3 | x4)))));
  assign n572 = x7 & ~x4 & ~x0 & x3 & x5;
  assign z021 = n574 | n579 | ~n586 | (~n582 & n585);
  assign n574 = ~x7 & (n576 | (~n575 & (~x3 ^ x4)));
  assign n575 = (~x0 | x1 | x2 | ~x5 | ~x6) & (x0 | x5 | (x1 ? (x2 | ~x6) : (~x2 | x6)));
  assign n576 = ~x0 & ((x1 & ~n577) | (n205 & ~n578));
  assign n577 = (~x2 | ~x4 | x6 | (x3 ^ x5)) & (x2 | x3 | x4 | ~x5 | ~x6);
  assign n578 = (~x2 | x4 | ~x5 | x6) & (x2 | x5 | ~x6);
  assign n579 = ~n416 & (n581 | (~x3 & ~n580));
  assign n580 = (x1 | ((~x4 | x6 | x0 | ~x2) & (~x0 | x4 | (x2 ^ x6)))) & (x0 | ~x1 | ((~x2 | x4 | x6) & (~x4 | (x2 & ~x6))));
  assign n581 = x6 & x3 & ~x2 & ~x0 & ~x1;
  assign n582 = (x1 | n583) & (~x1 | ~x3 | ~x6 | n584);
  assign n583 = (~x3 | x6 | ((x4 | ~x5) & (~x2 | (x4 & ~x5)))) & (x2 | x3 | ~x5 | ~x6);
  assign n584 = (x4 | x5) & (x2 | ~x4 | ~x5);
  assign n585 = ~x0 & x7;
  assign n586 = ~n587 & ~n589 & ~n592 & (n336 | n593);
  assign n587 = x3 & n155 & ~n588;
  assign n588 = (x2 | x4 | x5 | x6) & (~x5 | (x2 ? (~x4 | ~x6) : (~x4 ^ x6)));
  assign n589 = ~n591 & (x3 ? (n570 | (~x4 & n590)) : (x4 & n590));
  assign n590 = x5 & x7;
  assign n591 = (~x0 | x1 | x2) & (x0 | ~x1 | ~x2 | x6);
  assign n592 = n205 & ((x0 & x2 & ~x5 & ~x6) | (~x0 & x5 & (~x2 ^ x6)));
  assign n593 = (~n472 | ~n594) & (x0 | n283 | n595);
  assign n594 = x7 & x4 & ~x5;
  assign n595 = x1 ? (x3 | x4) : (~x3 | ~x4);
  assign z022 = n597 | ~n603 | ~n611 | (~n183 & ~n602);
  assign n597 = ~x1 & ((n598 & ~n601) | (~x3 & ~n599));
  assign n598 = x3 & x7;
  assign n599 = (~x5 | n600) & (x0 | x5 | ~n266 | ~n338);
  assign n600 = (x0 | ~x2 | x4 | ~x6 | x7) & (~x0 | ((~x6 | ~x7 | x2 | x4) & (~x2 | ~x4 | x6 | x7)));
  assign n601 = (~x0 | x2 | ~x4 | x5 | ~x6) & (x0 | x6 | (x2 ? (~x4 | x5) : (x4 | ~x5)));
  assign n602 = (~x0 | x1 | x2 | x3 | x4) & (x0 | ~x2 | (x1 ? (~x3 | ~x4) : (x3 ^ ~x4)));
  assign n603 = ~n606 & (n604 | ~n605) & (x0 | n608);
  assign n604 = (~x2 | ~x3 | x4 | (~x5 ^ ~x6)) & (x2 | x3 | ~x4 | x5 | ~x6);
  assign n605 = ~x7 & ~x0 & x1;
  assign n606 = n607 & (x2 ? ~x6 : (~x4 & x6));
  assign n607 = ~x3 & ~x0 & x1;
  assign n608 = x1 ? (~x7 | n610) : (~n293 | ~n609);
  assign n609 = ~x7 & ~x4 & ~x6;
  assign n610 = (~x2 | ~x3 | x4 | x6) & (x2 | x3 | ~x4 | ~x6);
  assign n611 = (n300 | n613) & (x1 | (n614 & (n300 | n612)));
  assign n612 = (x0 | x2 | x3 | x4 | ~x5) & (~x0 | ~x4 | (x2 ? (x3 | x5) : (~x3 | ~x5)));
  assign n613 = (~x0 | x1 | ~x2 | x3 | x4) & (x0 | x2 | (x1 ? ~x3 : (x3 | ~x4)));
  assign n614 = (x2 | ((~x4 | x6 | x0 | ~x3) & (~x0 | ~x6 | (~x3 ^ x4)))) & (x0 | ~x2 | (x3 ? (~x4 | ~x6) : (x4 | x6)));
  assign z023 = n618 | ~n625 | (~x1 & (~n616 | ~n624));
  assign n616 = (~x0 | ~x4 | x7 | n498) & (x0 | (n617 & (x4 | ~x7 | n498)));
  assign n617 = (x2 | x4 | x7 | (~x3 ^ x5)) & (~x2 | ~x3 | ~x4 | ~x5 | ~x7);
  assign n618 = ~x1 & (~n620 | (~n183 & ~n619));
  assign n619 = (~x0 | x2 | ~x3 | ~x4 | x5) & (x0 | ~x2 | x3 | x4 | ~x5);
  assign n620 = (n621 | n622) & (~x6 | ~n146 | n623);
  assign n621 = x0 ? (x3 | ~x5) : (~x3 | x5);
  assign n622 = (~x2 | ~x4 | x6 | x7) & (x2 | x4 | ~x6 | ~x7);
  assign n623 = (x2 | x3 | x4 | x7) & (~x2 | ~x3 | ~x4 | ~x7);
  assign n624 = x0 ? ((x3 | x4 | x7) & (x2 | ~x7 | (~x3 ^ x4))) : (x3 ? (x2 ? (x4 | x7) : (~x4 | ~x7)) : (~x4 | x7));
  assign n625 = (~n368 | ~n626) & (~n155 | (n627 & n628));
  assign n626 = ~x2 & ~x0 & x1 & ~x3;
  assign n627 = (x2 | x3 | ~x4 | x5 | ~x7) & (~x2 | ~x3 | x4 | (x5 ^ ~x7));
  assign n628 = x7 ? (x3 | (~x2 & x4)) : (~x3 | (x2 & ~x4));
  assign z024 = ~n642 | n639 | n637 | n630 | n634;
  assign n630 = ~x1 & ((n631 & n633) | (~x5 & ~n632));
  assign n631 = x6 & ~x4 & x5;
  assign n632 = x0 ? ((~x4 | ~x6 | x2 | ~x3) & (x4 | x6 | ~x2 | x3)) : ((~x2 | ~x3 | ~x4 | ~x6) & (x2 | x3 | (x4 ^ ~x6)));
  assign n633 = ~x3 & ~x0 & x2;
  assign n634 = n279 & ((n334 & ~n636) | (n448 & n635));
  assign n635 = ~x4 & ~x1 & ~x2;
  assign n636 = (x1 | x2 | ~x4 | x6) & (~x1 | (x2 ? (~x4 | x6) : (x4 | ~x6)));
  assign n637 = ~x0 & ~n638;
  assign n638 = (x5 | ((x1 | x2 | ~x3 | ~x4) & (~x1 | (x2 ? (~x3 | ~x4) : x4)))) & (x1 | x2 | x4 | ~x5);
  assign n639 = ~x3 & (n640 | (n382 & n383 & n462));
  assign n640 = ~n641 & (x2 ? n570 : n590);
  assign n641 = (~x0 | x1 | x4 | ~x6) & (x0 | ~x1 | ~x4 | x6);
  assign n642 = (n643 | ~n645) & (n644 | (x3 & ~x5));
  assign n643 = x3 ? (x4 | x6) : (~x4 | ~x6);
  assign n644 = (~x0 | x1 | x2 | ~x4) & (x0 | ~x2 | (~x1 ^ x4));
  assign n645 = ~x2 & ~x0 & x1 & x5;
  assign z025 = n652 | n656 | (~x1 & ~n647) | n661;
  assign n647 = x2 ? n650 : (x3 ? n649 : n648);
  assign n648 = (~x6 | ((x0 | ~x4 | ~x5 | x7) & (~x0 | (x4 ? (x5 | x7) : (~x5 | ~x7))))) & (x0 | x4 | x6 | (x5 ^ ~x7));
  assign n649 = (~x0 | x4 | ~x5 | x6 | x7) & (x0 | ~x7 | (x4 ? (~x5 | x6) : (x5 | ~x6)));
  assign n650 = x0 ? (~n448 | ~n158) : (x7 | n651);
  assign n651 = (x3 | ~x4 | x5 | ~x6) & (~x3 | ~x5 | (x4 ^ x6));
  assign n652 = n155 & ((n653 & ~n655) | (x5 & ~n654));
  assign n653 = x4 & ~x5;
  assign n654 = (~x7 | ((~x2 | ~x3 | ~x4 | x6) & (x2 | (x3 ? (x4 | ~x6) : (~x4 | x6))))) & (~x2 | x3 | x7 | (x4 ^ x6));
  assign n655 = (x2 | ~x3 | ~x6 | x7) & (~x2 | x6 | (~x3 ^ x7));
  assign n656 = ~x4 & (~n658 | (~x0 & ~n657));
  assign n657 = (~x1 | x2 | ~x3 | x5 | x6) & (x1 | x3 | (x2 ? (~x5 ^ ~x6) : (x5 | ~x6)));
  assign n658 = ~n659 & ~n660 & (x3 | ~n157 | ~n159);
  assign n659 = ~x1 & (x0 ? (x2 ? (~x3 & x5) : (x3 & ~x5)) : (x3 & (~x2 ^ ~x5)));
  assign n660 = ~x0 & x1 & (x2 ? (x3 ^ ~x5) : (~x3 & x5));
  assign n661 = x4 & (~n663 | (~x0 & ~n662));
  assign n662 = x1 ? ((~x2 | ~x3 | ~x5 | ~x6) & (x2 | (x3 ? (x5 | x6) : (~x5 | ~x6)))) : ((~x5 | ~x6 | x2 | ~x3) & (x5 | x6 | ~x2 | x3));
  assign n663 = x5 ? (x6 | n664) : ((~x6 | n664) & (x3 | x6 | ~n157));
  assign n664 = (~x0 | x1 | x2 | ~x3) & (x0 | (x1 ? (~x2 | x3) : (x2 ^ x3)));
  assign z026 = ~n666 | (x5 ? ~n682 : ~n674);
  assign n666 = ~n667 & n671 & (n413 | n670);
  assign n667 = ~x1 & ((n203 & ~n669) | (~x2 & ~n668));
  assign n668 = x3 ? ((~x4 | ~x5 | ~x6) & (~x0 | x4 | x5 | x6)) : ((x5 | ~x6 | x0 | ~x4) & (~x0 | (x4 ? (~x5 | x6) : (x5 | ~x6))));
  assign n669 = x3 ? (x5 | (x4 ^ x6)) : (x4 ? (~x5 | x6) : ~x6);
  assign n670 = (~x0 | x1 | x2 | ~x3 | x4) & (x0 | ((~x1 | ~x2 | x3 | x4) & (x1 | ~x3 | (x2 ^ ~x4))));
  assign n671 = (~n155 | n673) & (n223 | n672);
  assign n672 = (x1 | ((~x3 | x6 | x0 | x2) & (~x0 | (x2 ? (x3 | x6) : (~x3 | ~x6))))) & (x0 | ~x1 | x3 | (x2 ^ x6));
  assign n673 = (x4 | ((x2 | ~x3 | x5 | ~x6) & (~x2 | x6 | (x3 ^ x5)))) & (x2 | ~x3 | ~x4 | ~x5 | x6);
  assign n674 = ~n676 & ~n678 & (~n141 | ~n155 | ~n675);
  assign n675 = ~x6 & (x4 ^ ~x7);
  assign n676 = ~n300 & ~n677;
  assign n677 = (x0 | ~x1 | x2 | ~x3 | ~x4) & (x1 | ((~x3 | x4 | x0 | x2) & (x3 | (x0 ? (x2 ^ ~x4) : (~x2 | ~x4)))));
  assign n678 = ~x3 & ((n679 & ~n681) | (n231 & n680));
  assign n679 = ~x0 & ~x6;
  assign n680 = x4 & x6 & ~x7;
  assign n681 = (x1 | x2 | x4 | ~x7) & (~x1 | (x2 ? (~x4 | ~x7) : (x4 | x7)));
  assign n682 = (x0 | n683) & (~x0 | ~n266 | ~n209 | ~n158);
  assign n683 = (~x7 | n685) & (n684 | (x2 ^ x3));
  assign n684 = (x1 | x4 | ~x6 | x7) & (~x4 | (x1 ? (~x6 ^ x7) : (~x6 | ~x7)));
  assign n685 = (~x1 | ~x6 | (x2 ? (x3 | ~x4) : (~x3 | x4))) & (x1 | x2 | x3 | x4 | x6);
  assign z027 = n687 | ~n708 | (x2 ? ~n690 : ~n699);
  assign n687 = ~x0 & (x1 ? ~n688 : ~n689);
  assign n688 = (x4 | (x2 ? (x3 ? (~x5 | x7) : (x5 | ~x7)) : (x7 | (~x3 ^ x5)))) & (x2 | ~x4 | (x3 ? (x5 | ~x7) : (~x5 ^ ~x7)));
  assign n689 = (x2 | ~x3 | x4 | x5 | ~x7) & (x3 | (x2 ? (~x4 | (x5 ^ ~x7)) : (~x5 | ~x7)));
  assign n690 = ~n696 & (x3 | (~n691 & (~n155 | n695)));
  assign n691 = ~x1 & ((n692 & n693) | (n312 & n694));
  assign n692 = x0 & x4;
  assign n693 = ~x7 & ~x5 & ~x6;
  assign n694 = x5 & x6 & x7;
  assign n695 = (~x4 | x5 | x6 | ~x7) & (x4 | ~x5 | (~x6 ^ x7));
  assign n696 = ~n697 & n698;
  assign n697 = x4 ? (~x6 | x7) : (x6 | ~x7);
  assign n698 = ~x5 & x3 & ~x0 & x1;
  assign n699 = ~n705 & (x7 | (~n701 & (~x5 | n700)));
  assign n700 = (x0 | x1 | ~x3 | x4 | ~x6) & ((x0 ? (x1 | x3) : (~x1 | ~x3)) | (~x4 ^ ~x6));
  assign n701 = n510 & (n704 | (~x0 & (n702 | n703)));
  assign n702 = x3 & x4 & ~x6;
  assign n703 = x6 & ~x3 & ~x4;
  assign n704 = x6 & x4 & x0 & ~x3;
  assign n705 = n707 & (n706 | (~x3 & ~x5 & ~n446));
  assign n706 = ~x6 & x5 & x3 & ~x4;
  assign n707 = x7 & ~x0 & x1;
  assign n708 = ~n709 & ~n712 & n714 & (~x3 | n713);
  assign n709 = ~n244 & ((n169 & ~n711) | (n157 & n710));
  assign n710 = x7 & x3 & ~x4;
  assign n711 = (x1 | x2 | ~x3 | ~x7) & (x7 | (x1 ? (~x2 | x3) : (x2 ^ x3)));
  assign n712 = n254 & ((x2 & ((~x5 & x7) | (~x4 & x5 & ~x7))) | (x4 & ~x5 & x7) | (~x2 & ~x4 & (~x5 ^ x7)));
  assign n713 = (~x0 | x1 | x2 | ~x4 | x7) & (x0 | ~x2 | ~x7 | (x1 ^ x4));
  assign n714 = (~n193 | ~n715) & (n718 | (~n716 & ~n717));
  assign n715 = ~x7 & ~x3 & ~x4;
  assign n716 = x4 & x5 & x6 & x7;
  assign n717 = ~x7 & ~x6 & ~x4 & ~x5;
  assign n718 = (~x0 | x1 | x2 | ~x3) & (x0 | ~x2 | (~x1 ^ x3));
  assign z028 = n729 | n732 | (~x1 & ~n720);
  assign n720 = ~n721 & ~n724 & (x4 ? n728 : n727);
  assign n721 = x3 & ((n722 & n694) | (~x2 & ~n723));
  assign n722 = ~x4 & ~x0 & x2;
  assign n723 = (~x0 | ((~x4 | x5 | x6 | ~x7) & (~x5 | ~x6 | x7))) & (x0 | x4 | x5 | x6 | ~x7) & (~x5 | ((~x4 | ~x6 | x7) & (x0 | x6 | (~x4 ^ ~x7))));
  assign n724 = ~x3 & (x0 ? ~n726 : ~n725);
  assign n725 = (x6 | ((x2 | (x4 ? (~x5 | x7) : (x5 | ~x7))) & (~x2 | x4 | ~x5 | ~x7))) & (~x2 | ~x6 | (x4 ? (~x5 | ~x7) : x7));
  assign n726 = (~x4 | ~x5 | x6 | x7) & (x5 | ~x7 | (x2 ? (x4 | x6) : (~x4 ^ x6)));
  assign n727 = (~x0 | (x2 ? (x3 | ~x6) : (~x3 | x6))) & (x0 | x2 | x3 | ~x6);
  assign n728 = (x0 | ~x2 | x3 | x5 | ~x6) & (~x3 | ((x2 | (x0 ? (x5 ^ ~x6) : (x5 | x6))) & (x0 | ~x2 | ~x5 | x6)));
  assign n729 = ~n300 & ((n254 & ~n731) | (~x0 & ~n730));
  assign n730 = (x2 | ((~x1 | ~x3 | ~x5) & (~x4 | x5 | x1 | x3))) & (x1 | ~x3 | x5 | (~x2 & x4));
  assign n731 = (~x4 | x5) & (x2 | x4 | ~x5);
  assign n732 = n155 & (~n734 | ~n735 | (n176 & ~n733));
  assign n733 = x2 ? (x5 | x6) : (~x5 | ~x6);
  assign n734 = (x2 & ~x5 & (~x6 | x7)) | (x3 & ~x6) | (~x3 & x6) | (~x2 & x5);
  assign n735 = ~n738 & (x5 | x6 | ~n736 | n737);
  assign n736 = x2 & ~x4;
  assign n737 = x3 ^ x7;
  assign n738 = ~x2 & ~x3 & (x5 ? (~x6 & x7) : (x6 & ~x7));
  assign z029 = ~n748 | (~x1 & (~n740 | ~n745));
  assign n740 = x2 ? n743 : (n742 & (~x6 | n741));
  assign n741 = (~x0 | ~x4 | ~x7 | (~x3 ^ x5)) & (x4 | x5 | ((x3 | x7) & (x0 | (x3 & x7))));
  assign n742 = (~x0 | ((x3 | x5 | x6 | ~x7) & (~x3 | ~x5 | ~x6 | x7))) & (x0 | ~x3 | x5 | x6 | ~x7);
  assign n743 = x0 ? (~n174 | ~n176) : n744;
  assign n744 = (~x5 | (~x3 ^ x4) | (x6 ^ ~x7)) & (x3 | x5 | x6 | (x4 & x7));
  assign n745 = x0 ? n746 : n747;
  assign n746 = (x2 | ~x3 | x5 | (x4 ^ ~x7)) & (x3 | (x2 ? (x4 ? (x5 | x7) : (~x5 | ~x7)) : (~x5 | x7)));
  assign n747 = x3 ? ((~x5 | x7 | x2 | ~x4) & (~x2 | ((x5 | x7) & (~x4 | ~x5 | ~x7)))) : (x2 ? (x4 ? (x5 | ~x7) : (~x5 | x7)) : (x4 ? (x5 | x7) : (~x5 | ~x7)));
  assign n748 = ~n749 & ~n753 & (~n155 | n752);
  assign n749 = n155 & (x3 ? ~n751 : ~n750);
  assign n750 = x2 ? (x6 | ((~x5 | ~x7) & (~x4 | x5 | x7))) : (~x6 | ((~x4 | ~x5 | ~x7) & (x5 | x7)));
  assign n751 = (x2 | x4 | ~x5 | ~x6 | ~x7) & (~x2 | ((x6 | x7 | x4 | ~x5) & (~x4 | x5 | (x6 ^ ~x7))));
  assign n752 = (~x4 | ((x2 | ~x5 | x7) & (~x2 | x3 | x5 | ~x7))) & (~x3 | (x2 ? ((~x5 | ~x7) & (x4 | x5 | x7)) : (x5 ^ ~x7)));
  assign n753 = ~n300 & ((n231 & n351) | (~x0 & ~n754));
  assign n754 = (x1 | x2 | ~x3 | x4 | ~x5) & (x3 | ((x1 | x2 | ~x4 | ~x5) & (~x1 | x4 | (x2 ^ ~x5))));
  assign z030 = n766 | n771 | (~x1 & (n756 | ~n759));
  assign n756 = ~x0 & (n758 | (~x3 & ~n757));
  assign n757 = (~x2 | x4 | x5 | ~x6 | x7) & (~x4 | ((~x5 | ~x6 | ~x7) & (x6 | x7 | x2 | x5)));
  assign n758 = ~x7 & n305 & (x2 ? ~x6 : (~x4 & x6));
  assign n759 = ~n762 & (x2 | (n760 & n761)) & n765;
  assign n760 = (x3 | x4 | ~x5 | x6 | x7) & (~x3 | x5 | (x4 ? (~x6 | ~x7) : (x6 | x7)));
  assign n761 = (x0 | x3 | ~x4 | ~x6 | x7) & (~x0 | ~x7 | (x3 ? (x4 | x6) : (~x4 | ~x6)));
  assign n762 = x6 & n764 & (n763 | (n653 & n164));
  assign n763 = x5 & ~x2 & x3;
  assign n764 = x0 & ~x7;
  assign n765 = (~n174 | ~n464) & (x3 | ~n203 | n697);
  assign n766 = ~n281 & (~n768 | (n767 & ~n427));
  assign n767 = x3 & x5;
  assign n768 = ~n770 & (x1 ? (x0 | ~n763) : n769);
  assign n769 = x0 ? (x3 | x5) : (~x3 | ~x5);
  assign n770 = x7 & ~x5 & ~x0 & ~x3;
  assign n771 = n155 & (n772 | ~n776 | (~n219 & ~n775));
  assign n772 = n773 & n774;
  assign n773 = x3 & ~x4;
  assign n774 = ~x6 & (x2 ? ~x5 : (x5 & x7));
  assign n775 = (~x4 | ~x6) & (x2 | x4 | x6);
  assign n776 = ~n777 & (~n457 | ~n164) & (~n249 | ~n694);
  assign n777 = (x3 ^ x6) & (x2 ? (x5 & x7) : (~x5 & ~x7));
  assign z031 = ~n794 | n792 | n789 | n779 | n782;
  assign n779 = ~n300 & (~n781 | (x4 & ~n780));
  assign n780 = (x0 | ((~x2 | ~x3 | ~x5) & (x1 | (x2 ^ x5)))) & (x1 | x2 | ((~x3 | x5) & (~x0 | x3 | ~x5)));
  assign n781 = (~x0 | x1 | ~x2 | x3 | x5) & (x0 | ~x1 | ~x5 | (x2 & x3));
  assign n782 = ~x2 & (n783 | n786);
  assign n783 = ~x1 & ((x3 & ~n784) | (n238 & n785));
  assign n784 = x0 ? ((~x4 | ~x5 | ~x7) & (x6 | x7 | x4 | x5)) : ((~x6 | ~x7 | x4 | x5) & (~x4 | ~x5 | x6 | x7));
  assign n785 = x7 & (x4 ? (~x5 & ~x6) : (x5 ^ x6));
  assign n786 = n787 & n155 & (n788 | n158);
  assign n787 = x6 & ~x7;
  assign n788 = x3 & x4 & ~x5;
  assign n789 = ~x0 & (~n791 | (x7 & n510 & ~n790));
  assign n790 = x2 ? (x3 | ~x6) : (~x3 | x6);
  assign n791 = (x1 | ((~x2 | x5 | x6 | ~x7) & (~x5 | ~x6 | x7))) & (~x1 | x2 | x5 | x6 | ~x7);
  assign n792 = n203 & (x1 ? ~n793 : (n174 & n773));
  assign n793 = (~x3 | ((~x6 | ~x7 | x4 | ~x5) & (x6 | x7 | ~x4 | x5))) & (x3 | ~x4 | x5 | x6 | ~x7);
  assign n794 = (n413 | n796) & (~n191 | ~n795 | ~n157);
  assign n795 = ~x3 & ~x5;
  assign n796 = x0 ? (x1 | ((x3 | x4) & (x2 | (x3 & x4)))) : (~x1 | (~x2 & (~x3 | x4)));
  assign z032 = ~n806 | (~x1 & (n798 | n801 | ~n803));
  assign n798 = ~x2 & (x3 ? ~n799 : ~n800);
  assign n799 = (x6 | (~x4 ^ x5) | (~x0 ^ ~x7)) & (~x0 | ~x6 | (x4 ? ~x5 : (x5 | ~x7)));
  assign n800 = x0 ? ((~x6 | ~x7 | x4 | x5) & (~x4 | x6 | (x5 ^ ~x7))) : (~x5 | (x4 ? (~x6 | x7) : (~x6 ^ ~x7)));
  assign n801 = x2 & (x0 ? (n176 & n339) : ~n802);
  assign n802 = (x3 | ((x6 | x7 | x4 | ~x5) & (~x6 | ~x7 | ~x4 | x5))) & (~x7 | (x4 ? (~x5 | x6) : ((x5 | x6) & (~x3 | ~x5 | ~x6))));
  assign n803 = (n537 | n804) & (~x6 | n805);
  assign n804 = (x0 | x2 | ~x3 | ~x6) & (x3 | (x0 ? (~x2 | x6) : (x2 ^ x6)));
  assign n805 = x2 ? (x7 | (x3 ? x0 : x4)) : ((~x0 | x7 | (x3 & x4)) & (~x4 | ~x7 | (x0 & x3)));
  assign n806 = ~n155 | (n807 & (x2 ? n808 : n809));
  assign n807 = (x6 | ((x3 | (x2 ^ ~x7)) & (x2 | (x4 ^ x7)))) & (~x2 | ~x6 | ~x7 | (~x3 & x4));
  assign n808 = (~x3 | ~x4 | ~x5 | x6 | x7) & ((x5 ^ x6) | (x3 ? (x4 | x7) : (~x4 | ~x7)));
  assign n809 = x3 ? (x6 | (x4 ? (~x5 | x7) : (x5 | ~x7))) : (~x6 | x7 | (~x4 ^ x5));
  assign z033 = ~n812 | ~n816 | (~n811 & (n155 | n268));
  assign n811 = (x3 | ((~x2 | (x4 ? (x5 | ~x7) : x7)) & (x5 | x7 | x2 | ~x4))) & (x2 | (x4 ? (~x5 | ~x7) : ((x5 | ~x7) & (~x3 | ~x5 | x7))));
  assign n812 = ~n813 & (x5 | ~n279 | n815);
  assign n813 = ~n300 & (x0 ? (n788 & n209) : ~n814);
  assign n814 = (~x4 | x5 | x2 | ~x3) & (x1 | ~x2 | x3 | x4 | ~x5);
  assign n815 = (x1 | x2 | x4 | x6 | ~x7) & (~x2 | ~x4 | (x6 ^ ~x7));
  assign n816 = ~n820 & (x0 | (n818 & (x1 | n817)));
  assign n817 = ((x4 ^ x7) | (x2 ? (x3 | x5) : (~x3 | ~x5))) & (x2 | x3 | x4 | x5 | ~x7) & (~x2 | ~x3 | ~x4 | ~x5 | x7);
  assign n818 = (n283 | n819) & (~x1 | ~n141 | ~n534);
  assign n819 = (~x2 | ~x3 | x4) & (x1 | x2 | x3 | ~x4);
  assign n820 = n304 & ((~n537 & ~n821) | (x6 & ~n822));
  assign n821 = (x1 | x2 | x6) & (x0 | ((x2 | x6) & (~x1 | ~x2 | ~x6)));
  assign n822 = (~x0 | x1 | ~x2 | x4 | ~x7) & (x0 | x7 | ((x2 | x4) & (x1 | ~x2 | ~x4)));
  assign z034 = ~n832 | (~x1 & (~n827 | (x5 & ~n824)));
  assign n824 = (~x2 | n826) & (~x0 | x2 | n737 | ~n825);
  assign n825 = ~x4 & x6;
  assign n826 = (~x0 | x3 | x4 | ~x6 | x7) & (x0 | ~x3 | ~x4 | x6 | ~x7);
  assign n827 = ~n830 & (~n828 | ~n559) & (x3 | n829);
  assign n828 = x4 & ~x2 & x3;
  assign n829 = (~x2 | x4 | x5 | ~x6 | ~x7) & (~x4 | ~x5 | x6 | x7);
  assign n830 = x6 & n382 & n401 & ~n831;
  assign n831 = ~x3 ^ x7;
  assign n832 = ~n833 & ~n835 & (~x3 | (~n836 & ~n838));
  assign n833 = x5 & n155 & ~n834;
  assign n834 = x3 ? (~x7 | (~x4 ^ x6)) : (x7 | ((~x2 | x4 | ~x6) & (~x4 | x6)));
  assign n835 = ~x3 & (~x0 | ~x1) & ~n374;
  assign n836 = ~n837 & ((~x1 & n151) | (~x0 & (~x1 | x4)));
  assign n837 = x5 ^ x6;
  assign n838 = n382 & (~n839 | (n140 & n240));
  assign n839 = x0 ? (x1 | x2) : ~x1;
  assign z035 = ~n850 | n841 | n843;
  assign n841 = n268 & ((x7 & ~n842) | (~x2 & n534));
  assign n842 = (x6 | (x2 & x3) | (~x4 ^ x5)) & (x2 | ~x6 | ((x4 | x5) & (~x3 | ~x4 | ~x5)));
  assign n843 = ~x0 & (x1 ? (n785 | n844) : ~n847);
  assign n844 = ~x7 & ((n845 & n393) | (n141 & n846));
  assign n845 = ~x2 & ~x3;
  assign n846 = x4 & x5 & ~x6;
  assign n847 = n849 & (~x7 | ~n773 | n848);
  assign n848 = x2 ? (x5 | ~x6) : (~x5 | x6);
  assign n849 = (~x4 | x5 | x6 | ~x7) & (x4 | ((x5 | ~x6 | x7) & (x6 | ~x7 | ~x2 | ~x5)));
  assign n850 = (~x7 & ~n851 & ~n854 & ~n855) | (x7 & n857);
  assign n851 = ~n281 & ((~n852 & n155) | n853);
  assign n852 = ~x2 ^ x3;
  assign n853 = ~x3 & x2 & x0 & ~x1;
  assign n854 = ~x1 & ((~x0 & x4 & ~x6) | (x0 & ~x2 & ~x4 & x6));
  assign n855 = n155 & ((n845 & n856) | (n141 & n825));
  assign n856 = x4 & ~x6;
  assign n857 = (~x6 | ~n209 | x3 | ~x4) & (x0 | ((~x4 | ~x6) & (x3 | x4 | x6 | ~n209)));
  assign z036 = ~n870 | n867 | n859 | n862;
  assign n859 = ~x2 & ((n155 & ~n861) | (~x1 & ~n860));
  assign n860 = (~x4 | ((x6 | ~x7 | x0 | x5) & (~x0 | ((x6 | x7) & (~x5 | ~x6 | ~x7))))) & (x0 | x4 | (x5 ? (~x6 ^ ~x7) : (~x6 | x7)));
  assign n861 = (~x4 | x5 | (~x6 ^ x7)) & (~x5 | ~x6 | ~x7);
  assign n862 = n864 & ((n863 & n865) | (~x3 & ~n866));
  assign n863 = ~x6 & ~x4 & ~x5;
  assign n864 = ~x1 & x7;
  assign n865 = x3 & ~x0 & ~x2;
  assign n866 = (~x0 | x2 | ~x4 | x5 | x6) & (~x2 | x4 | ((x5 | x6) & (x0 | ~x5 | ~x6)));
  assign n867 = ~x4 & ((x7 & ~n869) | (~n416 & ~n868));
  assign n868 = (~x0 | x1 | x2 | x3) & (x0 | ~x1 | ~x2 | ~x3);
  assign n869 = (~x0 | x1 | x2 | ~x3 | x5) & (x0 | ((x1 | ~x2 | ~x3) & (x3 | x5 | ~x1 | x2)));
  assign n870 = n873 & (~n203 | n872) & (n852 | n871);
  assign n871 = x0 ? (x1 | (x4 ? (x5 | ~x7) : (~x5 | x7))) : ((~x4 | ~x5 | x7) & (~x1 | ((~x5 | x7) & (x4 | x5 | ~x7))));
  assign n872 = (x1 | x4 | ~x5 | x6 | x7) & (~x4 | ~x7 | ((x5 | x6) & (~x1 | ~x5 | ~x6)));
  assign n873 = (~n874 | ~n876) & (x7 | ~n169 | n875);
  assign n874 = ~x3 & x2 & ~x0 & x1;
  assign n875 = x2 ? (~x3 | (~x1 & ~x5)) : (x3 | ~x5);
  assign n876 = ~x7 & x6 & x4 & ~x5;
  assign z037 = n878 | n884 | ~n888 | (~n405 & ~n887);
  assign n878 = ~x1 & (n880 | (n879 & n383 & n883));
  assign n879 = x4 & x5;
  assign n880 = ~x0 & ((x2 & ~n882) | (~n852 & ~n881));
  assign n881 = (~x4 | x5 | ~x6 | x7) & (x4 | ~x5 | x6 | ~x7);
  assign n882 = (~x3 | x5 | ~x6 | x7) & (~x4 | ~x5 | x6 | ~x7);
  assign n883 = x3 & x0 & ~x2;
  assign n884 = ~x0 & ((x3 & ~n885) | (n205 & ~n886));
  assign n885 = x1 ? ((x2 | x4 | x5 | ~x6) & (~x2 | ~x4 | ~x5 | x6)) : (~x4 | (~x5 ^ ~x6));
  assign n886 = (x2 | x4 | ~x5 | x6) & (~x4 | ((~x5 | ~x6) & (~x2 | x5 | x6)));
  assign n887 = (x1 | (x0 ? (~x4 | (~x2 ^ x3)) : (x4 | (~x2 & ~x3)))) & (x0 | ~x1 | x2 | x3 | x4);
  assign n888 = ~n889 & ~n893 & n895 & (n183 | n891);
  assign n889 = ~n537 & (~n890 | (x3 & n159 & n327));
  assign n890 = (~x0 | x1 | x2 | x5 | x6) & (x0 | ~x1 | ~x2 | ~x5 | ~x6);
  assign n891 = (~n231 | ~n351) & (~x4 | ~n401 | n892);
  assign n892 = x1 ? ~x5 : (x3 | x5);
  assign n893 = ~n894 & (x2 ? n825 : n856);
  assign n894 = (~x0 | x1 | x3 | ~x5) & (x0 | ~x1 | x5);
  assign n895 = ~n898 & (~n327 | ~n897) & (~n896 | ~n626);
  assign n896 = ~x7 & x6 & ~x4 & ~x5;
  assign n897 = ~x6 & ~x3 & x4;
  assign n898 = x6 & ~x4 & ~x2 & x0 & ~x1;
  assign z038 = ~n911 | n908 | n900 | n903;
  assign n900 = ~x3 & (x4 ? ~n902 : ~n901);
  assign n901 = (x0 | ~x1 | ((x2 | ~x5 | x7) & (x5 | ~x7))) & (x1 | ~x2 | ((~x5 | ~x7) & (~x0 | x5 | x7)));
  assign n902 = (~x0 | x1 | x2 | x5 | x7) & (x0 | ((~x5 | ~x7 | x1 | x2) & (~x1 | (x2 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n903 = ~x1 & (n904 | (n203 & ~n907));
  assign n904 = ~x2 & ((~x4 & ~n906) | (~n281 & ~n905));
  assign n905 = (x0 | x3 | x5 | x7) & (~x0 | ~x3 | ~x5 | ~x7);
  assign n906 = (~x0 | x3 | x5 | x6 | x7) & (x0 | ~x6 | (x3 ? (x5 | x7) : (~x5 | ~x7)));
  assign n907 = x5 ? ((~x3 | x4 | x6 | x7) & (~x6 | ((~x4 | ~x7) & (~x3 | (~x4 & ~x7))))) : (x6 | ~x7);
  assign n908 = ~n244 & (~n910 | (~x1 & ~n909));
  assign n909 = x0 ? ((x2 | ~x3 | x4 | ~x7) & (~x4 | x7 | ~x2 | x3)) : ((~x3 | ~x4 | x7) & (x2 | ((~x4 | x7) & (x3 | x4 | ~x7))));
  assign n910 = (~x0 | x1 | x2 | x3 | ~x7) & (x0 | ~x2 | (x1 ? (~x3 | ~x7) : (x3 | x7)));
  assign n911 = ~n912 & (~n155 | (n915 & (x4 | n914)));
  assign n912 = n293 & ~n913;
  assign n913 = (~x0 | x1 | x5 | x7) & (x0 | (x1 ? ((x5 | ~x7) & (~x4 | ~x5 | x7)) : (~x5 | ~x7)));
  assign n914 = (x2 | ~x3 | ~x5 | ~x6) & (~x2 | x7 | ((x5 | x6) & (x3 | ~x5 | ~x6)));
  assign n915 = (~n301 | ~n252) & (n437 | n916);
  assign n916 = x2 ? (~x3 | x7) : (x3 | ~x7);
  assign z039 = ~n932 | n929 | n926 | n918 | n923;
  assign n918 = ~x0 & (n921 | (~x2 & ~n919));
  assign n919 = (x1 | ~x3 | ~x4 | ~n694) & (x4 | n920);
  assign n920 = x1 ? ((~x5 | ~x6 | ~x7) & (x6 | x7 | x3 | x5)) : (x5 | ~x7 | (~x3 ^ x6));
  assign n921 = x2 & (x1 ? ~n922 : (n457 & n158));
  assign n922 = (x3 | x4 | ~x5 | ~x6 | ~x7) & (~x4 | x5 | x7 | (~x3 & x6));
  assign n923 = ~n183 & ((n231 & n924) | (~x0 & ~n925));
  assign n924 = ~x5 & ~x3 & x4;
  assign n925 = (~x1 | ((~x2 | x3) & (x2 | ~x3 | x4 | ~x5))) & (~x2 | x3 | x4 | ~x5) & (x1 | x2 | ~x4 | (~x3 & ~x5));
  assign n926 = ~n300 & ((n924 & n928) | (~x1 & ~n927));
  assign n927 = (~x0 | x2 | x3 | (x4 ^ ~x5)) & (~x3 | (~x0 ^ x2) | (~x4 ^ ~x5));
  assign n928 = ~x2 & ~x0 & x1;
  assign n929 = ~x1 & ((n338 & ~n931) | (~n223 & ~n930));
  assign n930 = (~x0 | x2 | ~x3 | x6) & (x0 | (x2 ? (~x3 | ~x6) : (x3 | x6)));
  assign n931 = (~x0 | x3 | x5 | ~x6) & (x0 | ~x3 | ~x5 | x6);
  assign n932 = n935 & (~n155 | n933) & (x0 | n934);
  assign n933 = (~x2 | ~x3 | ~x4 | ~x5 | ~x6) & (x2 | x6 | (x3 ? (x4 | x5) : ~x5));
  assign n934 = (x1 | ~x2 | x3 | ~x4 | ~x6) & (~x1 | ~x3 | (x2 ? (x4 | ~x6) : (~x4 | x6)));
  assign n935 = (~n365 | ~n716) & (~n567 | ~n231);
  assign z040 = n946 | n950 | (x2 ? ~n937 : ~n942);
  assign n937 = x0 ? (~n205 | ~n938) : n939;
  assign n938 = x7 & x6 & ~x4 & x5;
  assign n939 = (x5 | n941) & (x4 | ~x5 | n183 | ~n940);
  assign n940 = x1 & ~x3;
  assign n941 = (~x1 | x3 | ~x4 | x6 | x7) & (~x6 | (x1 ? (x3 ? (x4 | x7) : (~x4 | ~x7)) : (x3 ? (~x4 | ~x7) : (x4 ^ ~x7))));
  assign n942 = x0 ? (x1 | n943) : (x1 ? n945 : n944);
  assign n943 = (x3 | ~x4 | x6 | (x5 ^ ~x7)) & (~x6 | ((~x3 | x4 | ~x5 | x7) & (x3 | (x4 ? (x5 ^ x7) : (x5 | ~x7)))));
  assign n944 = (x3 | x4 | ~x5 | ~x6 | x7) & (~x3 | ((~x6 | ~x7 | x4 | ~x5) & ((x4 ^ x5) | (x6 ^ ~x7))));
  assign n945 = (~x5 | ((~x6 | (x3 ? (~x4 | ~x7) : (x4 ^ ~x7))) & (x3 | x4 | x6 | x7))) & (x3 | x4 | x5 | (x6 ^ ~x7));
  assign n946 = ~x7 & (n948 | ~n949 | (~x1 & ~n947));
  assign n947 = (x5 | ((x0 | x2 | x3 | ~x4) & ((~x0 ^ x2) | (x3 ^ x4)))) & (x0 | ~x5 | ((~x3 | x4) & (~x2 | x3 | ~x4)));
  assign n948 = x3 & n155 & (x2 ? x5 : (~x4 & ~x5));
  assign n949 = (~x0 | x1 | ~x2 | x3 | x4) & (x0 | ~x1 | x2 | ~x3 | ~x4);
  assign n950 = x7 & (~n951 | (~n273 & ~n664));
  assign n951 = (n952 | n953) & (x0 | n954);
  assign n952 = x0 ? (x1 | x3) : (~x1 | ~x3);
  assign n953 = x2 ? (~x4 | x5) : (x4 | ~x5);
  assign n954 = (x1 | ((~x2 | x3 | x4 | ~x5) & (~x4 | x5 | x2 | ~x3))) & (~x1 | x2 | x3 | ~x4 | x5);
  assign z041 = n956 | n961 | ~n967 | (n268 & ~n959);
  assign n956 = ~x1 & ((n391 & ~n958) | (~x0 & ~n957));
  assign n957 = (x3 | (~x4 & ~x6) | (~x2 ^ ~x5)) & (x2 | ~x3 | x6 | (x4 ^ x5));
  assign n958 = x3 ? (x5 | ~x6) : (~x4 | x6);
  assign n959 = (x3 | n960) & (x2 | ~x3 | ~x5 | ~n675);
  assign n960 = (x2 | ~x4 | x5 | ~x6 | ~x7) & (x7 | ((~x2 | ~x5 | (~x4 ^ x6)) & (x2 | x4 | x5 | ~x6)));
  assign n961 = ~x0 & (~n963 | (~x4 & ~x7 & ~n962));
  assign n962 = (~x2 | x5 | (x1 ? (~x3 | x6) : (x3 | ~x6))) & (x1 | x2 | ~x5 | (x3 ^ x6));
  assign n963 = (~n716 | ~n966) & (n537 | n964 | n965);
  assign n964 = x3 ^ x6;
  assign n965 = x1 ? (x2 | ~x5) : (~x2 | x5);
  assign n966 = ~x3 & ~x1 & ~x2;
  assign n967 = ~n969 & (~n155 | n968) & (n837 | n970);
  assign n968 = x2 ? (x4 | (x3 ? (~x5 | ~x6) : (x5 ^ ~x6))) : ((~x3 | (x4 ? (~x5 | x6) : x5)) & (x5 | ((x3 | ~x4 | ~x6) & (x4 | x6))));
  assign n969 = ~n374 & (n853 | (n279 & (~x1 ^ x2)));
  assign n970 = (x0 | ~x1 | ~x2 | x3 | ~x4) & (x1 | ((~x3 | ~x4 | x0 | ~x2) & (~x0 | x2 | (~x3 ^ ~x4))));
  assign z042 = ~n980 | (~x1 & ~n972) | (~x0 & x1 & ~n977);
  assign n972 = n975 & (~n585 | n973) & (n964 | n974);
  assign n973 = (x2 | (x3 ? (~x4 | ~x5) : (x4 | ~x6))) & (~x5 | ~x6 | x3 | x4) & (~x3 | x5 | x6 | (~x2 & x4));
  assign n974 = x0 ? (x2 | ((x5 | ~x7) & (~x4 | (x5 & ~x7)))) : (~x2 | x4 | (~x5 & x7));
  assign n975 = (n419 | n976) & (~n243 | ~n883);
  assign n976 = (~x0 | x2 | ~x3 | x4) & (x0 | ~x2 | x3 | ~x4);
  assign n977 = ~n978 & ~n979 & (~n694 | (~n141 & ~n249));
  assign n978 = x3 & ((n538 & n675) | (n338 & n694));
  assign n979 = ~x3 & (x2 ? (x5 & x7) : (~x5 & (x6 ^ ~x7)));
  assign n980 = ~n981 & (n413 | n983);
  assign n981 = ~n416 & ((n155 & ~n964) | (~x1 & ~n982));
  assign n982 = ((x0 ? (~x2 | x3) : (x2 | ~x3)) | (x4 ^ ~x6)) & (~x0 | x2 | ~x3 | x4 | x6) & (x0 | x3 | ((~x4 | ~x6) & (x2 | x4 | x6)));
  assign n983 = (x1 | (x0 ? (x3 | x4) : (~x4 | (x2 ^ x3)))) & (x0 | x2 | ~x3 | (~x1 & x4));
  assign z043 = n985 | ~n994 | ~n1000 | (~x3 & ~n991);
  assign n985 = ~x0 & (n989 | (~x1 & (n986 | n988)));
  assign n986 = x7 & ~n987;
  assign n987 = (~x2 | x3 | x4 | ~x5 | x6) & ((~x2 ^ ~x6) | (x3 ? (~x4 | ~x5) : (x4 | x5)));
  assign n988 = n334 & ((x2 & x3 & x4 & ~x6) | (~x2 & x6 & (x3 ^ x4)));
  assign n989 = n990 & n215 & (x3 ? (x6 & ~x7) : (~x6 ^ x7));
  assign n990 = ~x4 & x5;
  assign n991 = n993 & (~n534 | ~n928) & (x1 | n992);
  assign n992 = (x0 | x2 | ~x4 | x5 | ~x7) & ((~x0 ^ x5) | (x2 ? (~x4 | ~x7) : (x4 | x7)));
  assign n993 = (~x0 | x1 | x2 | ~x5 | ~x7) & (x0 | ~x2 | x5 | (~x1 ^ ~x7));
  assign n994 = ~n998 & (n996 | ~n997) & (n995 | n999);
  assign n995 = x3 ? (~x6 | ~x7) : (x6 | x7);
  assign n996 = (~x2 | x3 | ~x4 | x6 | x7) & (x2 | (~x3 ^ x4) | (x6 ^ ~x7));
  assign n997 = ~x5 & x0 & ~x1;
  assign n998 = ~n416 & ((n155 & n828) | (n268 & (n828 | n464)));
  assign n999 = (~x0 | x1 | x2 | ~x5) & (x0 | ~x1 | ~x2 | x5);
  assign n1000 = (~x3 | n1001) & (x0 | (~n1003 & ~n1004));
  assign n1001 = (x4 | n1002) & (~x2 | ~x4 | ~n155 | n283);
  assign n1002 = (~x0 | x1 | x2 | ~x5 | x7) & (x0 | ((~x2 | ~x5 | ~x7) & (~x1 | x5 | (x2 ^ ~x7))));
  assign n1003 = n940 & (x2 ? (x5 & ~n183) : (~x5 & n383));
  assign n1004 = ~x5 & n201 & (x2 ? (x6 & ~x7) : (~x6 ^ x7));
  assign z044 = ~n1015 | (~x1 & (~n1006 | ~n1011));
  assign n1006 = ~n1008 & n1009 & (~x3 | n1007);
  assign n1007 = (x0 | ~x2 | x4 | ~x5 | ~x6) & (~x4 | ((x2 | (x0 ? (x5 ^ ~x6) : (x5 | x6))) & (x0 | ~x2 | ~x5 | x6)));
  assign n1008 = x0 & ~x4 & (x2 ? (~x3 & x6) : (x3 & ~x6));
  assign n1009 = ~n1010 & (x0 | ~n845 | ~n631);
  assign n1010 = x6 & ~x3 & ~x0 & x2 & x4;
  assign n1011 = ~n1012 & (~n293 | n723);
  assign n1012 = ~x3 & (x6 ? ~n1014 : ~n1013);
  assign n1013 = ((x0 ^ x2) | (x4 ? (~x5 | x7) : (x5 | ~x7))) & (~x7 | ((~x0 | x2 | ~x4 | x5) & (x0 | ~x2 | x4 | ~x5)));
  assign n1014 = (x5 | ((x0 | ((x2 | ~x4 | ~x7) & (x4 | x7))) & (~x0 | x2 | x4 | ~x7))) & (x0 | ~x2 | x4 | x7);
  assign n1015 = ~n1016 & (~n155 | (~n1019 & n1020));
  assign n1016 = ~n300 & ((n1017 & n928) | (~x1 & ~n1018));
  assign n1017 = x5 & x3 & ~x4;
  assign n1018 = x0 ? (x3 | (x5 ? x2 : ~x4)) : (~x3 | x5 | (~x2 & x4));
  assign n1019 = ~x5 & ~x7 & (x2 ? (~x3 ^ x6) : (~x3 & x6));
  assign n1020 = n1022 & (~n598 | n1021) & (~n845 | ~n559);
  assign n1021 = (~x2 | x4 | x5 | x6) & (x2 | ~x4 | ~x5 | ~x6);
  assign n1022 = (x2 | x3 | ~x4 | ~x5 | ~x6) & ((~x3 ^ ~x6) | (~x2 ^ ~x5));
  assign z045 = n1024 | n1029 | n1033 | (n155 & ~n1032);
  assign n1024 = ~x3 & (n1025 | (n155 & ~n1028));
  assign n1025 = ~x1 & ((x4 & ~n1026) | (n382 & ~n1027));
  assign n1026 = (x0 | x2 | ~x6 | (x5 ^ x7)) & (x6 | (x0 ? (x2 ? (~x5 | x7) : (x5 | ~x7)) : (x2 ? (x5 ^ x7) : (~x5 | x7))));
  assign n1027 = (~x0 | ~x7 | (x2 ^ x6)) & (x7 | ((x2 | ~x6) & (x0 | ~x2 | x6)));
  assign n1028 = ((~x2 ^ ~x7) | ((x5 | ~x6) & (x4 | ~x5 | x6))) & (~x2 | x5 | x6 | x7) & (x2 | ~x7 | ((~x5 | ~x6) & (~x4 | x5 | x6)));
  assign n1029 = ~x1 & (x5 ? ~n1031 : ~n1030);
  assign n1030 = ((x0 ^ ~x7) | (x2 ? x3 : (~x3 | ~x4))) & (~x3 | ((x0 | ~x2 | x7) & (~x0 | x2 | x4 | ~x7)));
  assign n1031 = (x3 | (x0 ? (x2 ? (x4 | ~x7) : x7) : (x4 | (x2 ^ ~x7)))) & (x0 | ~x3 | ~x4 | (~x2 ^ ~x7));
  assign n1032 = (~x5 | (x2 ? (~x7 | (~x3 & ~x4)) : (x7 | (~x3 ^ x4)))) & (~x3 | x5 | (x2 ? (x4 | x7) : ~x7));
  assign n1033 = x3 & (~n1037 | (x5 & (n1034 | n1036)));
  assign n1034 = n1035 & (x0 ? (~x1 & ~x7) : ((~x4 & x7) | (x1 & x4 & ~x7)));
  assign n1035 = ~x2 & x6;
  assign n1036 = n203 & n285 & (x1 ^ x7);
  assign n1037 = (n244 | n1038) & (~n146 | ~n383 | n220);
  assign n1038 = (~x0 | x1 | x2 | ~x4 | ~x7) & (x0 | x7 | (x1 ? (~x2 | ~x4) : (x2 | x4)));
  assign z046 = n1040 | n1044 | n1058 | (~x1 & ~n1049);
  assign n1040 = x6 & ~n1041;
  assign n1041 = n1043 & (x0 ? (~n209 | ~n351) : n1042);
  assign n1042 = (~x4 | ((x1 | x3 | (x2 ^ ~x5)) & (~x1 | ~x2 | ~x3 | ~x5))) & (x2 | ~x3 | x4 | (x1 & ~x5));
  assign n1043 = (~x0 | x1 | x2 | ~x3 | ~x5) & (x0 | ~x1 | x3 | x5);
  assign n1044 = ~x6 & (~n1046 | (~x1 & ~n1045));
  assign n1045 = x0 ? (x2 | x5 | (~x3 ^ x4)) : (x3 ? (~x4 | (~x2 & ~x5)) : (x4 | ~x5));
  assign n1046 = (~n155 | ~n1047) & (n223 | n1048);
  assign n1047 = ~x5 & x3 & ~x4;
  assign n1048 = (~x0 | x1 | ~x2 | x3) & (x0 | ~x1 | x2 | ~x3);
  assign n1049 = x6 ? (~n1053 & n1054) : (~n1050 & n1051);
  assign n1050 = n146 & (x4 ? (x7 & n845) : (~x7 & n141));
  assign n1051 = ~n1052 & (~n391 | ~n402) & (~n171 | ~n883);
  assign n1052 = ~x0 & ~x5 & (x2 ? (~x3 & x7) : (x3 & ~x7));
  assign n1053 = n795 & (((x2 ^ x4) & (x0 ^ ~x7)) | (x0 & x2 & x4 & ~x7));
  assign n1054 = (n1055 | n1057) & (x0 | ~n1056);
  assign n1055 = x4 ^ x7;
  assign n1056 = x2 & x3 & x5 & (~x4 ^ ~x7);
  assign n1057 = (~x0 | x2 | ~x3 | x5) & (x0 | ~x2 | x3 | ~x5);
  assign n1058 = n155 & (x5 ? ~n1060 : ~n1059);
  assign n1059 = (x2 | x3 | x4 | x6 | ~x7) & (~x2 | ~x3 | ~x4 | ~x6 | x7);
  assign n1060 = x6 ? (((x3 ^ ~x7) | (x2 ^ ~x4)) & (x2 | x3 | x4 | x7)) : ((~x3 | ~x4 | ~x7) & (~x2 | (~x3 ^ ~x7)));
  assign z047 = n1067 | ~n1072 | (x6 ? ~n1062 : ~n1069);
  assign n1062 = (x3 | n1063) & (x0 | ~x3 | n1066);
  assign n1063 = (x1 | n1064) & (x0 | ~x1 | n283 | n1065);
  assign n1064 = (~x4 | ((x0 | ~x2 | x5 | x7) & (~x0 | (x2 ? (x5 | ~x7) : (~x5 | x7))))) & (x0 | ~x5 | (x2 ? ~x7 : (x4 | x7)));
  assign n1065 = x2 & x4;
  assign n1066 = ((~x1 ^ x2) | (~x5 ^ ~x7)) & (~x2 | ~x7 | ((x4 | ~x5) & (~x1 | ~x4 | x5)));
  assign n1067 = ~n416 & ((n567 & n928) | (~x1 & ~n1068));
  assign n1068 = x0 ? (~x6 | (x2 ? (x3 | x4) : ~x3)) : ((x3 | x6) & (x2 | (x6 & (x3 | ~x4))));
  assign n1069 = x5 ? (~x7 | n1070) : ((~n201 | n1071) & (x7 | n1070));
  assign n1070 = x0 ? (x1 | x2 | (x3 & x4)) : (~x1 | (~x2 & (~x3 | ~x4)));
  assign n1071 = (~x0 | x2 | ~x4 | x7) & (x0 | ~x2 | x4 | ~x7);
  assign n1072 = (n848 | ~n1073) & (x1 | n335 | n769);
  assign n1073 = ~x0 & x1 & (x3 ^ x4);
  assign z048 = n1079 | ~n1082 | (~x0 & ~n1075) | ~n1086;
  assign n1075 = ~n1078 & (x4 | (~x1 & n1077) | (x1 & n1076));
  assign n1076 = (~x2 | ~x3 | ~x5 | ~x6 | ~x7) & (x2 | x3 | x5 | x6 | x7);
  assign n1077 = (~x5 | ((~x2 | x3 | x6 | x7) & (x2 | ~x7 | (~x3 ^ x6)))) & (~x2 | x5 | (x3 ? x6 : (~x6 | x7)));
  assign n1078 = n141 & n879 & (x1 ? (x6 ^ x7) : (~x6 & ~x7));
  assign n1079 = ~n300 & (n1081 | (~x1 & ~n1080));
  assign n1080 = (~x0 | x2 | ~x3 | ~x4 | ~x5) & (~x2 | (x0 ? (x3 | (x4 & x5)) : (~x3 | (x4 ^ ~x5))));
  assign n1081 = ~x2 & n155 & (x4 ? ~x3 : (x3 | n990));
  assign n1082 = n1085 & (x0 | (n1083 & (x4 | n1084)));
  assign n1083 = (x1 | ~x2 | x3 | ~x4 | x6) & (~x6 | ((~x1 | (x2 ? (x3 | x4) : (~x3 | ~x4))) & (x1 | x2 | x3 | ~x4)));
  assign n1084 = (x1 | ((~x2 | x3 | x6 | ~x7) & (~x6 | x7 | x2 | ~x3))) & (~x1 | x2 | x3 | x6 | ~x7);
  assign n1085 = x6 | ~n157 | (x3 ? x4 : (~x4 | ~x7));
  assign n1086 = (n183 | n1087) & (~x4 | ~n268 | n1088);
  assign n1087 = (x3 | x4 | x1 | x2) & (x0 | ((~x3 | ~x4 | x1 | x2) & (~x1 | ~x2 | (x3 ^ ~x4))));
  assign n1088 = (x6 | x7 | x3 | ~x5) & (x2 | x5 | (x3 ? x6 : (~x6 | x7)));
  assign z049 = n1094 | ~n1097 | (~x1 & ~n1090);
  assign n1090 = x3 ? (x0 | n1093) : (~n1091 & ~n1092);
  assign n1091 = n692 & (x2 ? (x5 & n191) : (~x5 & n266));
  assign n1092 = x6 & n312 & (x2 ? (~x5 & x7) : (~x5 ^ x7));
  assign n1093 = x2 ? (~x4 | ~x5 | (~x6 ^ ~x7)) : (x4 | x5 | (x6 ^ ~x7));
  assign n1094 = ~x3 & ((n1095 & n928) | (~x1 & ~n1096));
  assign n1095 = x7 & ~x4 & ~x5;
  assign n1096 = x0 ? (~x4 | ((x5 | x7) & (x2 | ~x5 | ~x7))) : (x4 | (x2 ? (~x5 ^ ~x7) : (~x5 | x7)));
  assign n1097 = ~n1101 & n1103 & (~x3 | (~n1098 & ~n1099));
  assign n1098 = ~n416 & ((~x0 & x2 & (~x1 ^ x4)) | (x0 & ~x1 & ~x2 & x4));
  assign n1099 = n1100 & (x1 ? (x2 & n382) : ~n953);
  assign n1100 = ~x0 & ~x7;
  assign n1101 = n990 & n155 & ~n1102;
  assign n1102 = (x2 | x3 | (~x6 ^ x7)) & (~x3 | ((~x6 | ~x7) & (~x2 | x6 | x7)));
  assign n1103 = (~x0 | x1 | x4 | n1104) & (x0 | (n1105 & (~x1 | ~x4 | n1104)));
  assign n1104 = (x3 | x7) & (x2 | ~x3 | ~x7);
  assign n1105 = x1 ? (x4 | (x2 ? (x3 | ~x7) : (~x3 | x7))) : (~x4 | ((x2 | ~x3 | x7) & (x3 | ~x7)));
  assign z050 = ~n1118 | (~x0 & (~n1107 | ~n1114));
  assign n1107 = ~n1110 & (x2 | (n1108 & n1109)) & n1111;
  assign n1108 = (x1 | ~x3 | x4 | ~x5 | ~x6) & (~x1 | x6 | (x3 ? (x4 | ~x5) : (~x4 | x5)));
  assign n1109 = x3 ? ((x5 & x6) | (x1 & (x5 | x6))) : (~x1 | (~x5 & ~x6));
  assign n1110 = x1 & x3 & (x2 ? (x4 & ~x6) : (~x4 & x6));
  assign n1111 = ~n1113 & (n204 | n1112) & (x1 | ~n249);
  assign n1112 = x1 ? (x2 | x5) : (~x2 | ~x5);
  assign n1113 = x6 & x1 & x2 & x3 & x5;
  assign n1114 = (x2 | ~x5 | n1117) & (~n1115 | ~n1116);
  assign n1115 = ~x3 & ~x1 & x2;
  assign n1116 = x7 & x6 & ~x4 & ~x5;
  assign n1117 = (~x1 | ~x3 | ~x4 | x6 | x7) & (x1 | ~x6 | (x3 ? (~x4 | x7) : (x4 | ~x7)));
  assign n1118 = ~n268 | x2 | (x3 & ~n139 & ~n1047);
  assign z051 = n1124 | ~n1127 | (x5 & ~n1120);
  assign n1120 = (x1 | n1122) & (x0 | ~x1 | ~x4 | ~n1121);
  assign n1121 = ~x6 & (x2 ? (~x3 & ~x7) : (x3 & x7));
  assign n1122 = (x2 | n1123) & (x0 | ~x2 | x7 | n643);
  assign n1123 = (x0 | ~x3 | ~x4 | ~x6 | ~x7) & (x4 | ((x0 | x3 | ~x6 | ~x7) & (~x0 | x6 | (~x3 ^ ~x7))));
  assign n1124 = ~x0 & (x1 ? ~n1126 : ~n1125);
  assign n1125 = (x4 | (x2 ? (x3 | (~x5 ^ ~x6)) : (~x3 | (x5 ^ ~x6)))) & (~x2 | ~x4 | ~x5 | (~x3 ^ ~x6));
  assign n1126 = (~x2 | ~x3 | ~x4 | x5 | x6) & (~x5 | (~x3 ^ ~x6) | (x2 ^ ~x4));
  assign n1127 = ~n1130 & ~n1131 & (x2 ? n1128 : n1129);
  assign n1128 = (~x0 | x1 | x3 | x4 | x5) & (x0 | ((x3 | ~x4 | x5) & (~x1 | (x3 ? (~x4 | ~x5) : x5))));
  assign n1129 = (x1 | (x0 ? (x3 ? ~x4 : (x4 | x5)) : (x3 | ~x4))) & (x0 | x3 | (x4 ? x5 : ~x1));
  assign n1130 = n157 & n773 & n247;
  assign n1131 = n1132 & n205 & ~n1133;
  assign n1132 = ~x5 & x6;
  assign n1133 = (~x0 | x2 | ~x4 | ~x7) & (x0 | ~x2 | x4 | x7);
  assign z052 = n1135 | n1142 | n1144 | (n159 & ~n1149);
  assign n1135 = ~x1 & (n1140 | (~x2 & (n1136 | ~n1137)));
  assign n1136 = ~n283 & ((x0 & ~x3 & ~x4 & ~x6) | (~x0 & x3 & x4 & x6));
  assign n1137 = (n1138 | n1139) & (x0 | ~n158 | ~n339);
  assign n1138 = x4 ? (x5 | x7) : (~x5 | ~x7);
  assign n1139 = x0 ? (~x3 | x6) : (x3 | ~x6);
  assign n1140 = x2 & (x0 ? (n176 & n693) : ~n1141);
  assign n1141 = (x4 | ((x5 | ~x6 | x7) & (x6 | ~x7 | ~x3 | ~x5))) & (x3 | ~x4 | ~x5 | ~x6 | ~x7);
  assign n1142 = n155 & (x6 ? (n338 & ~n250) : ~n1143);
  assign n1143 = x2 ? ((~x5 | ~x7 | x3 | ~x4) & (x5 | x7 | ~x3 | x4)) : (~x4 | ((x5 | x7) & (~x3 | ~x5 | ~x7)));
  assign n1144 = x5 & ((x6 & ~n1145) | n1146 | ~n1147);
  assign n1145 = (~x3 | x4 | x1 | x2) & (x0 | ((~x3 | ~x4 | x1 | ~x2) & (~x1 | x3 | (x2 & ~x4))));
  assign n1146 = ~x1 & ((x0 & ~x2 & x4) | (~x4 & x6 & ~x0 & x2));
  assign n1147 = (~x6 | n1148) & (~x2 | (n1148 & (x4 | ~x6 | ~n155)));
  assign n1148 = (~x0 | x1 | x3 | x4) & (x0 | ~x1 | ~x3 | ~x4);
  assign n1149 = (x2 & (x0 | (x1 & x3 & ~x4))) | (x0 & (x3 | ~x4)) | (~x3 & ~x4 & ~x1 & ~x2) | (x1 & x4 & (~x2 | ~x3));
  assign z053 = n1151 | n1159 | ~n1161 | (~x3 & ~n1156);
  assign n1151 = ~x2 & (n1152 | (n155 & ~n1155));
  assign n1152 = ~x1 & ((x6 & ~n1153) | (n191 & ~n1154));
  assign n1153 = (x3 | ((x4 | ~x5 | ~x7) & (x5 | x7 | ~x0 | ~x4))) & (~x7 | ((~x3 | ~x4 | x5) & (x0 | ((~x4 | x5) & (~x3 | (~x4 & x5))))));
  assign n1154 = (x0 | ~x4 | x5) & (~x3 | (x4 ^ x5));
  assign n1155 = (~x6 | ~x7 | (x3 ? (~x4 | ~x5) : x5)) & (x4 | x7 | ((~x5 | x6) & (x3 | (~x5 & x6))));
  assign n1156 = (x1 | x6 | n1157) & (x0 | (n1158 & (~x1 | ~x6 | n1157)));
  assign n1157 = x2 ? (x4 | x5) : (~x4 | ~x5);
  assign n1158 = (~x5 | ~x6 | ~x2 | x4) & (x5 | ((~x1 | ~x2 | ~x4 | x6) & (x1 | ~x6 | (x2 ^ x4))));
  assign n1159 = n279 & ~n1160;
  assign n1160 = (~x1 | ~x2 | ~x4 | ~x5 | x6) & (~x6 | ((x1 | ~x2 | ~x4) & (x4 | (x1 ? (x2 ^ x5) : (x2 | ~x5)))));
  assign n1161 = ~n1162 & (~x2 | (~n1167 & (x0 | n1165)));
  assign n1162 = ~n183 & ((n268 & ~n1164) | (~x0 & ~n1163));
  assign n1163 = (~x3 | (x1 ? (x2 ? (x4 | x5) : ~x4) : (x4 | (~x2 ^ ~x5)))) & (~x1 | ~x4 | (x2 ? (x3 | ~x5) : x5));
  assign n1164 = (x2 & (x3 | (~x4 & ~x5))) | (x4 & (x5 | (~x2 & ~x3)));
  assign n1165 = x1 ? (~n448 | ~n773) : (n300 | n1166);
  assign n1166 = x3 ? (x4 | x5) : (~x4 | ~x5);
  assign n1167 = n139 & n472;
  assign z054 = n1174 | n1177 | ~n1179 | (x7 & ~n1169);
  assign n1169 = ~n1170 & (n336 | n1173) & (~n226 | ~n702);
  assign n1170 = ~x4 & ((n1171 & n327) | (~x5 & ~n1172));
  assign n1171 = x6 & ~x3 & x5;
  assign n1172 = (~x0 | x1 | x2 | ~x3 | ~x6) & (x0 | ((~x1 | ~x3 | (x2 ^ ~x6)) & (x1 | ~x2 | x3 | ~x6)));
  assign n1173 = (~x0 | x1 | x3 | x4 | ~x5) & (x0 | ~x1 | ~x4 | (x3 ^ x5));
  assign n1174 = n1175 & ((n170 & n276) | (~x2 & ~n1176));
  assign n1175 = ~x1 & ~x7;
  assign n1176 = (~x0 | ~x3 | ~x4 | ~x6) & (x4 | (x0 ? (x3 ? (x5 | x6) : (~x5 | ~x6)) : (x3 | (x5 ^ ~x6))));
  assign n1177 = ~x4 & ((~n295 & ~n427) | (~x0 & ~n1178));
  assign n1178 = (~x1 | x2 | ~x3 | ~x5 | ~x7) & (x1 | x3 | (x2 ? (x5 | x7) : (~x5 | ~x7)));
  assign n1179 = n1182 & (n1055 | n1180) & (x0 | n1181);
  assign n1180 = (x1 | ((x0 | x2 | ~x3) & (x3 | x5 | ~x0 | ~x2))) & (x0 | (x2 ? (x3 | ~x5) : (~x3 | x5)));
  assign n1181 = (~x1 | x2 | x3 | x4 | ~x7) & (~x2 | ~x3 | ((~x4 | x7) & (x1 | x4 | ~x7)));
  assign n1182 = (~n157 | ~n1183) & (~x4 | ~n238 | n1184);
  assign n1183 = ~x7 & ~x3 & x4;
  assign n1184 = x2 ? (x5 | x7) : ((~x5 | x7) & (x1 | x5 | ~x7));
  assign z055 = n1186 | n1191 | ~n1195 | (~n273 & ~n1194);
  assign n1186 = ~x3 & (n1187 | (n312 & ~n1190));
  assign n1187 = x4 & ((n585 & ~n1189) | (~x7 & ~n1188));
  assign n1188 = (x0 | ~x1 | x5 | ~x6) & (~x0 | x1 | (x2 ? (~x5 | x6) : (x5 | ~x6)));
  assign n1189 = (x1 | x2 | x5 | x6) & (~x1 | ~x5 | ~x6);
  assign n1190 = (x1 | x2 | x6 | (x5 ^ ~x7)) & (~x6 | ((~x2 | x5 | ~x7) & (~x1 | ((x5 | ~x7) & (~x2 | ~x5 | x7)))));
  assign n1191 = ~x1 & (x6 ? ~n1192 : (n653 & ~n1193));
  assign n1192 = x0 ? ((~x2 | x3 | x5) & (x2 | ~x3 | x4 | ~x5)) : (x2 | (x3 ? (~x4 | ~x5) : (x4 | x5)));
  assign n1193 = x0 ? (x2 | ~x3) : (~x2 | x3);
  assign n1194 = (~x0 | x1 | x2 | x3 | ~x6) & (~x3 | ((x1 | x2 | x6) & (x0 | (x6 & (x1 | ~x2)))));
  assign n1195 = ~n1197 & n1199 & (x0 | n1196);
  assign n1196 = (x1 | ~x3 | x4 | ~x5) & (x3 | ((x5 | ~x6 | x1 | ~x4) & (~x1 | x6 | (~x4 ^ x5))));
  assign n1197 = x3 & x6 & n155 & ~n1198;
  assign n1198 = x4 ? (~x5 ^ x7) : ((x5 | x7) & (~x2 | ~x5 | ~x7));
  assign n1199 = (~n327 | ~n1200) & (~n276 | ~n472);
  assign n1200 = ~x6 & x3 & x4 & ~x5;
  assign z056 = ~n1207 | (~x3 & (n1203 | (n1202 & ~n1206)));
  assign n1202 = ~x0 & x6;
  assign n1203 = ~x6 & ((n707 & ~n1205) | (~x1 & ~n1204));
  assign n1204 = x0 ? ((x2 | x4 | x5 | ~x7) & (~x2 | ~x4 | ~x5 | x7)) : (x2 | x7 | (~x4 ^ x5));
  assign n1205 = ~x5 & ~x2 & x4;
  assign n1206 = (~x1 | x7 | (~x2 & ~x4 & x5)) & (x1 | x2 | x4 | ~x7);
  assign n1207 = ~n1208 & ~n1213 & (x0 | (~n1210 & ~n1212));
  assign n1208 = n279 & (x1 ? ~n1209 : (n448 & n338));
  assign n1209 = x7 ? (x6 | (x2 & x4 & ~x5)) : ~x6;
  assign n1210 = x1 & ((n141 & n1211) | (n845 & n631));
  assign n1211 = ~x6 & x4 & ~x5;
  assign n1212 = n357 & (x2 | n151 | (n990 & n293));
  assign n1213 = n310 & ((~x2 & (x3 | x4)) | (~x3 & (~n953 | (x2 & ~x4))));
  assign z057 = ~n1221 | (~x0 & (~n1215 | (x5 & ~n1220)));
  assign n1215 = x5 ? (~n1216 | n1219) : (~n1217 & ~n1218);
  assign n1216 = x1 & ~x4;
  assign n1217 = ~n183 & ((~x1 & ~x2 & x3 & ~x4) | (x1 & x4 & (~x2 ^ x3)));
  assign n1218 = n845 & ((~x1 & x4 & ~n300) | (~x4 & n787));
  assign n1219 = (~x2 | ~x3 | ~x6 | ~x7) & (x2 | x3 | (x6 ^ x7));
  assign n1220 = (x1 | x2 | x4 | (x3 ^ x7)) & (~x4 | ((x1 | x2 | x3 | ~x7) & (~x1 | x7 | (x2 ^ x3))));
  assign n1221 = n1222 & ~n1224 & (~n365 | ~n717) & n1225;
  assign n1222 = ~n231 | ((~n176 | ~n228) & ~n1223);
  assign n1223 = x7 & ~x3 & ~x4;
  assign n1224 = n279 & ((x1 & x2 & ~x4 & ~x7) | (~x1 & ~x2 & x4 & x7));
  assign n1225 = (~x0 | x1 | x2 | ~x7) & (x0 | (x1 ? (x7 | (~x2 ^ x3)) : (~x2 | ~x7)));
  assign z058 = n1227 | n1231 | ~n1236 | (~x1 & ~n1230);
  assign n1227 = ~x0 & ((x1 & ~n1228) | (n510 & ~n1229));
  assign n1228 = (x3 | (x2 ? (x5 | ~x6) : (x4 ? (x5 | x6) : (~x5 | ~x6)))) & (~x2 | ((~x4 | x5 | ~x6) & (~x5 | x6 | ~x3 | x4)));
  assign n1229 = (~x2 | x3 | ~x4 | ~x6) & (x2 | ((x4 | ~x6) & (x3 | ~x4 | x6)));
  assign n1230 = x2 ? (x0 ? (x3 | (x4 ^ ~x5)) : (~x3 & (~x4 | ~x5))) : ((~x4 | x5 | ~x0 | ~x3) & (x4 | ~x5 | x0 | x3));
  assign n1231 = ~x4 & (x6 ? ~n1232 : (n795 & ~n1235));
  assign n1232 = (~n1233 | n1234) & (~x3 | ~n157 | ~n590);
  assign n1233 = ~x7 & ~x0 & x2;
  assign n1234 = x1 ? (~x3 | ~x5) : (x3 | x5);
  assign n1235 = (x0 & (x1 | (~x2 & x7))) | (x1 & ~x2 & x7) | (~x7 & (x2 | (~x0 & ~x1)));
  assign n1236 = n1238 & (~x2 | ~n155 | n1237);
  assign n1237 = (x3 & ~x4 & x5) | (~x5 & (~x3 | x4));
  assign n1238 = (~n243 | ~n853) & (~n158 | ~n1132 | ~n231);
  assign z059 = (x3 | ~n1240) & (~x3 | n1248 | n1250 | ~n1251);
  assign n1240 = ~n1243 & ~n1247 & (x1 | (n1241 & n1246));
  assign n1241 = (~n693 | ~n722) & (~x0 | n1242);
  assign n1242 = (~x6 | ~x7 | x4 | ~x5) & (x7 | (x4 ? (x2 ? (~x5 | x6) : (x5 | ~x6)) : (x5 | x6)));
  assign n1243 = n1245 & ((n191 & n1244) | (x2 & ~n419));
  assign n1244 = ~x2 & ~x5;
  assign n1245 = ~x4 & ~x0 & x1;
  assign n1246 = (x0 | x4 | ~x5) & (~x4 | x5 | ((~x0 | ~x2) & x6));
  assign n1247 = n155 & ((n159 & n301) | (~x2 & ~n437));
  assign n1248 = ~x4 & ((n140 & n339) | (~n1249 & ~n839));
  assign n1249 = x5 ? (~x6 | x7) : (x6 | ~x7);
  assign n1250 = ~x0 & ((x4 & ~x5 & x6) | (x5 & ~x6 & x1 & ~x4));
  assign n1251 = (~x4 & (x6 ? x5 : ~n157)) | (x0 & ~n157) | (~x5 & (x4 | ~x6));
  assign z060 = ~n1260 | n1253 | n1257;
  assign n1253 = x5 & (n1254 | (n191 & n176 & n231));
  assign n1254 = x7 & (x6 ? (n312 & ~n1256) : ~n1255);
  assign n1255 = (x0 | (~x4 & (~x1 | x2 | x3))) & (x1 | x2 | (~x4 & (~x0 | x3)));
  assign n1256 = x1 ? x2 : (~x2 & ~x3);
  assign n1257 = ~n837 & ((n169 & ~n1259) | (~x4 & ~n1258));
  assign n1258 = (x0 | x1 | x2 | x3 | ~x7) & (x7 | (x0 ? (x1 | (x2 & x3)) : (~x1 | (~x2 & ~x3))));
  assign n1259 = (x1 | ~x2 | ~x3) & (x2 | x3 | ~x7);
  assign n1260 = ~n1261 & n1264 & (x5 | ~n312 | n1263);
  assign n1261 = ~n1262 & (x3 ? ~x2 : (x2 | ~x7));
  assign n1262 = x0 ? (x1 | (x4 ? (x5 | ~x6) : (~x5 | x6))) : ((~x4 | (~x5 ^ ~x6)) & (~x5 | x6 | ~x1 | x4));
  assign n1263 = (~x1 | x2 | x3 | x6 | x7) & (x1 | ((~x3 | x6 | x7) & (~x2 | ((x6 | x7) & (x3 | ~x6 | ~x7)))));
  assign n1264 = (~n327 | ~n706) & (~x6 | ((~n460 | ~n327) & ~n1265));
  assign n1265 = ~x1 & ~x2 & (x0 ? (x4 & x5) : (~x4 & ~x5));
  assign z061 = n1267 | ~n1271 | (n343 & ~n1269);
  assign n1267 = ~n1268 & ~x7 & n159;
  assign n1268 = (x1 | x2 | (~x0 ^ x4)) & (x0 | x4 | (~x1 & ~x2));
  assign n1269 = (x0 | x2 | ~x3 | ~n693) & (~x0 | ~x2 | x3 | n1270);
  assign n1270 = x5 ? (x6 | ~x7) : x7;
  assign n1271 = (n1272 | n1273) & (n416 | n281 | (~n853 & n1272));
  assign n1272 = x0 & (x1 | x2);
  assign n1273 = (~x4 | ~x5 | ~x6 | ~x7) & (x4 | (x5 ? (x6 | ~x7) : (~x6 | x7)));
  assign z062 = n1275 | n1278 | n1279 | (n205 & ~n1277);
  assign n1275 = ~n1276 & ~x7 & n343;
  assign n1276 = (~x0 | ~x2 | x3 | ~x5 | ~x6) & (x0 | x6 | (x2 ? (x3 | ~x5) : ~x3));
  assign n1277 = (x0 | x2 | ~x5 | x6 | x7) & (~x0 | ~x2 | x5 | (x6 & ~x7));
  assign n1278 = ~n1272 & (n228 | n252);
  assign n1279 = ~x7 & n159 & (~x0 ^ (~x1 & ~x2));
  assign z063 = (~n300 & ~n1282) | (~x1 & (~n1283 | (~n300 & ~n1281)));
  assign n1281 = (x0 | x2 | ~x3 | ~x4 | ~x5) & (x5 | ((~x0 | ~x2 | x3 | ~x4) & (x0 | x4 | (~x2 ^ x3))));
  assign n1282 = x0 ^ (~x1 & (~x2 | (~x3 & ~x4)));
  assign n1283 = (x3 | n1284) & (~x3 | ~x6 | ~n401 | n1286);
  assign n1284 = (~x5 | n1285) & (x0 | x2 | x5 | ~x6);
  assign n1285 = (~x0 | ~x2 | ~x4 | x6 | x7) & (x0 | ~x6 | ((x4 | ~x7) & (x2 | (x4 & ~x7))));
  assign n1286 = x4 ^ (~x5 & x7);
  assign z064 = ~n1293 | (~x1 & (~n1288 | ~n1290));
  assign n1288 = (x3 | x5 | ~x7 | ~n401) & (x7 | n1289);
  assign n1289 = (x0 | x2 | ~x3 | ~x4 | ~x5) & (~x2 | ((x4 | ~x5 | x0 | ~x3) & (~x0 | x3 | (x4 & x5))));
  assign n1290 = (~x7 | ~n312 | n852 | ~n1132) & (x7 | n1291);
  assign n1291 = (x3 | ~x5 | n1292) & (~x3 | x5 | ~n401 | n446);
  assign n1292 = (~x0 | ~x2 | ~x4 | x6) & (x0 | ~x6 | (~x2 ^ x4));
  assign n1293 = (~n171 | ~n462) & (x7 | n1294);
  assign n1294 = (x0 & (x1 | x2)) | (~x1 & (x2 ? (~x4 & x5) : ~x0));
  assign z065 = ~x0 & (n1296 | ~n1300 | (~x5 & ~n1299));
  assign n1296 = ~x3 & ((n559 & n1297) | (x2 & ~n1298));
  assign n1297 = x4 & ~x1 & ~x2;
  assign n1298 = (~x1 | ~x4 | ~x5 | ~x6 | x7) & (x4 | ((x5 | ~x6 | x7) & (x6 | ~x7 | x1 | ~x5)));
  assign n1299 = (x1 | x2 | ~x3 | x4 | x6) & (~x1 | ~x2 | (x3 ? (~x4 | ~x6) : x6));
  assign n1300 = ~n1301 & n1302 & (x1 | ~n293 | ~n341);
  assign n1301 = ~n244 & (x2 ? (x3 ? ~x1 : x4) : (x1 | (x3 & x4)));
  assign n1302 = (~x1 & ~x2 & (~x4 | ~x6)) | (x1 & x2) | (x5 & ~x6) | (~x5 & x6);
  assign z066 = n1304 | ~n1312 | (~x3 & ~n1307);
  assign n1304 = ~x0 & (x2 ? ~n1306 : ~n1305);
  assign n1305 = (x3 | ((~x5 | ~x6 | x1 | ~x4) & (~x1 | (x4 ? (x5 | x6) : (~x5 | ~x6))))) & (x1 | ~x3 | x5 | (x4 ^ x6));
  assign n1306 = (x1 | x3 | x4 | ~x5 | ~x6) & (x6 | ((~x1 | ~x3 | ~x4 | x5) & (x1 | ((x4 | x5) & (~x3 | ~x4 | ~x5)))));
  assign n1307 = (x1 | n1309) & (x0 | ~x1 | ~n240 | ~n1308);
  assign n1308 = x7 & (~x4 ^ x5);
  assign n1309 = (x5 | n1311) & (x0 | ~x5 | ~n383 | n1310);
  assign n1310 = ~x2 ^ x4;
  assign n1311 = (x0 | ~x2 | x4 | ~x6 | x7) & (~x0 | ((~x6 | ~x7 | x2 | ~x4) & (x6 | x7 | ~x2 | x4)));
  assign n1312 = n1314 & ~n1315 & ~n1316 & (~x5 | n1313);
  assign n1313 = (x1 | x2 | ~x4 | (~x0 & ~x3)) & (x0 | ~x2 | (x1 ? (~x3 ^ ~x4) : (~x3 | x4)));
  assign n1314 = (~x0 | x1 | x2 | x3 | x4) & (x0 | ~x2 | (x1 ? (~x3 | x4) : (x3 | ~x4)));
  assign n1315 = ~x5 & n201 & (x0 ? n338 : n301);
  assign n1316 = n209 & n1317 & ~n1318;
  assign n1317 = x3 & ~x6;
  assign n1318 = (~x0 | x4 | ~x5 | x7) & (x0 | ~x4 | x5 | ~x7);
  assign z067 = n1327 | (~x1 & (~n1320 | ~n1324)) | ~n1329;
  assign n1320 = n1323 & (x2 | n1321);
  assign n1321 = (~x3 | n1322) & (x0 | x3 | x6 | ~n1308);
  assign n1322 = (~x0 | ((x4 | ~x5 | x6 | ~x7) & (~x6 | x7 | ~x4 | x5))) & (x0 | x4 | x5 | ~x6 | x7);
  assign n1323 = (~n990 | ~n383 | ~n633) & (n524 | n1249);
  assign n1324 = n1326 & (n437 | n1193) & (x0 | n1325);
  assign n1325 = (~x2 | x3 | ~x4 | x5 | ~x6) & (x2 | ((~x5 | ~x6 | x3 | ~x4) & (x5 | x6 | ~x3 | x4)));
  assign n1326 = (~x0 | x2 | x3 | x5 | x6) & (x0 | ~x2 | ~x3 | ~x5 | ~x6);
  assign n1327 = ~n244 & ~n1328;
  assign n1328 = (x0 | ((~x1 | x2 | x3 | ~x4) & (~x2 | ~x3 | x4))) & (x1 | ((~x3 | ~x4 | x0 | x2) & (x3 | (x0 ? (x2 ^ ~x4) : (x2 | x4)))));
  assign n1329 = ~n155 | (n1331 & n1332 & (n1330 | n419));
  assign n1330 = x2 ? (x3 | ~x4) : (~x3 | x4);
  assign n1331 = x2 ? (x3 ? (x4 ? ~x5 : (x5 | x6)) : (x4 | ~x5)) : (x3 ? (~x4 | x5) : (x4 ? (~x5 | ~x6) : x5));
  assign n1332 = (~n174 | ~n828) & (~n448 | ~n464);
  assign z068 = ~n1346 | n1343 | n1334 | n1337;
  assign n1334 = ~x0 & (x1 ? ~n1336 : ~n1335);
  assign n1335 = x2 ? ((~x3 | ~x4 | ~x5 | ~x6) & (x5 | x6 | x3 | x4)) : (x3 ? (x4 ? (x5 | ~x6) : (~x5 | x6)) : ((~x4 | x5 | x6) & (~x5 | ~x6)));
  assign n1336 = x5 ? ((x3 | x4 | x6) & (x2 | (x3 ? (~x4 | ~x6) : x6))) : ((x3 | ~x4 | ~x6) & (~x2 | ~x3 | x4 | x6));
  assign n1337 = ~x0 & (n1340 | (~x4 & (n1338 | n1339)));
  assign n1338 = x2 & ~n831 & (x1 ? (~x5 & x6) : (x5 & ~x6));
  assign n1339 = ~x5 & n209 & (x3 ? (x6 & x7) : (x6 ^ x7));
  assign n1340 = x4 & ((n1341 & n559) | (~x1 & ~n1342));
  assign n1341 = x3 & x1 & ~x2;
  assign n1342 = (x2 | x3 | ~x5 | x6 | ~x7) & (~x2 | ~x6 | x7 | (~x3 ^ x5));
  assign n1343 = ~n837 & ((n605 & ~n1345) | (x7 & ~n1344));
  assign n1344 = (~x0 | x1 | ~x2 | x3 | x4) & (x0 | ((~x3 | ~x4 | x1 | x2) & (~x1 | (x2 ? (x3 | ~x4) : (~x3 | x4)))));
  assign n1345 = x2 ? (~x3 | ~x4) : (x3 | x4);
  assign n1346 = ~n1349 & (n281 | n1348) & (~n157 | ~n1347);
  assign n1347 = x6 & x5 & ~x3 & x4;
  assign n1348 = (x0 | ~x1 | ~x3 | (x2 ^ x5)) & (x1 | (x0 ? ((x3 | x5) & (x2 | ~x3 | ~x5)) : (~x2 | (x3 ^ ~x5))));
  assign n1349 = n226 & ((~n737 & ~n374) | (n773 & n693));
  assign z069 = n1357 | ~n1360 | (~x3 & ~n1351);
  assign n1351 = ~n1352 & n1356 & (~x7 | ~n268 | n1355);
  assign n1352 = ~x0 & ((n825 & ~n1354) | (n1353 & n774));
  assign n1353 = ~x1 & x4;
  assign n1354 = (x1 | x2 | x5 | ~x7) & (x7 | (x1 ? (x2 ^ x5) : (~x2 ^ x5)));
  assign n1355 = (x2 | x5 | (~x4 ^ x6)) & (~x2 | x4 | ~x5 | x6);
  assign n1356 = (~n157 | ~n200) & (~n206 | ~n327);
  assign n1357 = ~n300 & (x3 ? ~n1359 : ~n1358);
  assign n1358 = x0 ? (x1 | ((~x2 | x4 | ~x5) & (~x4 | (x2 & x5)))) : ((x2 | x4 | ~x5) & (~x2 | (~x4 ^ ~x5)) & (~x1 | ((x2 | ~x4 | x5) & (x4 | ~x5))));
  assign n1359 = (~x0 | x1 | x2 | ~x4 | x5) & (x0 | (x4 ? ((~x2 | ~x5) & (x1 | (~x2 & ~x5))) : (x1 ? (x2 ^ ~x5) : (x2 | x5))));
  assign n1360 = ~n1364 & (~n279 | n1361) & (n697 | n1363);
  assign n1361 = (~x2 | n1362) & (x1 | x2 | ~x5 | n375);
  assign n1362 = (~x1 | ((~x4 | x5 | x6 | ~x7) & (~x6 | x7 | x4 | ~x5))) & (x1 | x4 | x5 | ~x6 | x7);
  assign n1363 = (x1 | ((~x3 | ~x5 | x0 | ~x2) & (~x0 | (x2 ? (x3 | x5) : ~x5)))) & (x0 | ((x2 | x3 | x5) & (~x1 | ((x3 | x5) & (x2 | (x3 & x5))))));
  assign n1364 = ~n183 & ((n157 & n1047) | (~x0 & ~n1365));
  assign n1365 = (x1 | ((~x2 | x3 | x4 | ~x5) & (~x4 | x5 | x2 | ~x3))) & (~x1 | x2 | ~x3 | ~x4 | ~x5);
  assign z070 = n1367 | ~n1376 | (~n300 & ~n1372);
  assign n1367 = ~x1 & (n1368 | n1370);
  assign n1368 = ~x0 & (x4 ? (n164 & ~n283) : ~n1369);
  assign n1369 = x2 ? (x3 ? (~x6 | x7) : (~x5 | ~x7)) : (x5 | (x3 ? (x6 | x7) : (~x6 | ~x7)));
  assign n1370 = x0 & (x2 ? (n174 & n176) : ~n1371);
  assign n1371 = (~x3 | ~x4 | x5 | x6 | ~x7) & (x3 | ((x5 | ~x6 | x7) & (x4 | (x5 ^ x7))));
  assign n1372 = ~n1374 & (n952 | n1373) & (x1 | n1375);
  assign n1373 = x2 ? (x4 | ~x5) : (~x4 | x5);
  assign n1374 = n155 & (x2 ? ((x4 & x5) | (~x3 & ~x4 & ~x5)) : (~x3 & x5));
  assign n1375 = (x0 | ~x2 | ~x3 | x5) & (x2 | ((x0 | (x3 ? ~x5 : (~x4 | x5))) & (~x3 | (x5 ? ~x4 : ~x0))));
  assign n1376 = ~n1377 & ~n1380 & (n1249 | n1379);
  assign n1377 = ~n183 & ((n788 & n327) | (~x3 & ~n1378));
  assign n1378 = (x0 | (x1 ? (x2 ? (x4 | ~x5) : (~x4 | x5)) : (x2 | ~x5))) & (x1 | (x2 ? (x5 | (~x0 & x4)) : (~x4 | ~x5)));
  assign n1379 = (~x3 | x4 | x1 | x2) & (x0 | (x1 ? (~x2 | (x3 ^ ~x4)) : (~x3 | ~x4)));
  assign n1380 = n155 & (x7 ? ~n1381 : (n293 & ~n1382));
  assign n1381 = (x2 | (x3 ? (~x5 | x6) : (x4 | x5))) & (~x4 | ((~x3 | ~x5 | x6) & (~x2 | x3 | x5 | ~x6)));
  assign n1382 = (x5 | ~x6) & (x4 | ~x5 | x6);
  assign z071 = n1389 | ~n1392 | (~x1 & ~n1384);
  assign n1384 = n1387 & (~x3 | (n1386 & (x0 | n1385)));
  assign n1385 = (x2 | ~x6 | ~x7) & (x6 | (x2 ? (x4 | (x5 ^ x7)) : (~x4 | x7)));
  assign n1386 = (x0 | ~x2 | ~x4 | n183) & (~x0 | x2 | (x4 ? ~n457 : n183));
  assign n1387 = (~n896 | ~n633) & (n416 | n1388);
  assign n1388 = (x0 | ~x2 | ~x3 | x4 | ~x6) & (x2 | ((x4 | x6 | x0 | ~x3) & (~x0 | ~x4 | (x3 ^ ~x6))));
  assign n1389 = ~x3 & (~n1391 | (~x0 & ~n1390));
  assign n1390 = (x1 | ~x2 | x4 | ~x5 | x6) & (~x1 | ((x4 | ~x5 | ~x6) & (x2 | (x4 ? (x5 | ~x6) : ~x5))));
  assign n1391 = (~x4 | x6 | x0 | ~x2) & (x1 | (x0 ? (x4 | (x2 ^ x6)) : (x2 | ~x6)));
  assign n1392 = (~x0 | x1 | ~x4 | n1393) & (x0 | ~x1 | (n1394 & (x4 | n1393)));
  assign n1393 = (~x2 | x3 | x5 | ~x6) & (x2 | (x3 ? (~x5 | ~x6) : (x5 | x6)));
  assign n1394 = (n423 | n1395) & (~x3 | n1396);
  assign n1395 = (x3 | ~x4 | ~x5 | ~x6) & (~x3 | (x4 ? (~x5 | x6) : (x5 | ~x6)));
  assign n1396 = ((x4 ^ x6) | (x2 ^ ~x7)) & (~x2 | x4 | ~x5 | ~x6 | ~x7) & (x6 | x7 | ~x4 | x5);
  assign z072 = n1400 | ~n1401 | (n879 & (n1398 | n1399));
  assign n1398 = x7 & ~n839 & (x3 ^ x6);
  assign n1399 = ~x7 & n268 & ((~x3 & ~x6) | (~x2 & x3 & x6));
  assign n1400 = ~n737 & ((~x0 & ~x4 & (x1 | x2)) | (~x1 & (x0 ? (~x2 & ~x4) : x4)));
  assign n1401 = ~n1403 & ~n1404 & n1405 & (~n653 | n1402);
  assign n1402 = (~x0 | x1 | ((x3 | x7) & (x2 | ~x3 | ~x7))) & (x0 | ~x1 | ~x3 | ~x7);
  assign n1403 = ~x0 & ((n209 & n710) | (x1 & n1183));
  assign n1404 = n140 & n845 & n896;
  assign n1405 = (~n231 | ~n715) & (~n158 | ~n334 | ~n462);
  assign z073 = n1412 | (~x1 & (~n1407 | ~n1411)) | ~n1414;
  assign n1407 = ~n1409 & (x3 | ~n1408 | ~n276);
  assign n1408 = x0 & x2;
  assign n1409 = ~x5 & ((n1408 & n703) | (~x6 & ~n1410));
  assign n1410 = (~x0 | ~x2 | x3 | x4) & (x0 | x2 | x7 | (~x3 ^ x4));
  assign n1411 = (x0 & (x2 | (~x4 & x5 & x6))) | (~x0 & (x4 | (~x2 & ~x5 & ~x6))) | (x4 & (~x5 | ~x6));
  assign n1412 = ~x0 & (n1413 | (n635 & n339));
  assign n1413 = x1 & x5 & x6 & (x4 ^ ~x7);
  assign n1414 = (~n626 | ~n938) & ((x5 & x6) | ~n1245);
  assign z074 = n1418 | n1419 | (~x0 & ~n1416) | ~n1422;
  assign n1416 = (x2 | n1417) & (~x1 | ~x2 | ~x6 | n283);
  assign n1417 = x1 ? (~x6 | ((~x4 | ~x5 | ~x7) & (x5 | x7))) : (x6 | ((x4 | ~x5 | x7) & (x5 | ~x7)));
  assign n1418 = ~x1 & (x0 ? (~x2 & (x5 ^ ~x6)) : (~x5 & (x2 | x6)));
  assign n1419 = ~x1 & (n1420 | (~x3 & n1408 & n631));
  assign n1420 = n159 & (n170 | (n401 & n1421));
  assign n1421 = x3 & ~x7;
  assign n1422 = x0 | ~x1 | (~n159 & (~n293 | ~n938));
  assign z075 = n1424 | ~n1435 | (~x1 & ~n1432);
  assign n1424 = ~x0 & (n1425 | ~n1429 | (~x4 & ~n1428));
  assign n1425 = ~x2 & ((n205 & ~n1427) | (x1 & n1426));
  assign n1426 = x3 & ((x6 & x7 & ~x4 & x5) | (~x6 & ~x7 & x4 & ~x5));
  assign n1427 = (x4 | ~x5 | ~x6 | x7) & (x5 | ((x6 | ~x7) & (~x4 | ~x6 | x7)));
  assign n1428 = x1 ? (x6 ? (~x7 | (~x2 & x5)) : x7) : (x2 | (x5 ? (x6 | ~x7) : (~x6 | x7)));
  assign n1429 = ~n1431 & (~n191 | ~n653 | ~n1430);
  assign n1430 = x1 & x2 & ~x3;
  assign n1431 = x1 & x4 & ((x5 & ~x6 & ~x7) | (x6 & x7));
  assign n1432 = n1433 & n1434 & (x6 | ~n401 | n1166);
  assign n1433 = x0 ? (~x6 | (x2 & (x3 | x4))) : (~x2 | x6);
  assign n1434 = (~n401 | ~n702) & (~x4 | ~n170 | ~n1132);
  assign n1435 = (~n365 | ~n717) & (~n159 | ~n176 | ~n928);
  assign z076 = n1437 | n1441 | ~n1449 | (n279 & ~n1446);
  assign n1437 = ~x3 & (x7 ? (n401 & ~n1440) : ~n1438);
  assign n1438 = (x1 | n1439) & (x0 | ~x1 | x2 | n437);
  assign n1439 = (x0 | x2 | ~x4 | ~x5) & (~x0 | ((x2 | ~x4 | x5 | ~x6) & (~x5 | x6 | ~x2 | x4)));
  assign n1440 = (x1 | ~x4 | x5 | x6) & (~x1 | (x4 ? (~x5 | x6) : (x5 | ~x6)));
  assign n1441 = ~n446 & (~n1443 | (~x2 & ~n1442));
  assign n1442 = (x0 | ~x1 | x3 | x5 | x7) & (x1 | ((x5 | x7 | x0 | ~x3) & (~x0 | x3 | (x5 ^ ~x7))));
  assign n1443 = ~n1444 & ~n1445 & (x3 | ~n570 | ~n231);
  assign n1444 = ~x0 & (x1 ? x7 : (x2 & ~x7));
  assign n1445 = ~x7 & x3 & ~x2 & x0 & ~x1;
  assign n1446 = (x1 | x2 | ~x6 | n1447) & (~x1 | ~x2 | n1448);
  assign n1447 = (~x5 | x7) & (x4 | x5 | ~x7);
  assign n1448 = (x4 | x5 | ~x6 | ~x7) & (~x4 | x6 | (x5 ^ x7));
  assign n1449 = (x2 | ~n140 | n1451) & (n281 | n1450);
  assign n1450 = (x0 | (x1 ? (~x7 | (~x2 ^ x3)) : (~x2 | x7))) & (x1 | x7 | (x2 ? x3 : ~x0));
  assign n1451 = (~x3 | ~x4 | x6 | x7) & (x3 | x4 | ~x7);
  assign z077 = n1454 | ~n1455 | (~x0 & ~n1453) | ~n1456;
  assign n1453 = (~x1 | ((x2 | ~x3) & (~x4 | x5 | ~x2 | x3))) & (x1 | ~x2 | x3 | x4 | ~x5) & (x2 | ~x4 | (~x3 & ~x5));
  assign n1454 = n795 & n268 & (x2 ? (~x4 & ~x6) : (x4 ^ x6));
  assign n1455 = (~n365 | ~n876) & (~n226 | (~x5 & ~n1047));
  assign n1456 = x0 | (n1457 & n1460 & (~n266 | n1459));
  assign n1457 = x5 ? (~n338 | n286) : n1458;
  assign n1458 = x1 ? ((x2 | x3 | x4 | ~x6) & (~x2 | ~x3 | ~x4 | x6)) : (x6 | (x2 ? (x3 | ~x4) : (~x3 | x4)));
  assign n1459 = (x1 | ~x2 | x3 | x4 | x5) & (~x1 | ((~x4 | x5 | x2 | x3) & (~x2 | ~x3 | x4 | ~x5)));
  assign n1460 = (~n1115 | ~n717) & (n1461 | (~x2 ^ x7));
  assign n1461 = (~x1 | x3 | x4 | x5 | x6) & (x1 | ((x3 | ~x4 | x5 | ~x6) & (~x5 | x6 | ~x3 | x4)));
  assign z078 = n1468 | (~x0 & (~n1463 | ~n1467)) | ~n1469;
  assign n1463 = (x5 | n1464) & (x4 | ~x5 | n1466);
  assign n1464 = ~n1465 & (~x1 | ~x4 | ~n266 | ~n845);
  assign n1465 = (~x3 ^ ~x7) & ((~x4 & ~x6) | (~x1 & x4 & x6));
  assign n1466 = x1 ? (~x6 | ((~x3 | ~x7) & (~x2 | x3 | x7))) : (x6 | (x3 ^ x7));
  assign n1467 = (x1 | ~x3 | (x4 ? (x5 | x6) : (~x5 | ~x6))) & (x3 | x4 | ((x5 | ~x6) & (~x1 | ~x5 | x6)));
  assign n1468 = x4 & ((n305 & ~n839) | (n304 & (n140 | ~n839)));
  assign n1469 = n1472 & (~n302 | ~n1471) & (~n365 | ~n1470);
  assign n1470 = ~x7 & x6 & ~x4 & x5;
  assign n1471 = ~x6 & (x3 ^ x5);
  assign n1472 = (~n393 | ~n472) & (x3 | ~n990 | ~n231);
  assign z079 = n1474 | n1479 | (n155 & ~n1483);
  assign n1474 = ~x1 & (n1477 | n1478 | n1475 | n1476);
  assign n1475 = x6 & ((n1095 & n340) | (n534 & n386));
  assign n1476 = ~n183 & (x0 ? (~x2 & n460) : (x2 & n382));
  assign n1477 = ~n374 & (n585 | (~x3 & ~x7 & n1408));
  assign n1478 = n242 & ((n312 & n228) | (x0 & n334));
  assign n1479 = ~n281 & (n1480 | n1481 | ~n1482);
  assign n1480 = ~x0 & ((x1 & x2 & x3 & ~x5) | (x5 & (~x1 | (~x2 & ~x3))));
  assign n1481 = n155 & (x5 ? (x7 & (x2 | x3)) : ((~x2 | ~x3) & ~x7));
  assign n1482 = (x2 | ~n997) & (x3 | (~n997 & (~n157 | ~n590)));
  assign n1483 = ~n1484 & n1485 & (~x2 | ~n773 | ~n339);
  assign n1484 = n151 & ((n266 & n795) | (n191 & n767));
  assign n1485 = (~x5 | x7 | ~x2 | ~x4) & (x4 | x5 | (x2 & x3) | ~x7);
  assign z080 = ~n1495 | (~x0 & (~n1487 | ~n1493));
  assign n1487 = x3 ? (n1489 & (x6 | n1488)) : n1490;
  assign n1488 = (~x7 | ((~x1 | ~x2 | x4 | x5) & (x1 | (x2 ? (x4 | ~x5) : (~x4 | x5))))) & (~x1 | x7 | (x2 ? (~x4 | x5) : (x4 | ~x5)));
  assign n1489 = n791 & (~x1 | ~n151 | ~n252);
  assign n1490 = x4 ? n1491 : n1492;
  assign n1491 = (~x2 | x5 | x6 | ~x7) & (x2 | ~x5 | ~x6 | x7);
  assign n1492 = (x5 | ((x1 | x2 | ~x6 | ~x7) & (~x1 | ((x6 | ~x7) & (x2 | ~x6 | x7))))) & (x1 | ~x5 | ((~x6 | x7) & (~x2 | x6 | ~x7)));
  assign n1493 = (x1 | x2 | ~x3 | ~n1095) & (x3 | n1494);
  assign n1494 = x1 ? (x2 | (x4 ? (x5 | ~x7) : (~x5 | x7))) : (~x2 | (x4 ? (~x5 | x7) : (x5 | ~x7)));
  assign n1495 = ~n1497 & n1500 & (n413 | n1496);
  assign n1496 = (x1 | ((x2 | x4) & (~x0 | (x3 ? x2 : x4)))) & (x0 | x4 | (x2 ? ~x1 : ~x3));
  assign n1497 = ~n300 & (~n1499 | (n1353 & ~n1498));
  assign n1498 = (~x0 | x5 | (~x2 ^ x3)) & (x0 | ~x2 | ~x3 | ~x5);
  assign n1499 = (~x0 | x1 | x2 | ~x4 | ~x5) & (x0 | (x1 ? (~x5 | (~x2 & ~x4)) : (~x4 | x5)));
  assign n1500 = (~n365 | ~n938) & (~n157 | ~n1501);
  assign n1501 = ~x5 & ~x3 & x4 & ~x7;
  assign z081 = n1508 | ~n1518 | (x2 ? ~n1512 : ~n1503);
  assign n1503 = ~n1504 & (~n155 | n1507);
  assign n1504 = ~x1 & (x6 ? ~n1505 : ~n1506);
  assign n1505 = (~x0 | ((~x4 | x5 | x7) & (~x5 | ~x7 | x3 | x4))) & (~x3 | ~x4 | ~x5 | ~x7) & (x0 | ((x3 | ~x4 | ~x7) & (x4 | x5 | x7)));
  assign n1506 = (~x0 | x4 | x5 | x7) & (x0 | (x4 ? (x7 | (~x3 & x5)) : (~x5 | ~x7)));
  assign n1507 = (~x4 | ~x5 | x6 | ~x7) & (~x6 | ((~x4 | x5 | x7) & (~x3 | (x4 ? x7 : (~x5 | ~x7)))));
  assign n1508 = ~n416 & ((~n1509 & ~n1510) | (~x0 & ~n1511));
  assign n1509 = x2 & x3;
  assign n1510 = (~x0 | x1 | (~x4 ^ x6)) & (x0 | ~x1 | x4 | x6);
  assign n1511 = x1 ? ((~x4 | ~x6 | x2 | x3) & (~x2 | ~x3 | x4)) : ((~x2 | (~x4 ^ ~x6)) & (~x4 | ((~x3 | ~x6) & (x2 | x3 | x6))));
  assign n1512 = ~n1517 & (x0 | (~n1513 & ~n1515 & n1516));
  assign n1513 = x1 & ~n1514;
  assign n1514 = (~x3 | ~x4 | ~x5 | x6 | x7) & (x3 | x5 | ~x7 | (~x4 ^ x6));
  assign n1515 = x1 & x4 & (x5 ? (~x6 & x7) : (x6 & ~x7));
  assign n1516 = x1 ? (x4 | n419) : ((~n176 | n419) & (x4 | ~n457));
  assign n1517 = n990 & n383 & n472;
  assign n1518 = ~n1519 & (~n158 | ~n590 | ~n928);
  assign n1519 = ~x1 & (x3 ? (n203 & ~n1138) : ~n1520);
  assign n1520 = (x0 | ~x2 | x4 | ~x5 | ~x7) & (~x0 | ((~x5 | ~x7 | x2 | ~x4) & (x5 | x7 | ~x2 | x4)));
  assign z082 = n1535 | n1533 | ~n1527 | n1522 | n1524;
  assign n1522 = ~x0 & ((n863 & n1341) | (~x3 & ~n1523));
  assign n1523 = (x1 | x2 | ~x4 | ~x5 | ~x6) & (~x2 | ((x5 | ~x6 | x1 | x4) & (~x1 | ~x5 | (x4 ^ ~x6))));
  assign n1524 = ~n283 & ((n155 & ~n1526) | (~x1 & ~n1525));
  assign n1525 = (x2 | ((~x0 | x6 | (x3 & x4)) & (~x6 | (x3 ? x0 : x4)))) & (x0 | ~x2 | (x3 ? x6 : ~x4));
  assign n1526 = (x2 | x3 | x4 | x6) & (~x2 | ~x6 | (~x3 & ~x4));
  assign n1527 = n1531 & (x1 | (n1528 & (x3 | n1529)));
  assign n1528 = (x0 | x2 | ~x3 | ~x5 | x6) & (~x0 | x5 | (x2 ? (x3 | x6) : (~x3 | ~x6)));
  assign n1529 = (~n722 | ~n559) & (~x6 | ~n692 | n1530);
  assign n1530 = x2 ? (x5 | ~x7) : (~x5 | x7);
  assign n1531 = (~n1532 | ~n928) & (~n157 | ~n176 | ~n1132);
  assign n1532 = x3 & x5 & x6;
  assign n1533 = ~n416 & ((n231 & n703) | (~x0 & ~n1534));
  assign n1534 = x1 ? (x2 ? (x4 | x6) : (x6 ? x3 : ~x4)) : ((~x2 | ~x3 | ~x4 | ~x6) & (x2 | x3 | x6));
  assign n1535 = x3 & (n1538 | (~x1 & (n337 | n1536)));
  assign n1536 = ~x7 & (x0 ? (~x2 & n1537) : (x2 & n825));
  assign n1537 = x4 & (~x5 ^ x6);
  assign n1538 = n707 & ((n338 & n1132) | (x2 & n856));
  assign z083 = n1546 | n1551 | (~x1 & ~n1540) | ~n1554;
  assign n1540 = x7 ? n1544 : (n1542 & (x6 | n1541));
  assign n1541 = x0 ? ((x4 | x5 | x2 | ~x3) & (~x4 | ~x5 | ~x2 | x3)) : (x3 | x4 | (x2 ^ ~x5));
  assign n1542 = x5 ? ((x6 | n1543) & (~x4 | ~x6 | ~n633)) : (~x6 | n1543);
  assign n1543 = (~x0 | x2 | x3 | ~x4) & (x0 | ~x2 | ~x3 | x4);
  assign n1544 = (~n386 | ~n846) & (~n317 | n1545);
  assign n1545 = (x2 & ~x5 & ~x6) | (x5 & (~x2 | x6));
  assign n1546 = ~n183 & (n1548 | ~n1549 | (~x0 & ~n1547));
  assign n1547 = x1 ? ((x2 | x3 | x4 | ~x5) & (~x2 | ~x3 | ~x4 | x5)) : (~x2 | x3 | (x4 ^ ~x5));
  assign n1548 = ~x0 & ((~x1 & ~x2 & ~x3 & x4) | (x1 & (x2 ? (~x3 & ~x4) : (x3 & x4))));
  assign n1549 = (~n788 | ~n157) & (~n268 | ~n1550);
  assign n1550 = ~x4 & ~x2 & x3;
  assign n1551 = n155 & (~n1553 | (~x7 & ~n1552));
  assign n1552 = (~x2 | x3 | ~x4 | ~x5 | x6) & (x2 | ((x3 | ~x4 | x5 | ~x6) & (~x5 | x6 | ~x3 | x4)));
  assign n1553 = (~x2 | ~x3 | ~x4 | ~x5 | ~x6) & (x2 | x3 | x4 | x5 | x6);
  assign n1554 = ~n1555 & n1559 & (~x7 | ~n238 | n1558);
  assign n1555 = ~n300 & ((n155 & ~n1557) | (~x1 & ~n1556));
  assign n1556 = (~x0 | ~x2 | x3 | (x4 & x5)) & (x2 | ~x3 | ((~x4 | ~x5) & (x0 | (~x4 & ~x5))));
  assign n1557 = x2 ? (~x4 | x5) : (x4 | (~x3 ^ x5));
  assign n1558 = (~x1 | x2 | ~x4 | ~x6) & (x1 | (x2 ? (~x4 | ~x6) : (x4 | x6)));
  assign n1559 = (~n157 | ~n703) & (~n1560 | (~x1 ^ x4));
  assign n1560 = ~x6 & x3 & ~x0 & x2;
  assign z084 = n1562 | ~n1566 | (x2 ? ~n1565 : ~n1564);
  assign n1562 = n176 & (x0 ? (n174 & n274) : ~n1563);
  assign n1563 = (x1 | ~x2 | x5 | x6 | x7) & (~x6 | ((~x1 | ~x5 | (~x2 ^ ~x7)) & (x1 | ~x2 | x5 | ~x7)));
  assign n1564 = (x7 | ((x1 | ~x3 | ~x4) & (x0 | (~x3 & (x1 | ~x4))))) & (x3 | ~x7 | (x0 ? x1 : x4));
  assign n1565 = (x4 | x7 | x1 | x3) & (x0 | ((~x3 | ~x7) & (~x1 | x3 | x7)));
  assign n1566 = n1568 & (x1 | (~n1567 & (~n471 | ~n633)));
  assign n1567 = n764 & ((n653 & n164) | (n990 & n293));
  assign n1568 = (~n1571 | ~n928) & (x4 | ~n1569 | ~n1570);
  assign n1569 = ~x5 & (x6 ^ x7);
  assign n1570 = x3 & ~x2 & x0 & ~x1;
  assign n1571 = ~x5 & ~x3 & x4 & x7;
  assign z085 = n1573 | ~n1574 | n1579 | (n510 & ~n1578);
  assign n1573 = ~x0 & ((~x1 & ~x2 & ~x3 & x4) | (x3 & ((x1 & x2) | ~x4)));
  assign n1574 = ~n1575 & ~n1576 & ~n1577 & (~n157 | ~n1017);
  assign n1575 = x4 & x3 & ~x2 & x0 & ~x1;
  assign n1576 = x5 & n151 & n155 & (~x3 ^ ~x6);
  assign n1577 = n169 & ((n305 & n215) | (n304 & n274));
  assign n1578 = x0 ? (x4 | (x2 ? (x3 | x6) : (~x3 | ~x6))) : (~x2 | ~x4 | (x3 ^ ~x6));
  assign n1579 = ~n336 & ((n523 & n472) | (n169 & ~n1580));
  assign n1580 = (~x1 | x3 | ~x5 | ~x7) & (x1 | ~x3 | x5 | x7);
  assign z086 = n1582 | n1585 | ~n1590 | (n155 & ~n1589);
  assign n1582 = x3 & ((n157 & n1470) | (~x0 & ~n1583));
  assign n1583 = (x2 | n1584) & (x1 | ~x2 | ~x4 | ~n448);
  assign n1584 = (~x1 | ((~x6 | ~x7 | x4 | ~x5) & (x6 | x7 | ~x4 | x5))) & (x1 | ~x4 | x5 | x6 | ~x7);
  assign n1585 = ~x3 & (n1588 | (~x1 & (n1586 | ~n1587)));
  assign n1586 = ~n336 & (x0 ? (~x4 & n228) : (x4 & n334));
  assign n1587 = (~x0 | x2 | ~x4 | n405) & (x0 | x4 | (x2 ? n405 : ~n339));
  assign n1588 = ~n336 & n155 & ~n229;
  assign n1589 = (x5 | ((x2 | ~x3 | x4 | x6) & (~x2 | (x3 ? (~x4 | ~x6) : x6)))) & (x2 | ~x5 | ~x6 | (x3 & ~x4));
  assign n1590 = n1593 & (x1 | (~n1591 & (~x3 | n1592)));
  assign n1591 = ~n244 & (x0 ? (~x2 & ~x4) : (x4 & (x2 ^ x3)));
  assign n1592 = (~x0 | x2 | ~x4 | ~x5 | x6) & (x0 | x4 | (x2 ? (~x5 | x6) : (x5 | ~x6)));
  assign n1593 = (~x0 | x3 | ~n990 | ~n274) & (x0 | n1594);
  assign n1594 = (~x1 | ~x2 | ~x3 | x4 | x5) & (x1 | ~x4 | (x2 ? (~x3 | ~x5) : (x3 | x5)));
  assign z087 = ~n1600 | (~x0 & (x3 ? ~n1599 : ~n1596));
  assign n1596 = (x6 | n1598) & (x2 | ~x6 | x7 | n1597);
  assign n1597 = (~x4 | ~x5) & (~x1 | x4 | x5);
  assign n1598 = (~x5 | ~x7 | x2 | ~x4) & (x4 | ((~x1 | x2 | x5 | ~x7) & (x1 | (x2 ? (~x5 ^ ~x7) : (~x5 | x7)))));
  assign n1599 = (~x1 | ~x2 | x4 | ~n252) & (x2 | ~x4 | ~n1569);
  assign n1600 = ~n1601 & n1606 & (n300 | n1604);
  assign n1601 = ~x1 & (x2 ? ~n1602 : ~n1603);
  assign n1602 = (x6 | (x0 ? (x3 | (~x4 ^ x5)) : (~x3 | (x4 ^ x5)))) & (x0 | ~x6 | ((x4 | ~x5) & (x3 | ~x4 | x5)));
  assign n1603 = x5 ? ((~x0 | x3 | x4 | ~x6) & (~x3 | ((~x4 | ~x6) & (x0 | x4 | x6)))) : ((x0 ^ x3) | (x4 ^ ~x6));
  assign n1604 = (x1 | n1605) & (x0 | ~x1 | ~n164 | n273);
  assign n1605 = x0 ? (x4 | (x2 ? (x3 | x5) : (~x3 | ~x5))) : (~x2 | ~x4 | (x3 ^ ~x5));
  assign n1606 = (~n155 | n1607) & (~n254 | n1608);
  assign n1607 = (~x4 | ((~x2 | x3 | x5 | ~x6) & (x2 | (x3 ? (~x5 | ~x6) : (x5 | x6))))) & (x2 | ~x3 | x4 | x5 | ~x6) & (~x2 | x6 | ((x4 | ~x5) & (~x3 | (x4 & ~x5))));
  assign n1608 = (~x2 | ~x4 | x5 | ~x6 | x7) & (x2 | (x4 ^ x5) | (x6 ^ ~x7));
  assign z088 = ~n1615 | n1623 | (~x1 & (~n1610 | ~n1620));
  assign n1610 = n1613 & (x3 | n1611);
  assign n1611 = (x7 | n1612) & (x0 | ~n448 | ~n338);
  assign n1612 = (x0 | x2 | x4 | x5 | ~x6) & (~x0 | ((~x5 | ~x6 | x2 | x4) & (~x2 | ~x4 | x5 | x6)));
  assign n1613 = (~n865 | ~n717) & (n964 | n1614);
  assign n1614 = (~x0 | x2 | ~x4 | x5 | x7) & (~x5 | ~x7 | x0 | x4);
  assign n1615 = n1617 & (n273 | n1616);
  assign n1616 = x0 ? (x1 | x2 | (x3 ^ ~x7)) : ((~x2 | x3 | ~x7) & (~x1 | ((x3 | ~x7) & (~x2 | ~x3 | x7))));
  assign n1617 = (n416 | n1618) & (~n155 | n1619);
  assign n1618 = (~x0 | x1 | ~x2 | x3 | x4) & (x0 | ~x3 | (x1 & x2) | ~x4);
  assign n1619 = (x5 | x7 | x3 | ~x4) & (~x3 | x4 | ((~x5 | ~x7) & (x2 | x5 | x7)));
  assign n1620 = ~n1622 & (x0 ? (~n164 | ~n594) : n1621);
  assign n1621 = (x2 | x3 | ~x4 | ~x5 | ~x7) & (~x2 | ~x3 | x4 | x5 | x7);
  assign n1622 = (n924 | n1017) & (x0 ? (~x2 & x7) : ~x7);
  assign n1623 = n155 & (n1624 | (x2 & n448 & n176));
  assign n1624 = ~x7 & n990 & ((x3 & ~x6) | (x2 & ~x3 & x6));
  assign z089 = n1626 | n1629 | n1631 | (n155 & ~n1635);
  assign n1626 = ~x1 & (x3 ? (x6 & ~n1628) : ~n1627);
  assign n1627 = x0 ? ((x4 | ~x6 | ~x7) & (~x2 | ~x4 | x6 | x7)) : ((~x4 | ~x6) & (x2 | ((~x6 | x7) & (x4 | x6 | ~x7))));
  assign n1628 = x0 ? (x2 | ~x7) : (~x4 & (x2 | x7));
  assign n1629 = n1630 & ((x2 & ~x4 & x7) | (x4 & (~x2 | ~x7)));
  assign n1630 = x6 & ~x0 & x1;
  assign n1631 = ~x1 & ((n203 & ~n695) | n1632 | ~n1633);
  assign n1632 = ~x4 & ~n848 & (x0 ? (~x3 & ~x7) : (x3 & x7));
  assign n1633 = x7 ? (n508 | ~n704) : (~n391 | n1634);
  assign n1634 = x4 ? (x5 ^ x6) : (x5 | ~x6);
  assign n1635 = n1638 & (x5 ? (~n787 | ~n1636) : n1637);
  assign n1636 = ~x4 & ~x2 & ~x3;
  assign n1637 = (~x2 | ~x4 | x6 | (x3 ^ ~x7)) & (x2 | ~x3 | x4 | ~x6 | x7);
  assign n1638 = x6 ? ((x2 | x4 | x5 | ~x7) & (~x2 | (x4 ? (~x5 | ~x7) : (x5 | x7)))) : ((x4 | ~x5 | x7) & (x2 | ~x4 | x5 | ~x7));
  assign z090 = x7 ? ~n1644 : (~n1641 | (~n281 & ~n1640));
  assign n1640 = (x3 | x5 | x0 | x2) & (x1 | (x0 ? (~x5 | (x2 & x3)) : x5));
  assign n1641 = n1643 & (~n653 | n1048) & (~n845 | n1642);
  assign n1642 = (~x0 | x1 | x4 | ~x5 | x6) & (x0 | ~x1 | ~x4 | x5 | ~x6);
  assign n1643 = (~x0 | x1 | x2 | ~x4 | x5) & (x0 | ((x4 | ~x5) & (~x1 | ~x2 | ~x4 | x5)));
  assign n1644 = ~n1646 & ~n1647 & n1648 & (~n146 | n1645);
  assign n1645 = x1 ? ((x3 | x4 | x6) & (x2 | (~x4 ^ ~x6))) : (~x2 | ((~x3 | x4 | x6) & (~x4 | ~x6)));
  assign n1646 = ~x0 & x4 & (x2 ? x5 : ~x1);
  assign n1647 = x5 & n151 & (x0 ? n201 : n940);
  assign n1648 = (~x2 | x4 | x5 | n952) & (x2 | (x4 ? (~x5 | n952) : (x5 | ~n268)));
  assign z091 = ~n1650 | (~x3 & ~n1656) | (~x2 & ~n1655);
  assign n1650 = n1653 & (x0 | (~n1651 & n1652));
  assign n1651 = n334 & ((x1 & ~x2 & ~x3 & x6) | (~x1 & ~x6 & (~x2 ^ x3)));
  assign n1652 = x1 ? (~x5 | (x2 ? ~x3 : (x3 | x6))) : (x5 | ~x6 | (x2 ^ x3));
  assign n1653 = (~n193 | ~n559) & (n852 | n1654);
  assign n1654 = (~x0 | x1 | x5 | x6 | x7) & (x0 | ((x1 | x5 | ~x6) & (~x5 | ((x6 | x7) & (~x1 | (x6 & x7))))));
  assign n1655 = (x0 | ~x1 | x5 | ~x6 | ~x7) & (x1 | ((x6 | ~x7 | x0 | x5) & (~x0 | ~x5 | (~x6 & ~x7))));
  assign n1656 = (~n327 | ~n716) & (x4 | (~n1657 & ~n1658));
  assign n1657 = ~n423 & (x5 ? (~x6 & n268) : (x6 & n155));
  assign n1658 = n274 & ((n146 & n383) | (x0 & n247));
  assign z092 = n1665 | (~x1 & (~n1661 | (~n183 & ~n1660)));
  assign n1660 = (x0 & ~x2 & ~x3 & (~x4 | ~x5)) | (x2 & ((~x0 & (x4 | x5)) | x3 | (x4 & x5)));
  assign n1661 = ~n1663 & n1664 & (x3 | n1662);
  assign n1662 = (~x0 | x2 | ~x4 | x5 | x6) & (x0 | ~x2 | x4 | ~x5 | ~x6);
  assign n1663 = ~x0 & x2 & x6 & (x3 | x4);
  assign n1664 = (~n567 | ~n391) & (~n633 | ~n1116);
  assign n1665 = n155 & (n1666 | ~n1667);
  assign n1666 = ~x3 & ((x2 & x7 & (x4 ^ x6)) | (~x6 & ~x7 & ~x2 & x4));
  assign n1667 = n1668 & (~n457 | ~n1636) & (~x3 | ~n1669);
  assign n1668 = x2 ? (x6 | x7) : (~x6 | ~x7);
  assign n1669 = ~x6 & (x2 ^ ~x7);
  assign z093 = ~n1676 | (~x3 & (~n1671 | ~n1673 | ~n1675));
  assign n1671 = (x7 | n1672) & (~x4 | ~x7 | ~n268 | n508);
  assign n1672 = (~x0 | x1 | x2 | ~x4 | x5) & (x0 | x4 | (x1 ? (x2 | x5) : (~x2 | ~x5)));
  assign n1673 = (~n312 | n1674) & (~n266 | ~n653 | ~n157);
  assign n1674 = (x1 | ~x2 | x5 | x6 | ~x7) & (~x1 | x2 | ~x5 | (~x6 ^ ~x7));
  assign n1675 = (x4 | ((x0 | ~x1 | ~x2 | ~x7) & (~x0 | x1 | (x2 ^ x7)))) & (x0 | ~x4 | ((~x2 | x7) & (~x1 | x2 | ~x7)));
  assign n1676 = (~x3 | x7 | x0 | ~x2) & (x2 | ~x7 | ((x1 | ~x3) & (x0 | (x1 & ~x3))));
  assign z094 = ~n1682 | n1678 | (~x7 & n205 & ~n1681);
  assign n1678 = ~x0 & ((x1 & ~n1680) | (n343 & n1679));
  assign n1679 = ~x5 & (x2 ? (~x3 & ~x6) : (x3 & x6));
  assign n1680 = (x2 | x3 | x4 | ~x5 | x6) & (~x2 | ~x3 | ~x4 | x5 | ~x6);
  assign n1681 = (~x0 | ~x4 | (x2 ? (~x5 | x6) : (x5 | ~x6))) & (x0 | ~x2 | x4 | x5 | ~x6);
  assign n1682 = n1685 & (x1 ? (x0 | n1684) : n1683);
  assign n1683 = (~x0 | x3 | (x4 & (~x2 | x5))) & (~x3 | ((x0 | (~x4 & ~x5)) & (x2 | ~x4 | ~x5)));
  assign n1684 = x4 ? (~x3 | (x2 & ~x5)) : (x3 | (~x2 & x5));
  assign n1685 = (~n938 | ~n1686) & (~n157 | ~n159 | ~n176);
  assign n1686 = ~x2 & ~x0 & x1 & x3;
  assign z095 = ~n1690 | n1693 | (~x0 & ~n1688) | ~n1694;
  assign n1688 = x6 ? (n1689 | (~x4 ^ ~x7)) : (~x7 | n1594);
  assign n1689 = (~x1 | x2 | ~x3 | ~x5) & (x1 | ~x2 | x3 | x5);
  assign n1690 = (~x5 & ((x2 & x3) | ~n1245)) | (n1691 & (~n1245 | (~x2 & x5)));
  assign n1691 = (~x6 | n1692) & (x2 | x4 | x6 | ~n155);
  assign n1692 = (~x0 | x1 | ~x2 | x3 | x4) & (x0 | ~x4 | (x1 ? (x2 | x3) : (~x2 | ~x3)));
  assign n1693 = n268 & ((n448 & n1550) | (~x3 & ~n147));
  assign n1694 = ~n1695 & (x5 | (~n1697 & (n281 | n868)));
  assign n1695 = ~x1 & ~n1696;
  assign n1696 = x5 ? (x0 ? (x2 | x4) : (~x4 | (x2 & x3))) : ((x0 | ~x2 | ~x3 | x4) & (~x0 | ~x4 | (~x2 ^ x3)));
  assign n1697 = n140 & ((x2 & ~x3 & ~x4 & ~x6) | (~x2 & ((x4 & x6) | (x3 & ~x4 & ~x6))));
  assign z096 = ~n1699 | n1707 | n1711 | (~x1 & ~n1709);
  assign n1699 = ~n1702 & (x0 | (n1700 & n1701)) & n1703;
  assign n1700 = (x1 | ~x3 | x5 | (~x2 ^ ~x6)) & (x3 | ((x1 | x2 | ~x5 | ~x6) & (~x1 | (x2 ? (~x5 | x6) : (x5 | ~x6)))));
  assign n1701 = (x1 | ~x2 | x5 | x6) & (~x1 | ~x5 | (x2 ^ x6));
  assign n1702 = n767 & n155 & (x2 ? n383 : n787);
  assign n1703 = ~n1705 & (~n231 | ~n1704) & (n1668 | n1706);
  assign n1704 = x6 & ~x3 & ~x5;
  assign n1705 = ~x6 & ~x5 & ~x2 & x0 & ~x1;
  assign n1706 = (~x0 | x1 | x3 | ~x5) & (x0 | ~x1 | ~x3 | x5);
  assign n1707 = n268 & ((n693 & n464) | (n1035 & ~n1708));
  assign n1708 = (~x3 | ~x4 | x5 | ~x7) & (x3 | x7 | (~x4 ^ x5));
  assign n1709 = (x5 | n1710) & (~x5 | ~x7 | ~n401 | n964);
  assign n1710 = (x0 | ~x2 | x3 | ~x6 | x7) & (~x0 | ((~x2 | x3 | x6 | ~x7) & (~x6 | x7 | x2 | ~x3)));
  assign n1711 = ~x0 & (n1713 | (n343 & n247 & ~n1712));
  assign n1712 = x2 ? (x3 | ~x7) : (~x3 | x7);
  assign n1713 = ~x6 & ((n1714 & n966) | (~n1345 & ~n1715));
  assign n1714 = ~x7 & x4 & ~x5;
  assign n1715 = x1 ? (x5 | ~x7) : (~x5 | x7);
  assign z097 = n1717 | n1721 | ~n1726 | (~n183 & ~n1724);
  assign n1717 = ~x2 & (n1720 | (~x1 & ~n1718));
  assign n1718 = (~x5 | n1719) & (x0 | x5 | ~n773 | ~n383);
  assign n1719 = x0 ? ((~x3 | x4 | x6 | ~x7) & (~x6 | x7 | x3 | ~x4)) : ((~x3 | ~x4 | ~x6 | x7) & (x3 | (x4 ? (x6 | x7) : (~x6 | ~x7))));
  assign n1720 = n1245 & ((n304 & n383) | (n787 & n305));
  assign n1721 = ~x1 & ((n240 & ~n1723) | (~x2 & ~n1722));
  assign n1722 = (x0 | x3 | x4 | x5 | ~x6) & (~x5 | ((x0 | ~x3 | x4 | x6) & (~x0 | (x3 ? (x4 | ~x6) : (~x4 | x6)))));
  assign n1723 = (~x0 | x3 | x4 | x5) & (x0 | ~x4 | (~x3 ^ x5));
  assign n1724 = (x1 | n1725) & (~n1686 | (~x4 & ~x5));
  assign n1725 = (x0 | ~x2 | x3 | x4) & (x5 | (x0 ? (x2 | (~x3 ^ x4)) : (~x2 | x3)));
  assign n1726 = ~n1728 & ~n1731 & (x1 | n1727) & n1733;
  assign n1727 = (x0 | ~x2 | ~x3 | x4 | ~x6) & (x2 | ((~x4 | x6 | x0 | ~x3) & (~x0 | (x3 ? (~x4 | ~x6) : (x4 | x6)))));
  assign n1728 = ~n300 & ((n401 & ~n1730) | (x2 & ~n1729));
  assign n1729 = (x1 | ((~x4 | ~x5 | x0 | ~x3) & (~x0 | x3 | (x4 ^ ~x5)))) & (x0 | ~x1 | ~x3 | (x4 & x5));
  assign n1730 = x1 ? (x3 | x4) : (x5 | (~x3 ^ x4));
  assign n1731 = ~n1732 & ~x6 & n301;
  assign n1732 = (~x0 | x1 | x3 | ~x5 | x7) & (x0 | ~x1 | ~x3 | (x5 ^ ~x7));
  assign n1733 = (~n607 | n1734) & (~n159 | ~n773 | ~n928);
  assign n1734 = x2 ? ~x6 : (~x4 | x6);
  assign z098 = n1736 | n1740 | n1743 | (n155 & ~n1748);
  assign n1736 = x5 & (n1738 | (x3 & (n299 | n1737)));
  assign n1737 = n401 & (x1 ? (~x4 & n266) : (x4 & ~n183));
  assign n1738 = ~x3 & ((n297 & n231) | (~x2 & ~n1739));
  assign n1739 = (x1 | (x4 ? (~x6 | (x0 ^ ~x7)) : (x6 | ~x7))) & (x0 | x4 | (x6 ^ ~x7));
  assign n1740 = ~x5 & (n1741 | (n266 & n157 & n176));
  assign n1741 = ~x0 & ((n293 & n200) | (~x6 & ~n1742));
  assign n1742 = (~x3 | ~x7 | (x2 ^ x4)) & (~x1 | x3 | x7 | (~x2 ^ x4));
  assign n1743 = ~x1 & (n1746 | n1747 | n1744 | n1745);
  assign n1744 = ~n1055 & ~n1057;
  assign n1745 = ~n537 & ((~x0 & x2 & n767) | ((x0 | ~x2) & n795));
  assign n1746 = ~n508 & ~x0 & ~n198;
  assign n1747 = ~n166 & (x4 ? (x7 & n293) : (~x7 & n164));
  assign n1748 = (~x7 & ((~x3 & (x4 | x5)) | (x2 & (~x3 | (x4 & x5))))) | (x3 & x7) | (~x2 & ~x4 & (x7 | (x3 & ~x5)));
  assign z099 = ~n1756 | (~x0 & (x4 ? ~n1750 : ~n1753));
  assign n1750 = x1 ? (x5 | n1752) : n1751;
  assign n1751 = (x2 | x3 | ~x5 | ~x6 | ~x7) & (~x3 | ((x6 | x7 | x2 | x5) & (~x2 | ~x6 | (x5 ^ ~x7))));
  assign n1752 = (~x2 | (x3 ? (x6 | ~x7) : (~x6 | x7))) & (x2 | x3 | x6 | ~x7);
  assign n1753 = (x1 | ~x2 | x5 | n1754) & (~x1 | n1755);
  assign n1754 = x3 ? (x6 | x7) : (~x6 | ~x7);
  assign n1755 = (x2 | ~x3 | ~x5 | ~x6 | x7) & (~x2 | x3 | x5 | x6 | ~x7);
  assign n1756 = ~n1757 & ~n1759 & n1763 & (~n203 | n1762);
  assign n1757 = n268 & (x2 ? (n176 & n693) : ~n1758);
  assign n1758 = (x4 | ((~x3 | x5 | x6 | x7) & (~x6 | ~x7 | x3 | ~x5))) & (x3 | ((x5 | ~x6 | x7) & (~x4 | ~x5 | x6 | ~x7)));
  assign n1759 = ~x2 & ((n155 & ~n1761) | (~x1 & ~n1760));
  assign n1760 = (x0 | ((~x5 | ~x6 | x3 | x4) & (~x3 | (x4 ? (~x5 | ~x6) : (x5 | x6))))) & (x5 | x6 | x3 | ~x4) & (~x0 | ((x3 | ((x5 | x6) & (~x4 | ~x5 | ~x6))) & (~x4 | x5 | x6) & (~x5 | ~x6 | ~x3 | x4)));
  assign n1761 = (x3 & x4) | (~x5 & ~x6) | (x6 & (x5 | (~x3 & ~x4)));
  assign n1762 = (x6 | ((x1 | ~x3 | ~x5) & (x3 | (x1 ? (~x4 ^ x5) : (x4 | x5))))) & (~x1 | ~x6 | (x3 ? (~x4 | ~x5) : (x4 | x5)));
  assign n1763 = (x1 | ~x5 | n1764) & (n1310 | ~n698);
  assign n1764 = (x0 | (x2 ? x3 : (~x3 | x4))) & (~x0 | x2 | ~x3 | ~x4) & (~x2 | x3 | x4);
  assign z100 = n1766 | ~n1772 | (x5 & ~n1770);
  assign n1766 = ~n183 & (n1768 | n1769 | (~x1 & ~n1767));
  assign n1767 = (x0 | ~x2 | ~x3 | x4 | x5) & (x2 | ((~x0 | (x3 ? (x4 | x5) : (~x4 | ~x5))) & (x4 | x5 | x0 | x3)));
  assign n1768 = ~n223 & (n853 | (n401 & (n940 | n201)));
  assign n1769 = n155 & ((~x2 & x3 & x4 & x5) | (x2 & ~x5 & (~x3 ^ x4)));
  assign n1770 = (~x6 | ~x7 | ~n176 | ~n462) & (x6 | x7 | n1771);
  assign n1771 = (x0 | ~x1 | x2 | (~x3 & x4)) & (x1 | ((~x0 | ((x3 | x4) & (x2 | ~x3 | ~x4))) & (~x2 | x3 | x4) & (x0 | ~x4 | (x2 ^ x3))));
  assign n1772 = ~n1773 & ~n1777 & n1779 & (~n155 | n1776);
  assign n1773 = ~x1 & ((x6 & ~n1774) | (~x3 & ~x6 & ~n1775));
  assign n1774 = (x0 | ~x2 | x4 | (x3 ^ x5)) & (x2 | ((~x4 | ~x5 | x0 | ~x3) & ((x4 ^ ~x5) | (~x0 ^ ~x3))));
  assign n1775 = x0 ? (x5 | (~x2 ^ x4)) : (~x2 | ~x4);
  assign n1776 = x3 ? (x2 ? (x4 ? (~x5 | ~x6) : x6) : (x5 | (x4 ^ ~x6))) : ((x2 | (x4 ? (~x5 | ~x6) : (x5 | x6))) & (~x2 | x4 | ~x5 | ~x6));
  assign n1777 = ~x0 & ((n297 & n1430) | (n201 & ~n1778));
  assign n1778 = (x2 | x4 | x6 | x7) & (~x2 | ~x4 | ~x6 | ~x7);
  assign n1779 = ~n266 | ((~n146 | n1780) & (~n157 | ~n158));
  assign n1780 = (x1 | x2 | x3 | x4) & (~x1 | ~x4 | (~x2 & x3));
  assign z101 = n1782 | n1787 | n1792 | (n155 & ~n1798);
  assign n1782 = ~x4 & (n1783 | (n279 & ~n1786));
  assign n1783 = ~x3 & (x5 ? ~n1784 : ~n1785);
  assign n1784 = (x0 | ~x2 | (x1 ? (~x6 | x7) : (x6 | ~x7))) & ((x0 ? (x1 | ~x2) : (~x1 | x2)) | (~x6 ^ ~x7));
  assign n1785 = (~x0 | x1 | x2 | x6 | x7) & (x0 | ((x1 | ~x7 | (x2 ^ x6)) & (~x6 | x7 | ~x1 | x2)));
  assign n1786 = (~x1 | ~x2 | ~x5 | ~x6 | ~x7) & (x2 | ((x6 | ~x7 | x1 | x5) & ((~x5 ^ x6) | (~x1 ^ ~x7))));
  assign n1787 = x4 & (x3 ? (n1788 | ~n1789) : ~n1790);
  assign n1788 = n1100 & ((~x1 & (x2 ? (~x5 & ~x6) : (x5 & x6))) | (x1 & ~x2 & x5 & ~x6));
  assign n1789 = (~n448 | ~n157) & (n183 | n999);
  assign n1790 = (~n457 | ~n157) & (~n1791 | (~x1 ^ x6));
  assign n1791 = ~x0 & x7 & (~x2 ^ x5);
  assign n1792 = ~x1 & (n1794 | ~n1795 | (~x0 & ~n1793));
  assign n1793 = (~x2 | x3 | ~x4 | ~x5 | x7) & (x2 | ((x5 | x7 | x3 | ~x4) & (~x3 | ~x7 | (~x4 ^ x5))));
  assign n1794 = n391 & ((x3 & ~x7 & (x4 ^ x5)) | (~x4 & ~x5 & x7));
  assign n1795 = n1797 & (n1055 | n1796);
  assign n1796 = (~x0 | ~x2 | x3 | x5) & (x0 | ~x5 | (x2 ^ x3));
  assign n1797 = (~x0 | x2 | x3 | ~x5 | ~x7) & (x0 | ~x2 | x5 | (x3 ^ x7));
  assign n1798 = (~x2 | (x3 ? (~x5 | x7) : (x5 | ~x7))) & (x5 | x7 | ~x3 | x4) & (x2 | ((~x5 | x7 | x3 | ~x4) & (~x3 | ((x5 | x7) & (~x4 | ~x5 | ~x7)))));
  assign z102 = n1800 | ~n1805 | n1811 | (n279 & ~n1813);
  assign n1800 = ~x3 & (n1801 | (n155 & ~n1804));
  assign n1801 = ~x1 & (x5 ? ~n1803 : ~n1802);
  assign n1802 = (x0 | ~x7 | ((x4 | x6) & (~x2 | ~x4 | ~x6))) & (x2 | ((~x6 | x7 | x0 | x4) & (~x0 | (x4 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n1803 = (~x0 | ~x2 | ~x4 | x6 | x7) & (x0 | ~x6 | (x2 ? x7 : (~x4 | ~x7)));
  assign n1804 = (x2 & (~x5 ^ x7)) | (~x2 & (~x5 ^ ~x7)) | (x4 & ~x6) | (x6 & (~x4 | (~x5 & ~x7)));
  assign n1805 = x0 ? (x1 | n1810) : (n1807 & (x1 | n1806));
  assign n1806 = (~x2 | x3 | ~x5 | x6) & (~x6 | ((x2 | ~x3 | x4 | x5) & (~x2 | (x3 ? ~x5 : (x4 | x5)))));
  assign n1807 = (~n1430 | ~n393) & (n1808 | n1809);
  assign n1808 = x3 ? (x4 ^ x6) : (~x4 | x6);
  assign n1809 = (x2 | x5) & (~x1 | ~x2 | ~x5);
  assign n1810 = (x3 | ((~x5 | ~x6 | x2 | x4) & (~x2 | ((x4 | ~x5 | x6) & (x5 | ~x6))))) & (x2 | ~x3 | (x4 ? x6 : x5));
  assign n1811 = ~n1138 & ~n1812;
  assign n1812 = (x3 | ~x6 | x0 | x2) & (x1 | ((~x3 | x6 | x0 | ~x2) & (~x0 | x2 | (~x3 ^ ~x6))));
  assign n1813 = ~n1815 & (x1 ? (~n457 | ~n338) : n1814);
  assign n1814 = (x2 | x4 | ~x5 | x6 | x7) & (~x2 | ~x7 | (x4 ? (~x5 | x6) : (x5 | ~x6)));
  assign n1815 = ~n416 & ((~x2 & n856) | (x1 & x2 & n825));
  assign z103 = ~n1828 | ~n1823 | n1817 | n1820;
  assign n1817 = ~n183 & ((n155 & ~n1819) | (~x1 & ~n1818));
  assign n1818 = (x2 | ((x0 | x3) & (~x4 | x5 | ~x0 | ~x3))) & (x0 | ((~x4 & ~x5) ? (~x2 | ~x3) : x3));
  assign n1819 = x4 ? (x3 | (x2 & ~x5)) : (~x3 | (~x2 & x5));
  assign n1820 = x5 & ((n254 & ~n1821) | (x3 & ~n1822));
  assign n1821 = x2 ? (x4 | x6) : (~x4 | ~x6);
  assign n1822 = (~x0 | x1 | x2 | ~x4 | x6) & (x0 | ~x1 | (x2 ? (~x4 | x6) : (x4 | ~x6)));
  assign n1823 = ~n1824 & (n300 | (~n1825 & ~n1826 & n1827));
  assign n1824 = n997 & (x2 ? (~x3 & ~x6) : (x3 & n825));
  assign n1825 = ~x0 & ((x1 & x2 & ~x3 & ~x4) | (x3 & (~x1 | ~x2) & x4));
  assign n1826 = n312 & ((n795 & n215) | (~x1 & n767));
  assign n1827 = (~n268 | ~n1636) & (~n157 | ~n924);
  assign n1828 = x7 ? (~n279 | n1832) : (~n1829 & ~n1831);
  assign n1829 = x5 & ((n155 & n1636) | (n268 & ~n1830));
  assign n1830 = (~x2 | x3 | ~x4 | x6) & (x2 | ~x3 | x4 | ~x6);
  assign n1831 = n795 & n203 & (x1 ? (x4 & x6) : (~x4 & ~x6));
  assign n1832 = (x1 | x2 | x4 | x5) & (~x1 | x6 | (x2 ? (~x4 | x5) : (x4 | ~x5)));
  assign z104 = n1834 | n1837 | ~n1842 | (n155 & ~n1841);
  assign n1834 = ~x1 & ((n1421 & ~n1836) | (~x3 & ~n1835));
  assign n1835 = (~x0 | ~x4 | ~x7 | (~x2 ^ x5)) & (x7 | ((x0 | ((x4 | ~x5) & (~x2 | ~x4 | x5))) & (x2 | ((x4 | ~x5) & (~x0 | ~x4 | x5)))));
  assign n1836 = (x2 | ~x4 | x5) & (x0 | (~x4 ^ x5));
  assign n1837 = ~x5 & (n1840 | (~x3 & (n1838 | n1839)));
  assign n1838 = n206 & n327;
  assign n1839 = x6 & n209 & ((~x4 & ~x7) | (x0 & x4 & x7));
  assign n1840 = x4 & n141 & n155 & ~n300;
  assign n1841 = (~x2 | ~x3 | ~x4 | ~x5 | ~x7) & (x7 | ((x3 | x4 | ~x5) & (x2 | (~x4 ^ x5))));
  assign n1842 = ~n1844 & n1845 & (n273 | n1843);
  assign n1843 = (~x3 | ((~x0 | x1 | x2 | ~x7) & (x0 | (x1 & x2) | x7))) & (x0 | x3 | x7 | (~x1 & ~x2));
  assign n1844 = n1100 & (x1 ? (x2 & n773) : (~x2 & n176));
  assign n1845 = (~n231 | ~n1223) & (~n990 | ~n383 | ~n1570);
  assign z105 = n1851 | ~n1854 | (~x3 & ~n1847);
  assign n1847 = ~n1850 & (x5 | (~n1849 & (x1 | n1848)));
  assign n1848 = (x0 | ~x2 | ~x6 | (x4 ^ x7)) & (x2 | ((x6 | ~x7 | x0 | x4) & (~x0 | (x4 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n1849 = n155 & ((n338 & n383) | (n787 & n301));
  assign n1850 = n231 & n243;
  assign n1851 = ~x0 & ((x4 & ~n1852) | (n343 & ~n1853));
  assign n1852 = (~x2 | (x1 ? (x3 ? (~x5 | ~x6) : (x5 | x6)) : (x3 | ~x5))) & (x1 | x2 | (~x5 ^ ~x6));
  assign n1853 = (x2 | ~x5 | ~x6) & (x5 | ((~x3 | x6) & (~x2 | (~x3 & x6))));
  assign n1854 = ~n1857 & (n244 | n1855) & (~n268 | n1856);
  assign n1855 = (x1 | (x0 ? (x4 | (~x2 ^ x3)) : (x2 | ~x4))) & (x0 | ((x2 | x3 | x4) & (~x1 | ~x2 | ~x3 | ~x4)));
  assign n1856 = x2 ? (x3 | ((x4 | ~x5 | ~x6) & (x5 | (~x4 & x6)))) : ((~x4 | ~x5) & (x5 | x6 | ~x3 | x4));
  assign n1857 = n209 & n1858 & (x0 ? n787 : n383);
  assign n1858 = x5 & x3 & ~x4;
  assign z106 = ~n1865 | (~x3 & ~n1860) | (~x1 & ~n1864);
  assign n1860 = (x1 | n1861) & (x0 | ~x1 | x5 | n1863);
  assign n1861 = (x5 | n1862) & (~x0 | ~x5 | ~n191 | ~n301);
  assign n1862 = x2 ? ((x4 | x6 | ~x7) & (~x6 | x7 | x0 | ~x4)) : ((~x4 | ~x6 | ~x7) & (~x0 | x4 | x6 | x7));
  assign n1863 = x2 ? (x4 ? (~x6 | x7) : (x6 | ~x7)) : (x4 ? (~x6 | ~x7) : (x6 | x7));
  assign n1864 = x2 ? ((x0 | ~x3 | ~x4) & (x3 | ((x4 | ~x5) & (~x0 | ~x4 | x5)))) : (x3 ? (x4 | x5) : (~x4 | ~x5));
  assign n1865 = n1866 & (~n1858 | n1871) & (x4 | n1868);
  assign n1866 = (~n155 | n1867) & (x3 | ~n1211 | ~n203);
  assign n1867 = x2 ? (x3 ? ~x4 : (x4 | ~x5)) : (x3 ? (x4 | x5) : (~x4 | ~x5));
  assign n1868 = x0 ? (x1 | n1870) : (x1 ? n1870 : (~x2 | ~n1869));
  assign n1869 = x6 & (~x3 ^ x5);
  assign n1870 = (~x2 | x3 | x5 | ~x6) & (x2 | ~x3 | ~x5 | x6);
  assign n1871 = (~x0 | x1 | x2 | ~x6 | x7) & (x0 | (x1 ^ x6) | (x2 ^ x7));
  assign z107 = x3 ? ~n1879 : (~n1875 | (~x7 & ~n1873));
  assign n1873 = (x1 | n1874) & (x0 | ~x1 | x5 | n446);
  assign n1874 = (~x4 | x5 | (x0 & x2) | ~x6) & (x6 | ((~x2 | x4 | x5) & (~x0 | ((x4 | x5) & (~x2 | ~x4 | ~x5)))));
  assign n1875 = ~n1247 & ~n1877 & (x1 | n1876);
  assign n1876 = (~x5 | ~x6 | x0 | x4) & (~x4 | x5 | ((~x0 | ~x2) & x6));
  assign n1877 = x7 & n990 & ~n1878;
  assign n1878 = x0 ? (x1 | ~x6) : (x1 ? (~x2 | ~x6) : x6);
  assign n1879 = ~n1880 & n1881 & (x6 | ~n990 | n839);
  assign n1880 = ~x4 & ((n140 & n359) | (~n1249 & ~n839));
  assign n1881 = (~n448 | ~n169) & (n1272 | (~n879 & ~n393));
  assign z108 = n1883 | n1887 | n1893 | (~n374 & ~n1892);
  assign n1883 = ~x6 & ((n317 & ~n530) | (~x3 & ~n1884));
  assign n1884 = (x5 | x7 | ~n312 | n1885) & (~x5 | n1886);
  assign n1885 = ~x1 ^ x2;
  assign n1886 = (x0 | ~x1 | x4 | ~x7) & (~x0 | x1 | (x2 ? (~x4 | x7) : (x4 | ~x7)));
  assign n1887 = ~n837 & (n1888 | n1889 | ~n1890);
  assign n1888 = ~x7 & ((~x0 & ((~x2 & x4) | (x1 & x2 & ~x4))) | (~x1 & (x0 ? (~x2 & ~x4) : x4)));
  assign n1889 = n155 & ((x2 & ~x3 & x4) | (~x2 & x3 & ~x4 & ~x7));
  assign n1890 = (~n231 | ~n715) & ~n1891;
  assign n1891 = ~x0 & x4 & (~x1 | ~x2) & x7;
  assign n1892 = (x0 & (x1 | (x2 & x3))) | (x7 & (~x0 | (~x2 & ~x3)));
  assign n1893 = x6 & ((n460 & n327) | n1265 | n1894);
  assign n1894 = n158 & n228 & n193;
  assign z109 = n1896 | ~n1900 | (n155 & ~n1899);
  assign n1896 = ~n416 & ((~n281 & ~n1897) | (~x4 & ~n1898));
  assign n1897 = (x1 | ~x2 | x3) & (x0 | (x1 & (x2 | x3)));
  assign n1898 = (~x0 | x1 | x2 | ~x6) & (x0 | ((x3 | x6 | x1 | x2) & (~x1 | ~x6 | (~x2 & ~x3))));
  assign n1899 = (x2 | ((x5 | ~x6 | x7) & (x4 | ~x5 | ~x7))) & (x6 | x7 | x4 | x5) & (~x4 | (x5 ? (x6 | ~x7) : (~x6 | x7)));
  assign n1900 = ~n1901 & (~n717 | ~n853) & (x0 | n1904);
  assign n1901 = ~x1 & ((n1202 & ~n1903) | (~x6 & ~n1902));
  assign n1902 = x0 ? (x2 | (x4 ? ~x7 : (x5 | x7))) : ((~x4 | ~x5 | ~x7) & (~x2 | x4 | x7));
  assign n1903 = x7 ? ~x5 : (x5 | (~x2 & ~x4));
  assign n1904 = (n1905 | ~n1906) & (~x3 | ~n209 | ~n609);
  assign n1905 = (~x2 | ~x3 | x5 | x6) & (x2 | x3 | ~x5 | ~x6);
  assign n1906 = x1 & x4 & x7;
  assign z110 = n1912 | ~n1915 | (~x6 & ~n1908);
  assign n1908 = ~n1911 & (x5 | (~n1910 & (x1 | n1909)));
  assign n1909 = (x2 | (x0 ? (x3 | x7) : (~x3 | x4))) & (x0 | x3 | (x7 ? x4 : ~x2));
  assign n1910 = x4 & n155 & ((x3 & x7) | (x2 & (x3 | x7)));
  assign n1911 = n158 & n590 & n193;
  assign n1912 = ~n300 & ((n155 & ~n1914) | (~x1 & ~n1913));
  assign n1913 = (~x4 | ((~x0 | (x2 ? (x3 | x5) : ~x5)) & (x2 | x5 | (x0 & ~x3)))) & (x0 | x4 | ((~x2 | ~x3) & ~x5));
  assign n1914 = x5 ? (~x4 | (~x2 & ~x3)) : x4;
  assign n1915 = (n413 | n1916) & (~x6 | ~n424 | n1917);
  assign n1916 = (x0 | ((~x1 | ~x2) & ~x4)) & (x1 | x4 | (x2 & (~x0 | x3)));
  assign n1917 = (x2 | (x1 ? (x4 | ~x7) : (~x4 | x7))) & (~x1 | x4 | x7 | (~x2 & ~x3));
  assign z111 = ~n1927 | (~x1 & (n1919 | n1925));
  assign n1919 = ~x2 & (n1921 | n1923 | (~x0 & ~n1920));
  assign n1920 = (~x3 | x4 | (x5 ? (x6 | x7) : (~x6 | ~x7))) & (~x6 | ((~x4 | x5 | x7) & (x3 | ~x5 | ~x7)));
  assign n1921 = ~n1922 & ((x3 & n825) | n897);
  assign n1922 = x0 ? (x5 | x7) : (~x5 | ~x7);
  assign n1923 = n1924 & ((x3 & x4 & ~x5) | ((~x3 | ~x4) & x5));
  assign n1924 = x7 & x0 & ~x6;
  assign n1925 = x2 & (x0 ? (n158 & n693) : ~n1926);
  assign n1926 = ((~x3 & ~x6) | (x4 ? (x5 | x7) : (~x5 | ~x7))) & (x4 | ((~x3 | ~x6 | ~x7) & (x6 | x7 | x3 | ~x5)));
  assign n1927 = ~n1928 & ~n1931 & (n229 | n1934);
  assign n1928 = n155 & (x2 ? ~n1929 : ~n1930);
  assign n1929 = (~x4 | x6 | x7 | (~x3 & x5)) & (~x7 | ((x4 | ~x5 | x6) & (x3 | (x4 ? (x5 | ~x6) : ~x5))));
  assign n1930 = (x6 | x7 | x3 | x5) & (~x4 | ((x5 | x6 | x7) & (~x6 | ~x7 | ~x3 | ~x5)));
  assign n1931 = ~n416 & (x3 ? ~n1933 : ~n1932);
  assign n1932 = (x1 | ((~x0 & x2) ? (~x4 | ~x6) : (x4 ^ ~x6))) & (x0 | ((x2 | x4 | x6) & (~x1 | (x2 ? x6 : (~x4 | ~x6)))));
  assign n1933 = (~x0 | x1 | x2 | x4 | ~x6) & (x0 | (x1 ? (x2 | (~x4 & x6)) : (~x2 | (~x4 ^ ~x6))));
  assign n1934 = (x1 | x2 | ((~x3 | x6) & (~x0 | x3 | ~x6))) & (x0 | ~x2 | (~x1 ^ ~x6));
  assign z112 = n1944 | n1936 | n1941;
  assign n1936 = x5 & (x2 ? ~n1939 : (n1937 | n1938));
  assign n1937 = ~n375 & (x0 ? ~x1 : x3);
  assign n1938 = n585 & ((x1 & x3 & ~x4 & x6) | (~x3 & ~x6 & (~x1 | x4)));
  assign n1939 = (~x0 | x4 | ~n383 | ~n205) & (x0 | n1940);
  assign n1940 = (x4 | x6 | (~x1 & ~x3) | ~x7) & (~x6 | x7 | (~x4 & (x1 | x3)));
  assign n1941 = ~n300 & ((n155 & ~n1943) | (~x1 & ~n1942));
  assign n1942 = x5 ? ((x2 | (x3 ^ x4)) & (x0 | (x2 ? (x3 | ~x4) : x4))) : (x0 ? (x2 ? (x3 | ~x4) : ~x3) : (~x2 | (x3 ^ x4)));
  assign n1943 = (x2 | ~x3 | x4 | x5) & (~x5 | (x2 ? (~x3 ^ x4) : (x3 ^ x4)));
  assign n1944 = ~x5 & (n1949 | (~x3 & (n1945 | ~n1946)));
  assign n1945 = ~x1 & (x0 ? (x2 ? (~x4 & ~x7) : x7) : (x4 & (~x2 ^ x7)));
  assign n1946 = ~n1948 & (x0 ? (~n209 | ~n680) : n1947);
  assign n1947 = (~x1 | ~x2 | ~x4 | x6 | ~x7) & (x1 | x4 | ((~x6 | x7) & (x2 | x6 | ~x7)));
  assign n1948 = ~x0 & x1 & (x2 ? (~x4 & ~x7) : (~x4 ^ ~x7));
  assign n1949 = x3 & ((n157 & n206) | (~x0 & ~n1950));
  assign n1950 = ((~x2 ^ x4) | (x6 ^ ~x7)) & (~x1 | ~x2 | ~x4 | ~x6 | ~x7) & (x1 | x2 | x4 | x6 | x7);
  assign z113 = n1962 | n1965 | (x3 ? ~n1952 : ~n1958);
  assign n1952 = ~n1953 & ~n1956 & (~n155 | n1957);
  assign n1953 = ~x1 & (x5 ? ~n1955 : ~n1954);
  assign n1954 = (~x0 | x2 | ~x4 | ~x6) & (x0 | x4 | x6);
  assign n1955 = (~x0 | x2 | ~x4 | x6 | x7) & (x0 | x4 | ((~x6 | x7) & (~x2 | x6 | ~x7)));
  assign n1956 = ~n419 & ((~x1 & (n169 | (x0 & ~x2))) | (~x2 & n169) | (~x0 & x1 & x2));
  assign n1957 = (x2 | x4 | x5 | x6 | x7) & (~x4 | ((x5 | ~x6 | ~x7) & (x6 | x7 | ~x2 | ~x5)));
  assign n1958 = ~n1961 & (x1 | (~n1960 & (x2 | n1959)));
  assign n1959 = (x0 | x4 | ~x6 | ~x7) & (~x0 | ~x4 | ((x6 | ~x7) & (~x5 | ~x6 | x7)));
  assign n1960 = ~x4 & n203 & ((x5 & ~x6 & ~x7) | (x6 & (~x5 | x7)));
  assign n1961 = n1630 & (x2 ? (x4 & n334) : (~x4 & x7));
  assign n1962 = ~n416 & ((n155 & ~n1964) | (~x1 & ~n1963));
  assign n1963 = (x6 | (x0 ? (x2 ? (x3 | ~x4) : (~x3 | x4)) : ((~x3 | ~x4) & (x2 | x3 | x4)))) & (x3 | ~x6 | (~x0 ^ x4));
  assign n1964 = (~x3 & ~x6) | (x2 & x4) | (x6 & (x3 | (~x2 & ~x4)));
  assign n1965 = ~n413 & ~n1966;
  assign n1966 = (x1 | x4 | (x0 ? x3 : (x2 | ~x3))) & (x0 | x3 | (~x1 & ~x4));
  assign z114 = n1976 | n1974 | ~n1972 | n1968 | n1971;
  assign n1968 = ~x1 & (~n1970 | (~x3 & ~n1969));
  assign n1969 = (~x5 | x7 | x0 | ~x4) & (~x0 | x4 | (x2 ? (x5 | ~x7) : (~x5 | x7)));
  assign n1970 = (n535 | (~x2 ^ x3)) & (x0 | (n535 & (x2 | ~x3 | ~n534)));
  assign n1971 = n155 & ((n141 & n1211) | (~x2 & n631));
  assign n1972 = n1973 & (n216 | ((~n140 | ~n141) & n839));
  assign n1973 = (~n1571 | ~n928) & (~n157 | ~n159 | ~n176);
  assign n1974 = ~n852 & (n1975 | (~x0 & n343 & n694));
  assign n1975 = n159 & ((~x0 & x7 & (~x1 ^ x4)) | (x0 & ~x1 & x4 & ~x7));
  assign n1976 = n312 & ((n247 & ~n1977) | (n339 & n966));
  assign n1977 = x1 ? (~x2 | x7) : (~x7 | (x2 ^ x3));
  assign z115 = ~n1984 | (~x1 & ~n1979);
  assign n1979 = x7 ? (~n1981 & (~x4 | n1980)) : n1982;
  assign n1980 = (x5 | ((x0 | x6 | (~x2 & ~x3)) & (~x0 | ~x2 | x3 | ~x6))) & (~x0 | x2 | ~x5 | (x3 ^ ~x6));
  assign n1981 = n312 & ((x3 & x5 & ~x6) | (x2 & ((x5 & ~x6) | (x3 & ~x5 & x6))));
  assign n1982 = ~n1983 & (~n203 | ~n631) & (~n170 | ~n393);
  assign n1983 = x0 & ~x2 & (x4 ? (x5 ^ ~x6) : (~x5 & x6));
  assign n1984 = ~n1626 & ~n1987 & (~n155 | n1985);
  assign n1985 = n1638 & (~n457 | ~n1550) & (~x4 | n1986);
  assign n1986 = (x2 | ~x3 | ~x5 | ~x6 | ~x7) & (~x2 | x5 | x6 | (x3 ^ ~x7));
  assign n1987 = n1630 & ((x4 & (~x7 | n845)) | (~x7 & n845) | (x2 & ~x4 & x7));
  assign z116 = ~n1993 | (~x0 & (n1989 | (n795 & ~n1992)));
  assign n1989 = x3 & (n1991 | (~x6 & ~n1990));
  assign n1990 = x1 ? ((x2 | x4 | x5 | ~x7) & (~x2 | ~x4 | ~x5 | x7)) : (x5 | (x2 ? (x4 | ~x7) : (~x4 | x7)));
  assign n1991 = ~x1 & ~x5 & x6 & (x4 ^ ~x7);
  assign n1992 = (~x7 | (~x1 ^ x2) | (x4 ^ x6)) & (x1 | x7 | (~x4 ^ x6));
  assign n1993 = x5 ? (n1997 & (~n268 | n1998)) : n1994;
  assign n1994 = n1996 & (x1 | n1995);
  assign n1995 = (x0 | x2 | x3 | ~x4 | ~x7) & (~x2 | ((~x4 | x7 | x0 | ~x3) & (~x0 | x3 | (x4 ^ ~x7))));
  assign n1996 = x0 ? (x1 | x2 | (x4 ^ ~x7)) : (~x1 | ((~x4 | x7) & (~x2 | x4 | ~x7)));
  assign n1997 = (~x7 | ~n209 | x3 | ~x4) & (x0 | (x4 ^ x7));
  assign n1998 = x7 ? ((~x2 | x3 | x4 | x6) & (x2 | ~x3 | ~x4 | ~x6)) : ((x2 & x3) | (~x4 ^ x6));
  assign z117 = ~n2005 | (~x0 & (n2000 | n2003 | ~n2004));
  assign n2000 = x7 & (n2002 | (x3 & ~n2001));
  assign n2001 = x1 ? ((x2 | x4 | x5 | ~x6) & (~x2 | ~x4 | ~x5 | x6)) : (x5 | (x2 ? (~x4 | ~x6) : (x4 | x6)));
  assign n2002 = ~x2 & ~x3 & ~x5 & (x1 ^ ~x6);
  assign n2003 = n334 & ((x1 & ~x2 & ~x3 & x6) | (~x1 & (x2 ? (x3 & x6) : (~x3 & ~x6))));
  assign n2004 = (x1 | ~x2 | x3 | x5 | ~x6) & (~x5 | ((x1 | x2 | ~x3 | x6) & (~x1 | (x2 ? (x3 | x6) : (~x3 | ~x6)))));
  assign n2005 = ~n2006 & ~n2008 & n2010 & (~n736 | n2007);
  assign n2006 = ~x0 & ((~x1 & ~x2 & ~x5 & x6) | (x5 & (x1 ? (~x2 ^ x6) : (x2 & ~x6))));
  assign n2007 = (~x0 | x1 | x3 | ~x5 | ~x6) & (x0 | ~x3 | (x1 ? (~x5 | x6) : (x5 | ~x6)));
  assign n2008 = n268 & n242 & ~n2009;
  assign n2009 = x7 ? ((x3 & x4) | ~x5) : x5;
  assign n2010 = ~n2011 & (x3 | ~n159 | ~n231);
  assign n2011 = x6 & x5 & ~x2 & x0 & ~x1;
  assign z118 = n2018 | n2021 | (~x0 & ~n2013) | ~n2022;
  assign n2013 = ~n2015 & (n300 | n2014) & (~x3 | n2016);
  assign n2014 = x1 ? (x2 | (x3 & (x4 | x5))) : (~x2 | ~x3 | (~x4 & ~x5));
  assign n2015 = ~n183 & (x1 ? (x2 & n460) : (~x2 & ~x3));
  assign n2016 = (~n635 | ~n339) & (~x1 | x7 | n2017);
  assign n2017 = (x2 | x4 | ~x5 | x6) & (~x2 | ~x4 | x5 | ~x6);
  assign n2018 = x2 & ((n169 & ~n2020) | (~x4 & ~n2019));
  assign n2019 = (x1 | x3 | ~x6 | (~x0 & ~x5)) & (x0 | ((~x1 | x6) & (x1 | ~x3 | x5 | ~x6)));
  assign n2020 = (~x1 | x6 | (~x3 ^ x5)) & (x1 | x3 | ~x5 | ~x6);
  assign n2021 = ~n498 & ((~x1 & x4 & x6) | (~x0 & (x1 ? (x4 & ~x6) : x6)));
  assign n2022 = ~n2023 & (~n445 | (~n357 & (~x1 | ~n856)));
  assign n2023 = ~n183 & n226 & (~x3 | n653 | n773);
  assign z119 = n2025 | ~n2027;
  assign n2025 = x3 & ((n155 & n521) | (~x1 & ~n2026));
  assign n2026 = (x0 | ~x2 | x4 | (~x5 ^ ~x7)) & (x2 | ((~x5 | x7 | x0 | x4) & (~x0 | ~x4 | (x5 ^ ~x7))));
  assign n2027 = ~n2029 & n2032 & (x3 ? n2028 : n2031);
  assign n2028 = (x1 | ~x7 | (x0 ? (x2 | x4) : (~x2 | ~x4))) & (x0 | x7 | ((x2 | ~x4) & (~x1 | ~x2 | x4)));
  assign n2029 = ~x6 & ((n279 & ~n2030) | (n217 & n231));
  assign n2030 = (x1 | x2 | x4 | x5 | ~x7) & (~x1 | ((~x5 | ~x7 | x2 | x4) & (~x2 | ~x4 | x5 | x7)));
  assign n2031 = (x2 & x7) | (~x2 & ~x7) | (x0 & (x1 | (x4 & ~x7)));
  assign n2032 = (~n231 | ~n1501) & (~n279 | ~n1132 | n2033);
  assign n2033 = (x1 | x2 | x4 | x7) & (~x1 | ~x2 | ~x4 | ~x7);
  assign z120 = ~n2036 | n2038 | (~x1 & ~n2035) | n2040;
  assign n2035 = (x0 | ((~x4 & ~x5) ? (~x2 | ~x3) : x3)) & (x2 | ((x3 | ~x4 | ~x5) & (~x0 | ~x3 | (x4 & x5))));
  assign n2036 = (~n155 | n2037) & (~n266 | ~n653 | ~n365);
  assign n2037 = x4 ? x3 : (~x3 | (~x2 & x5));
  assign n2038 = ~x0 & (n2039 | (x1 & n141 & n1211));
  assign n2039 = n338 & (x3 ^ x6) & (x1 ^ ~x5);
  assign n2040 = n312 & (n2041 | (n252 & n1341));
  assign n2041 = ~n336 & n205 & ~x5 & x7;
  assign z122 = z121;
  assign z123 = z121;
  assign z124 = z121;
  assign z125 = z121;
  assign z126 = z121;
  assign z127 = z121;
  assign z128 = z121;
endmodule


