// Benchmark "X_5_64" written by ABC on Tue Jun 27 01:56:52 2023

module X_5_64 ( 
    x0, x1, x2, x3, x4,
    z0, z1, z2, z3, z4, z5, z6, z7, z8  );
  input  x0, x1, x2, x3, x4;
  output z0, z1, z2, z3, z4, z5, z6, z7, z8;
  assign z0 = x2;
  assign z1 = x3;
  assign z2 = x4;
  assign z3 = 1'b0;
  assign z4 = x0;
  assign z5 = x1;
  assign z6 = 1'b0;
  assign z7 = x0;
  assign z8 = x1;
endmodule


