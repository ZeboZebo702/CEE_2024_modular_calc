module x_300_mod_997_reg(
    input [300:1] X,
    output [10:1] R
    );


assign R = X % 997;

endmodule
