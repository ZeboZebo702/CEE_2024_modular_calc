module x_400_mod_53(
    input [400:1] X,
    output [6:1] R
    );

wire [6:1] r1,r2,r3,r4,r5,r6,r7,r8,r9,r10,r11,r12,r13,r14,r15,r16,r17,
        r18,r19,r20,r21,r22,r23,r24,r25,r26,r27,r28,r29,r30,r31,r32,r33,
	r34,r35,r36,r37,r38,r39,r40,r41,r42,r43,r44,r45,r46,r47,r48,r49,
	r50,r51,r52,r53,r54,r55,r56,r57,r58,r59,r60,r61,r62,r63,r64,r65,r66;   

X_2 label2 (.x0(X[12]),.x1(X[11]),.x2(X[10]),.x3(X[9]),.x4(X[8]),.x5(X[7]),
.z0(r1[6]),.z1(r1[5]),.z2(r1[4]),.z3(r1[3]),.z4(r1[2]),.z5(r1[1]));

X_3 label3 (.x0(X[18]),.x1(X[17]),.x2(X[16]),.x3(X[15]),.x4(X[14]),.x5(X[13]),
.z0(r2[6]),.z1(r2[5]),.z2(r2[4]),.z3(r2[3]),.z4(r2[2]),.z5(r2[1]));

X_4 label4 (.x0(X[24]),.x1(X[23]),.x2(X[22]),.x3(X[21]),.x4(X[20]),.x5(X[19]),
.z0(r3[6]),.z1(r3[5]),.z2(r3[4]),.z3(r3[3]),.z4(r3[2]),.z5(r3[1]));

X_5 label5 (.x0(X[30]),.x1(X[29]),.x2(X[28]),.x3(X[27]),.x4(X[26]),.x5(X[25]),
.z0(r4[6]),.z1(r4[5]),.z2(r4[4]),.z3(r4[3]),.z4(r4[2]),.z5(r4[1]));

X_6 label6 (.x0(X[36]),.x1(X[35]),.x2(X[34]),.x3(X[33]),.x4(X[32]),.x5(X[31]),
.z0(r5[6]),.z1(r5[5]),.z2(r5[4]),.z3(r5[3]),.z4(r5[2]),.z5(r5[1]));

X_7 label7 (.x0(X[42]),.x1(X[41]),.x2(X[40]),.x3(X[39]),.x4(X[38]),.x5(X[37]),
.z0(r6[6]),.z1(r6[5]),.z2(r6[4]),.z3(r6[3]),.z4(r6[2]),.z5(r6[1]));

X_8 label8 (.x0(X[48]),.x1(X[47]),.x2(X[46]),.x3(X[45]),.x4(X[44]),.x5(X[43]),
.z0(r7[6]),.z1(r7[5]),.z2(r7[4]),.z3(r7[3]),.z4(r7[2]),.z5(r7[1]));

X_9 label9 (.x0(X[54]),.x1(X[53]),.x2(X[52]),.x3(X[51]),.x4(X[50]),.x5(X[49]),
.z0(r8[6]),.z1(r8[5]),.z2(r8[4]),.z3(r8[3]),.z4(r8[2]),.z5(r8[1]));

X_10 label10 (.x0(X[60]),.x1(X[59]),.x2(X[58]),.x3(X[57]),.x4(X[56]),.x5(X[55]),
.z0(r9[6]),.z1(r9[5]),.z2(r9[4]),.z3(r9[3]),.z4(r9[2]),.z5(r9[1]));

X_11 label11 (.x0(X[66]),.x1(X[65]),.x2(X[64]),.x3(X[63]),.x4(X[62]),.x5(X[61]),
.z0(r10[6]),.z1(r10[5]),.z2(r10[4]),.z3(r10[3]),.z4(r10[2]),.z5(r10[1]));

X_12 label12 (.x0(X[72]),.x1(X[71]),.x2(X[70]),.x3(X[69]),.x4(X[68]),.x5(X[67]),
.z0(r11[6]),.z1(r11[5]),.z2(r11[4]),.z3(r11[3]),.z4(r11[2]),.z5(r11[1]));

X_13 label13 (.x0(X[78]),.x1(X[77]),.x2(X[76]),.x3(X[75]),.x4(X[74]),.x5(X[73]),
.z0(r12[6]),.z1(r12[5]),.z2(r12[4]),.z3(r12[3]),.z4(r12[2]),.z5(r12[1]));

X_14 label14 (.x0(X[84]),.x1(X[83]),.x2(X[82]),.x3(X[81]),.x4(X[80]),.x5(X[79]),
.z0(r13[6]),.z1(r13[5]),.z2(r13[4]),.z3(r13[3]),.z4(r13[2]),.z5(r13[1]));

X_15 label15 (.x0(X[90]),.x1(X[89]),.x2(X[88]),.x3(X[87]),.x4(X[86]),.x5(X[85]),
.z0(r14[6]),.z1(r14[5]),.z2(r14[4]),.z3(r14[3]),.z4(r14[2]),.z5(r14[1]));

X_16 label16 (.x0(X[96]),.x1(X[95]),.x2(X[94]),.x3(X[93]),.x4(X[92]),.x5(X[91]),
.z0(r15[6]),.z1(r15[5]),.z2(r15[4]),.z3(r15[3]),.z4(r15[2]),.z5(r15[1]));

X_17 label17 (.x0(X[102]),.x1(X[101]),.x2(X[100]),.x3(X[99]),.x4(X[98]),.x5(X[97]),
.z0(r16[6]),.z1(r16[5]),.z2(r16[4]),.z3(r16[3]),.z4(r16[2]),.z5(r16[1]));

X_18 label18 (.x0(X[108]),.x1(X[107]),.x2(X[106]),.x3(X[105]),.x4(X[104]),.x5(X[103]),
.z0(r17[6]),.z1(r17[5]),.z2(r17[4]),.z3(r17[3]),.z4(r17[2]),.z5(r17[1]));

X_19 label19 (.x0(X[114]),.x1(X[113]),.x2(X[112]),.x3(X[111]),.x4(X[110]),.x5(X[109]),
.z0(r18[6]),.z1(r18[5]),.z2(r18[4]),.z3(r18[3]),.z4(r18[2]),.z5(r18[1]));

X_20 label20 (.x0(X[120]),.x1(X[119]),.x2(X[118]),.x3(X[117]),.x4(X[116]),.x5(X[115]),
.z0(r19[6]),.z1(r19[5]),.z2(r19[4]),.z3(r19[3]),.z4(r19[2]),.z5(r19[1]));

X_21 label21 (.x0(X[126]),.x1(X[125]),.x2(X[124]),.x3(X[123]),.x4(X[122]),.x5(X[121]),
.z0(r20[6]),.z1(r20[5]),.z2(r20[4]),.z3(r20[3]),.z4(r20[2]),.z5(r20[1]));

X_22 label22 (.x0(X[132]),.x1(X[131]),.x2(X[130]),.x3(X[129]),.x4(X[128]),.x5(X[127]),
.z0(r21[6]),.z1(r21[5]),.z2(r21[4]),.z3(r21[3]),.z4(r21[2]),.z5(r21[1]));

X_23 label23 (.x0(X[138]),.x1(X[137]),.x2(X[136]),.x3(X[135]),.x4(X[134]),.x5(X[133]),
.z0(r22[6]),.z1(r22[5]),.z2(r22[4]),.z3(r22[3]),.z4(r22[2]),.z5(r22[1]));

X_24 label24 (.x0(X[144]),.x1(X[143]),.x2(X[142]),.x3(X[141]),.x4(X[140]),.x5(X[139]),
.z0(r23[6]),.z1(r23[5]),.z2(r23[4]),.z3(r23[3]),.z4(r23[2]),.z5(r23[1]));

X_25 label25 (.x0(X[150]),.x1(X[149]),.x2(X[148]),.x3(X[147]),.x4(X[146]),.x5(X[145]),
.z0(r24[6]),.z1(r24[5]),.z2(r24[4]),.z3(r24[3]),.z4(r24[2]),.z5(r24[1]));

X_26 label26 (.x0(X[156]),.x1(X[155]),.x2(X[154]),.x3(X[153]),.x4(X[152]),.x5(X[151]),
.z0(r25[6]),.z1(r25[5]),.z2(r25[4]),.z3(r25[3]),.z4(r25[2]),.z5(r25[1]));

X_27 label27 (.x0(X[162]),.x1(X[161]),.x2(X[160]),.x3(X[159]),.x4(X[158]),.x5(X[157]),
.z0(r26[6]),.z1(r26[5]),.z2(r26[4]),.z3(r26[3]),.z4(r26[2]),.z5(r26[1]));

X_28 label28 (.x0(X[168]),.x1(X[167]),.x2(X[166]),.x3(X[165]),.x4(X[164]),.x5(X[163]),
.z0(r27[6]),.z1(r27[5]),.z2(r27[4]),.z3(r27[3]),.z4(r27[2]),.z5(r27[1]));

X_29 label29 (.x0(X[174]),.x1(X[173]),.x2(X[172]),.x3(X[171]),.x4(X[170]),.x5(X[169]),
.z0(r28[6]),.z1(r28[5]),.z2(r28[4]),.z3(r28[3]),.z4(r28[2]),.z5(r28[1]));

X_30 label30 (.x0(X[180]),.x1(X[179]),.x2(X[178]),.x3(X[177]),.x4(X[176]),.x5(X[175]),
.z0(r29[6]),.z1(r29[5]),.z2(r29[4]),.z3(r29[3]),.z4(r29[2]),.z5(r29[1]));

X_31 label31 (.x0(X[186]),.x1(X[185]),.x2(X[184]),.x3(X[183]),.x4(X[182]),.x5(X[181]),
.z0(r30[6]),.z1(r30[5]),.z2(r30[4]),.z3(r30[3]),.z4(r30[2]),.z5(r30[1]));

X_32 label32 (.x0(X[192]),.x1(X[191]),.x2(X[190]),.x3(X[189]),.x4(X[188]),.x5(X[187]),
.z0(r31[6]),.z1(r31[5]),.z2(r31[4]),.z3(r31[3]),.z4(r31[2]),.z5(r31[1]));

X_33 label33 (.x0(X[198]),.x1(X[197]),.x2(X[196]),.x3(X[195]),.x4(X[194]),.x5(X[193]),
.z0(r32[6]),.z1(r32[5]),.z2(r32[4]),.z3(r32[3]),.z4(r32[2]),.z5(r32[1]));

X_34 label34 (.x0(X[204]),.x1(X[203]),.x2(X[202]),.x3(X[201]),.x4(X[200]),.x5(X[199]),
.z0(r33[6]),.z1(r33[5]),.z2(r33[4]),.z3(r33[3]),.z4(r33[2]),.z5(r33[1]));

X_35 label35 (.x0(X[210]),.x1(X[209]),.x2(X[208]),.x3(X[207]),.x4(X[206]),.x5(X[205]),
.z0(r34[6]),.z1(r34[5]),.z2(r34[4]),.z3(r34[3]),.z4(r34[2]),.z5(r34[1]));

X_36 label36 (.x0(X[216]),.x1(X[215]),.x2(X[214]),.x3(X[213]),.x4(X[212]),.x5(X[211]),
.z0(r35[6]),.z1(r35[5]),.z2(r35[4]),.z3(r35[3]),.z4(r35[2]),.z5(r35[1]));

X_37 label37 (.x0(X[222]),.x1(X[221]),.x2(X[220]),.x3(X[219]),.x4(X[218]),.x5(X[217]),
.z0(r36[6]),.z1(r36[5]),.z2(r36[4]),.z3(r36[3]),.z4(r36[2]),.z5(r36[1]));

X_38 label38 (.x0(X[228]),.x1(X[227]),.x2(X[226]),.x3(X[225]),.x4(X[224]),.x5(X[223]),
.z0(r37[6]),.z1(r37[5]),.z2(r37[4]),.z3(r37[3]),.z4(r37[2]),.z5(r37[1]));

X_39 label39 (.x0(X[234]),.x1(X[233]),.x2(X[232]),.x3(X[231]),.x4(X[230]),.x5(X[229]),
.z0(r38[6]),.z1(r38[5]),.z2(r38[4]),.z3(r38[3]),.z4(r38[2]),.z5(r38[1]));

X_40 label40 (.x0(X[240]),.x1(X[239]),.x2(X[238]),.x3(X[237]),.x4(X[236]),.x5(X[235]),
.z0(r39[6]),.z1(r39[5]),.z2(r39[4]),.z3(r39[3]),.z4(r39[2]),.z5(r39[1]));

X_41 label41 (.x0(X[246]),.x1(X[245]),.x2(X[244]),.x3(X[243]),.x4(X[242]),.x5(X[241]),
.z0(r40[6]),.z1(r40[5]),.z2(r40[4]),.z3(r40[3]),.z4(r40[2]),.z5(r40[1]));

X_42 label42 (.x0(X[252]),.x1(X[251]),.x2(X[250]),.x3(X[249]),.x4(X[248]),.x5(X[247]),
.z0(r41[6]),.z1(r41[5]),.z2(r41[4]),.z3(r41[3]),.z4(r41[2]),.z5(r41[1]));

X_43 label43 (.x0(X[258]),.x1(X[257]),.x2(X[256]),.x3(X[255]),.x4(X[254]),.x5(X[253]),
.z0(r42[6]),.z1(r42[5]),.z2(r42[4]),.z3(r42[3]),.z4(r42[2]),.z5(r42[1]));

X_44 label44 (.x0(X[264]),.x1(X[263]),.x2(X[262]),.x3(X[261]),.x4(X[260]),.x5(X[259]),
.z0(r43[6]),.z1(r43[5]),.z2(r43[4]),.z3(r43[3]),.z4(r43[2]),.z5(r43[1]));

X_45 label45 (.x0(X[270]),.x1(X[269]),.x2(X[268]),.x3(X[267]),.x4(X[266]),.x5(X[265]),
.z0(r44[6]),.z1(r44[5]),.z2(r44[4]),.z3(r44[3]),.z4(r44[2]),.z5(r44[1]));

X_46 label46 (.x0(X[276]),.x1(X[275]),.x2(X[274]),.x3(X[273]),.x4(X[272]),.x5(X[271]),
.z0(r45[6]),.z1(r45[5]),.z2(r45[4]),.z3(r45[3]),.z4(r45[2]),.z5(r45[1]));

X_47 label47 (.x0(X[282]),.x1(X[281]),.x2(X[280]),.x3(X[279]),.x4(X[278]),.x5(X[277]),
.z0(r46[6]),.z1(r46[5]),.z2(r46[4]),.z3(r46[3]),.z4(r46[2]),.z5(r46[1]));

X_48 label48 (.x0(X[288]),.x1(X[287]),.x2(X[286]),.x3(X[285]),.x4(X[284]),.x5(X[283]),
.z0(r47[6]),.z1(r47[5]),.z2(r47[4]),.z3(r47[3]),.z4(r47[2]),.z5(r47[1]));

X_49 label49 (.x0(X[294]),.x1(X[293]),.x2(X[292]),.x3(X[291]),.x4(X[290]),.x5(X[289]),
.z0(r48[6]),.z1(r48[5]),.z2(r48[4]),.z3(r48[3]),.z4(r48[2]),.z5(r48[1]));

X_50 label50 (.x0(X[300]),.x1(X[299]),.x2(X[298]),.x3(X[297]),.x4(X[296]),.x5(X[295]),
.z0(r49[6]),.z1(r49[5]),.z2(r49[4]),.z3(r49[3]),.z4(r49[2]),.z5(r49[1]));

X_51 label51 (.x0(X[306]),.x1(X[305]),.x2(X[304]),.x3(X[303]),.x4(X[302]),.x5(X[301]),
.z0(r50[6]),.z1(r50[5]),.z2(r50[4]),.z3(r50[3]),.z4(r50[2]),.z5(r50[1]));

X_52 label52 (.x0(X[312]),.x1(X[311]),.x2(X[310]),.x3(X[309]),.x4(X[308]),.x5(X[307]),
.z0(r51[6]),.z1(r51[5]),.z2(r51[4]),.z3(r51[3]),.z4(r51[2]),.z5(r51[1]));

X_53 label53 (.x0(X[318]),.x1(X[317]),.x2(X[316]),.x3(X[315]),.x4(X[314]),.x5(X[313]),
.z0(r52[6]),.z1(r52[5]),.z2(r52[4]),.z3(r52[3]),.z4(r52[2]),.z5(r52[1]));

X_54 label54 (.x0(X[324]),.x1(X[323]),.x2(X[322]),.x3(X[321]),.x4(X[320]),.x5(X[319]),
.z0(r53[6]),.z1(r53[5]),.z2(r53[4]),.z3(r53[3]),.z4(r53[2]),.z5(r53[1]));

X_55 label55 (.x0(X[330]),.x1(X[329]),.x2(X[328]),.x3(X[327]),.x4(X[326]),.x5(X[325]),
.z0(r54[6]),.z1(r54[5]),.z2(r54[4]),.z3(r54[3]),.z4(r54[2]),.z5(r54[1]));

X_56 label56 (.x0(X[336]),.x1(X[335]),.x2(X[334]),.x3(X[333]),.x4(X[332]),.x5(X[331]),
.z0(r55[6]),.z1(r55[5]),.z2(r55[4]),.z3(r55[3]),.z4(r55[2]),.z5(r55[1]));

X_57 label57 (.x0(X[342]),.x1(X[341]),.x2(X[340]),.x3(X[339]),.x4(X[338]),.x5(X[337]),
.z0(r56[6]),.z1(r56[5]),.z2(r56[4]),.z3(r56[3]),.z4(r56[2]),.z5(r56[1]));

X_58 label58 (.x0(X[348]),.x1(X[347]),.x2(X[346]),.x3(X[345]),.x4(X[344]),.x5(X[343]),
.z0(r57[6]),.z1(r57[5]),.z2(r57[4]),.z3(r57[3]),.z4(r57[2]),.z5(r57[1]));

X_59 label59 (.x0(X[354]),.x1(X[353]),.x2(X[352]),.x3(X[351]),.x4(X[350]),.x5(X[349]),
.z0(r58[6]),.z1(r58[5]),.z2(r58[4]),.z3(r58[3]),.z4(r58[2]),.z5(r58[1]));

X_60 label60 (.x0(X[360]),.x1(X[359]),.x2(X[358]),.x3(X[357]),.x4(X[356]),.x5(X[355]),
.z0(r59[6]),.z1(r59[5]),.z2(r59[4]),.z3(r59[3]),.z4(r59[2]),.z5(r59[1]));

X_61 label61 (.x0(X[366]),.x1(X[365]),.x2(X[364]),.x3(X[363]),.x4(X[362]),.x5(X[361]),
.z0(r60[6]),.z1(r60[5]),.z2(r60[4]),.z3(r60[3]),.z4(r60[2]),.z5(r60[1]));

X_62 label62 (.x0(X[372]),.x1(X[371]),.x2(X[370]),.x3(X[369]),.x4(X[368]),.x5(X[367]),
.z0(r61[6]),.z1(r61[5]),.z2(r61[4]),.z3(r61[3]),.z4(r61[2]),.z5(r61[1]));

X_63 label63 (.x0(X[378]),.x1(X[377]),.x2(X[376]),.x3(X[375]),.x4(X[374]),.x5(X[373]),
.z0(r62[6]),.z1(r62[5]),.z2(r62[4]),.z3(r62[3]),.z4(r62[2]),.z5(r62[1]));

X_64 label64 (.x0(X[384]),.x1(X[383]),.x2(X[382]),.x3(X[381]),.x4(X[380]),.x5(X[379]),
.z0(r63[6]),.z1(r63[5]),.z2(r63[4]),.z3(r63[3]),.z4(r63[2]),.z5(r63[1]));

X_65 label65 (.x0(X[390]),.x1(X[389]),.x2(X[388]),.x3(X[387]),.x4(X[386]),.x5(X[385]),
.z0(r64[6]),.z1(r64[5]),.z2(r64[4]),.z3(r64[3]),.z4(r64[2]),.z5(r64[1]));

X_66 label66 (.x0(X[396]),.x1(X[395]),.x2(X[394]),.x3(X[393]),.x4(X[392]),.x5(X[391]),
.z0(r65[6]),.z1(r65[5]),.z2(r65[4]),.z3(r65[3]),.z4(r65[2]),.z5(r65[1]));

X_67 label67 (.x0(X[400]),.x1(X[399]),.x2(X[398]),.x3(X[397]),
.z0(r66[6]),.z1(r66[5]),.z2(r66[4]),.z3(r66[3]),.z4(r66[2]),.z5(r66[1]));


wire [8:1] R_temp_1,R_temp_2,R_temp_3,R_temp_4,R_temp_5,R_temp_6,R_temp_7,R_temp_8,R_temp_9,R_temp_10,R_temp_11,
	R_temp_12,R_temp_13,R_temp_14,R_temp_15,R_temp_16,R_temp_17,R_temp_18,R_temp_19,R_temp_20,R_temp_21,R_temp_22;

assign R_temp_1 = r1 + r2 + r3;
assign R_temp_2 = r4 + r5 + r6;
assign R_temp_3 = r7 + r8 + r9;
assign R_temp_4 = r10 + r11 + r12;
assign R_temp_5 = r13 + r14 + r15;
assign R_temp_6 = r16 + r17 + r18;
assign R_temp_7 = r19 + r20 + r21;
assign R_temp_8 = r22 + r23 + r24;
assign R_temp_9 = r25 + r26 + r27;
assign R_temp_10 = r28 + r29 + r30;
assign R_temp_11 = r31 + r32 + r33;
assign R_temp_12 = r34 + r35 + r36;
assign R_temp_13 = r37 + r38 + r39;
assign R_temp_14 = r40 + r41 + r42;
assign R_temp_15 = r43 + r44 + r45;
assign R_temp_16 = r46 + r47 + r48;
assign R_temp_17 = r49 + r50 + r51;
assign R_temp_18 = r52 + r53 + r54;
assign R_temp_19 = r55 + r56 + r57;
assign R_temp_20 = r58 + r59 + r60;
assign R_temp_21 = r61 + r62 + r63;
assign R_temp_22 = r64 + r65 + r66;

wire [9:1] R_temp_23,R_temp_24,R_temp_25,R_temp_26,R_temp_27,R_temp_28,R_temp_29;

assign R_temp_23 = R_temp_1 + R_temp_2 + R_temp_3;
assign R_temp_24 = R_temp_4 + R_temp_5 + R_temp_6;
assign R_temp_25 = R_temp_7 + R_temp_8 + R_temp_9;
assign R_temp_26 = R_temp_10 + R_temp_11 + R_temp_12;
assign R_temp_27 = R_temp_13 + R_temp_14 + R_temp_15;
assign R_temp_28 = R_temp_16 + R_temp_17 + R_temp_18;
assign R_temp_29 = R_temp_19 + R_temp_20 + R_temp_21;

wire [10:1] R_temp_30,R_temp_31,R_temp_32;

assign R_temp_30 = R_temp_23 + R_temp_24 + R_temp_25;
assign R_temp_31 = R_temp_26 + R_temp_27 + R_temp_28;
assign R_temp_32 = R_temp_29 + R_temp_22 + X[6:1];

wire [8:1] R_temp_33,R_temp_34,R_temp_35;

assign R_temp_33 = R_temp_30 [6:1] + 11 * R_temp_30 [7] +  22 * R_temp_30 [10:8]; 

assign R_temp_34 = 11 * R_temp_32 [7] + 22 * R_temp_32 [10:8] + R_temp_32 [6:1]; 

assign R_temp_35 = R_temp_31 [6:1] + 11* R_temp_31 [7] + 22 * R_temp_31 [10:8]; 


wire [8:1] R_temp_36,R_temp_37;

assign R_temp_36 = R_temp_33 [6:1] + 11 * R_temp_33 [7] + 22 * R_temp_33 [8] + R_temp_34 [6:1] + 22 * R_temp_34 [8]; 

assign R_temp_37 = R_temp_35 [6:1] + 11* R_temp_35 [7] + 22 * R_temp_35 [8] + 11 * R_temp_34 [7]; 


wire [7:1] R_temp_38;

assign R_temp_38 = R_temp_36 [6:1] + 11 * R_temp_36 [7] + 22 * R_temp_36 [8] + R_temp_37 [6:1] + 11 * R_temp_37 [7] + 22 * R_temp_37 [8];



reg [6:1]  R_temp;

always @(R_temp_38)
begin
  if (R_temp_38 >= 6'b110101  )
    R_temp <= R_temp_38 - 6'b110101;
  else
    R_temp <= R_temp_38;
end

assign R = R_temp;

endmodule