// Benchmark "128_128_mod" written by ABC on Thu Dec 01 02:19:21 2022

module const_128_128_mod ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z000, z001, z002, z003, z004, z005, z006, z007, z008, z009, z010, z011,
    z012, z013, z014, z015, z016, z017, z018, z019, z020, z021, z022, z023,
    z024, z025, z026, z027, z028, z029, z030, z031, z032, z033, z034, z035,
    z036, z037, z038, z039, z040, z041, z042, z043, z044, z045, z046, z047,
    z048, z049, z050, z051, z052, z053, z054, z055, z056, z057, z058, z059,
    z060, z061, z062, z063, z064, z065, z066, z067, z068, z069, z070, z071,
    z072, z073, z074, z075, z076, z077, z078, z079, z080, z081, z082, z083,
    z084, z085, z086, z087, z088, z089, z090, z091, z092, z093, z094, z095,
    z096, z097, z098, z099, z100, z101, z102, z103, z104, z105, z106, z107,
    z108, z109, z110, z111, z112, z113, z114, z115, z116, z117, z118, z119,
    z120, z121, z122, z123, z124, z125, z126, z127, z128, z129, z130, z131,
    z132, z133, z134, z135, z136, z137, z138, z139, z140, z141, z142, z143,
    z144, z145, z146, z147, z148, z149, z150, z151, z152, z153, z154, z155,
    z156, z157, z158, z159, z160, z161, z162, z163, z164, z165, z166, z167,
    z168, z169, z170, z171, z172, z173, z174, z175, z176, z177, z178, z179,
    z180, z181, z182, z183, z184, z185, z186, z187, z188, z189, z190, z191,
    z192, z193, z194, z195, z196, z197, z198, z199, z200, z201, z202, z203,
    z204, z205, z206, z207, z208, z209, z210, z211, z212, z213, z214, z215,
    z216, z217, z218, z219, z220, z221, z222, z223, z224, z225, z226, z227,
    z228, z229, z230, z231, z232, z233, z234, z235, z236, z237, z238, z239,
    z240, z241, z242, z243, z244, z245, z246, z247, z248, z249, z250, z251,
    z252, z253, z254, z255, z256, z257  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z000, z001, z002, z003, z004, z005, z006, z007, z008, z009, z010,
    z011, z012, z013, z014, z015, z016, z017, z018, z019, z020, z021, z022,
    z023, z024, z025, z026, z027, z028, z029, z030, z031, z032, z033, z034,
    z035, z036, z037, z038, z039, z040, z041, z042, z043, z044, z045, z046,
    z047, z048, z049, z050, z051, z052, z053, z054, z055, z056, z057, z058,
    z059, z060, z061, z062, z063, z064, z065, z066, z067, z068, z069, z070,
    z071, z072, z073, z074, z075, z076, z077, z078, z079, z080, z081, z082,
    z083, z084, z085, z086, z087, z088, z089, z090, z091, z092, z093, z094,
    z095, z096, z097, z098, z099, z100, z101, z102, z103, z104, z105, z106,
    z107, z108, z109, z110, z111, z112, z113, z114, z115, z116, z117, z118,
    z119, z120, z121, z122, z123, z124, z125, z126, z127, z128, z129, z130,
    z131, z132, z133, z134, z135, z136, z137, z138, z139, z140, z141, z142,
    z143, z144, z145, z146, z147, z148, z149, z150, z151, z152, z153, z154,
    z155, z156, z157, z158, z159, z160, z161, z162, z163, z164, z165, z166,
    z167, z168, z169, z170, z171, z172, z173, z174, z175, z176, z177, z178,
    z179, z180, z181, z182, z183, z184, z185, z186, z187, z188, z189, z190,
    z191, z192, z193, z194, z195, z196, z197, z198, z199, z200, z201, z202,
    z203, z204, z205, z206, z207, z208, z209, z210, z211, z212, z213, z214,
    z215, z216, z217, z218, z219, z220, z221, z222, z223, z224, z225, z226,
    z227, z228, z229, z230, z231, z232, z233, z234, z235, z236, z237, z238,
    z239, z240, z241, z242, z243, z244, z245, z246, z247, z248, z249, z250,
    z251, z252, z253, z254, z255, z256, z257;
  wire n268, n269, n270, n271, n272, n273, n274, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n291, n292,
    n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n322, n323, n324, n325, n326, n327, n328, n329, n330,
    n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
    n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n354, n355,
    n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n392, n393,
    n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n410, n411, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
    n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n455, n456,
    n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
    n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n487, n488, n489, n490, n491, n492, n493,
    n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512, n513, n514, n516, n517, n518,
    n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n542, n543,
    n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
    n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574, n575, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648, n649, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
    n679, n680, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n708, n709, n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735, n736, n737, n739, n740, n741,
    n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
    n766, n767, n768, n769, n770, n771, n772, n774, n775, n776, n777, n778,
    n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n828, n829,
    n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
    n842, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
    n855, n857, n858, n859, n860, n861, n862, n863, n864, n866, n867, n868,
    n869, n870, n871, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n906, n907,
    n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
    n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n931, n932,
    n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
    n945, n946, n947, n948, n950, n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n970,
    n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
    n983, n984, n985, n986, n987, n988, n989, n990, n992, n993, n994, n995,
    n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
    n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
    n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1067, n1068,
    n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
    n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
    n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1150, n1151, n1152,
    n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
    n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
    n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
    n1194, n1195, n1196, n1197, n1198, n1199, n1201, n1202, n1203, n1204,
    n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1221, n1222, n1223, n1224, n1225,
    n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
    n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1274, n1275, n1276, n1277,
    n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
    n1298, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
    n1319, n1320, n1321, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
    n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
    n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
    n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
    n1372, n1373, n1374, n1375, n1376, n1378, n1379, n1380, n1381, n1382,
    n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
    n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
    n1404, n1405, n1406, n1407, n1408, n1410, n1411, n1412, n1413, n1414,
    n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
    n1425, n1426, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1445, n1446,
    n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
    n1457, n1458, n1459, n1460, n1461, n1462, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
    n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
    n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
    n1499, n1500, n1501, n1502, n1503, n1504, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
    n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
    n1562, n1563, n1564, n1565, n1567, n1568, n1569, n1570, n1571, n1572,
    n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
    n1583, n1584, n1585, n1586, n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1613, n1614,
    n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
    n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
    n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1654, n1655, n1656,
    n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
    n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
    n1688, n1689, n1690, n1691, n1692, n1693, n1695, n1696, n1697, n1698,
    n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
    n1709, n1710, n1711, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1736, n1737, n1738, n1739, n1740, n1741,
    n1742, n1743, n1744, n1745, n1746, n1747, n1749, n1750, n1751, n1752,
    n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
    n1763, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1779, n1780, n1781, n1782, n1783, n1784,
    n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1795, n1796,
    n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
    n1807, n1808, n1809, n1810, n1811, n1813, n1814, n1815, n1816, n1817,
    n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
    n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
    n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
    n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1891,
    n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
    n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
    n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
    n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
    n1933, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
    n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
    n1975, n1976, n1977, n1978, n1979, n1981, n1982, n1983, n1984, n1985,
    n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
    n2007, n2008, n2009, n2010, n2011, n2012, n2014, n2015, n2016, n2017,
    n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
    n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
    n2039, n2040, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2062, n2063, n2064, n2065, n2066, n2068, n2069, n2070, n2071, n2072,
    n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2082, n2083,
    n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
    n2094, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
    n2105, n2106, n2107, n2108, n2109, n2110, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
    n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
    n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2147,
    n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
    n2158, n2159, n2160, n2161, n2163, n2164, n2165, n2166, n2167, n2168,
    n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
    n2179, n2180, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
    n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2226, n2227, n2228, n2229, n2230, n2231,
    n2232, n2233, n2234, n2235, n2236, n2237, n2239, n2240, n2241, n2242,
    n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
    n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2272, n2273, n2274,
    n2275, n2276, n2277, n2278, n2279, n2280, n2282, n2283, n2284, n2285,
    n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2297, n2298, n2299, n2301, n2302, n2303, n2304, n2305, n2306,
    n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2315, n2316, n2317,
    n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2328,
    n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
    n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
    n2360, n2361, n2362, n2363, n2364, n2365, n2367, n2368, n2369, n2370,
    n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
    n2381, n2382, n2383, n2384, n2385, n2387, n2388, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
    n2402, n2403, n2404, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2423,
    n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
    n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
    n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
    n2465, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
    n2486, n2487, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
    n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
    n2507, n2508, n2509, n2510, n2511, n2513, n2514, n2515, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
    n2528, n2529, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
    n2539, n2540, n2541, n2542, n2543, n2544, n2546, n2547, n2548, n2549,
    n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2566, n2567, n2568, n2569, n2570,
    n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
    n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2600, n2601, n2602,
    n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
    n2613, n2614, n2615, n2616, n2618, n2619, n2620, n2621, n2622, n2623,
    n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
    n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
    n2645, n2646, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661, n2663, n2664, n2665, n2666,
    n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
    n2677, n2678, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
    n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
    n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
    n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
    n2719, n2720, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
    n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2739, n2740,
    n2741, n2742, n2743, n2744, n2745, n2746, n2748, n2749, n2750, n2751,
    n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2760, n2761, n2762,
    n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2772, n2773,
    n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2782, n2783, n2784,
    n2785, n2786, n2787, n2788, n2790, n2791, n2792, n2793, n2794, n2795,
    n2796, n2797, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
    n2808, n2809, n2810, n2811, n2812, n2814, n2815, n2816, n2817, n2818,
    n2819, n2820, n2821, n2822, n2823, n2824, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2836, n2837, n2838, n2839, n2840,
    n2841, n2842, n2843, n2845, n2846, n2847, n2848, n2849, n2850, n2852,
    n2853, n2854, n2855, n2856, n2857, n2859, n2860, n2861, n2862, n2863,
    n2865, n2866, n2867, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
    n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
    n2887, n2888, n2889, n2890, n2892, n2893, n2894, n2895, n2896, n2897,
    n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
    n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
    n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2929,
    n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
    n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2955, n2956, n2957, n2958, n2959, n2960,
    n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
    n2971, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
    n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2990, n2991, n2992,
    n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
    n3003, n3004, n3005, n3006, n3007, n3009, n3010, n3011, n3012, n3013,
    n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
    n3024, n3025, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
    n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
    n3045, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
    n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
    n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
    n3077, n3078, n3079, n3080, n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
    n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
    n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3117, n3118, n3119,
    n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
    n3130, n3131, n3132, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
    n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3151,
    n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
    n3162, n3163, n3164, n3165, n3167, n3168, n3169, n3170, n3171, n3172,
    n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3182, n3183,
    n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3194,
    n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210, n3212, n3213, n3214, n3215,
    n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
    n3226, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
    n3237, n3238, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3248,
    n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3259,
    n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3268, n3269, n3270,
    n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3279, n3280, n3281,
    n3282, n3283, n3284, n3285, n3287, n3288, n3289, n3290, n3291, n3292,
    n3293, n3294, n3295, n3296, n3297, n3298, n3300, n3301, n3302, n3303,
    n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3314,
    n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
    n3325, n3326, n3327, n3328, n3330, n3331, n3332, n3333, n3334, n3335,
    n3336, n3337, n3338, n3339, n3341, n3342, n3343, n3344, n3345, n3346,
    n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3356, n3357,
    n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
    n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
    n3389, n3390, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
    n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
    n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3430, n3431,
    n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
    n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
    n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
    n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3471, n3472, n3473,
    n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
    n3484, n3485, n3486, n3487, n3489, n3490, n3491, n3492, n3493, n3494,
    n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
    n3505, n3506, n3507, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
    n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3526,
    n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
    n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
    n3548, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
    n3559, n3560, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
    n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3579, n3580,
    n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
    n3601, n3602, n3604, n3605, n3607, n3608, n3609, n3610, n3611, n3612,
    n3613, n3614, n3615, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
    n3624, n3625, n3626, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
    n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3643, n3644, n3645,
    n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
    n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3665, n3666,
    n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
    n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3685, n3686, n3687,
    n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
    n3698, n3699, n3700, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
    n3709, n3710, n3711, n3712, n3713, n3714, n3716, n3717, n3718, n3719,
    n3720, n3721, n3722, n3723, n3725, n3726, n3727, n3728, n3729, n3730,
    n3732, n3733, n3734, n3735, n3736, n3737, n3739, n3740, n3741, n3742,
    n3743, n3744, n3745, n3746, n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3756, n3757, n3758, n3759, n3760, n3762, n3763, n3764, n3765,
    n3766, n3767, n3768, n3769, n3770, n3771, n3773, n3774, n3775, n3776,
    n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3786, n3787,
    n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
    n3798, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
    n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
    n3819, n3820, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
    n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
    n3840, n3841, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
    n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
    n3861, n3862, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
    n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3882,
    n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
    n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3903,
    n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
    n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3923, n3924,
    n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
    n3935, n3936, n3937, n3938, n3939, n3941, n3942, n3943, n3944, n3945,
    n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
    n3956, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
    n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3977,
    n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
    n3988, n3989, n3990, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
    n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4008, n4009,
    n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
    n4020, n4021, n4022, n4023, n4024, n4025, n4027, n4028, n4029, n4030,
    n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
    n4041, n4042, n4043, n4044, n4046, n4047, n4048, n4049, n4050, n4051,
    n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
    n4062, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
    n4073, n4074, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
    n4084, n4086, n4087, n4088, n4089, n4090, n4092, n4093, n4094, n4095,
    n4096, n4097, n4099, n4101, n4102, n4103, n4106, n4108, n4109, n4110,
    n4112, n4113, n4114, n4115, n4116, n4118, n4119, n4120, n4121, n4122,
    n4123, n4124, n4125, n4126, n4128, n4129, n4130, n4131, n4132, n4133,
    n4134, n4135, n4136, n4137, n4138, n4139, n4141, n4142, n4143, n4144,
    n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
    n4155, n4156, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
    n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
    n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
    n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4197,
    n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
    n4208, n4209, n4210, n4211, n4213, n4214, n4215, n4216, n4217, n4218,
    n4219, n4220, n4221, n4222, n4224, n4225, n4226, n4227, n4228, n4229,
    n4230, n4231, n4232, n4233, n4234, n4236, n4237, n4238, n4239, n4240,
    n4241, n4242, n4243, n4244, n4245, n4247, n4248, n4249, n4250, n4251,
    n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4262, n4263,
    n4264, n4265, n4266, n4268, n4269, n4271, n4273, n4274, n4275, n4276,
    n4277, n4278, n4279, n4281, n4283, n4284, n4285, n4286, n4287, n4288;
  assign z250 = 1'b0;
  assign z000 = ~x0 & (~n268 | ~n274);
  assign n268 = n271 & ~n272 & (~n269 | (~n270 & ~n273));
  assign n269 = ~x3 & ~x1 & ~x2;
  assign n270 = x7 & ~x6 & ~x4 & ~x5;
  assign n271 = x1 ^ ~x2;
  assign n272 = x3 & ~x1 & ~x2;
  assign n273 = x6 & ~x4 & ~x5;
  assign n274 = x3 | (x1 ? (~x2 | (x4 & x5)) : (x2 | (~x4 & ~x5)));
  assign z001 = n281 | ~n286 | (n276 & ~n277);
  assign n276 = ~x1 & ~x3;
  assign n277 = x0 ? (~n278 | ~n280) : (x6 | n279);
  assign n278 = x2 & x4;
  assign n279 = (~x2 | ~x4 | ~x5 | x7) & (x2 | x4 | x5 | ~x7);
  assign n280 = ~x7 & ~x5 & x6;
  assign n281 = n285 & ((~x1 & ~n283) | (n282 & n284));
  assign n282 = x1 & x2;
  assign n283 = x2 ? (~x4 | x5) : (x4 | ~x5);
  assign n284 = x4 & x5;
  assign n285 = ~x0 & ~x3;
  assign n286 = n289 & (~n276 | (n287 & (x5 | n288)));
  assign n287 = (~x2 | x4) & (x0 | x2 | ~x4);
  assign n288 = (~x0 | ~x2 | ~x4 | x6) & (x0 | x2 | x4 | ~x6);
  assign n289 = (x1 | x2 | (~x0 & ~x3)) & (x0 | ~x1 | ~x2 | ~x3);
  assign z002 = n298 | (~x3 & (~n291 | ~n297)) | ~n302;
  assign n291 = (x1 | n292) & (~n295 | ~n296);
  assign n292 = (~x4 | n293) & (x0 | x2 | x4 | ~n294);
  assign n293 = (~x0 | x5 | ~x6 | (~x2 ^ ~x7)) & (x0 | ~x2 | ~x5 | x6 | ~x7);
  assign n294 = x7 & ~x5 & ~x6;
  assign n295 = ~x2 & ~x0 & x1;
  assign n296 = ~x7 & ~x6 & x4 & x5;
  assign n297 = (~x5 | ((x0 | (x1 ? (~x2 | ~x4) : (x2 | x4))) & (~x0 | x1 | ~x2 | ~x4))) & (x0 | x2 | ~x4 | x5);
  assign n298 = ~x3 & ((n300 & n301) | (~x2 & ~n299));
  assign n299 = (x0 | x1 | (x4 ? (~x5 | x6) : (x5 | ~x6))) & (x5 | x6 | ~x0 | ~x4);
  assign n300 = x2 & ~x0 & ~x1;
  assign n301 = x6 & x4 & x5;
  assign n302 = x2 ? (~x3 | (x0 & x1)) : (x3 | x4 | (~x0 & ~x1));
  assign z003 = n304 | n307 | n317 | (~n315 & ~n316);
  assign n304 = x0 & ((x4 & ~n305) | (~x1 & n306));
  assign n305 = (x1 | ((~x2 | (x3 ? (x5 | x6) : ~x5)) & (x3 | ~x5 | x6))) & (~x1 | x2 | x3 | x5 | ~x6);
  assign n306 = ~x4 & x2 & x3;
  assign n307 = x4 & (n309 | (n308 & n295 & n314));
  assign n308 = ~x6 & x7;
  assign n309 = ~x1 & ((n312 & n313) | (~n310 & ~n311));
  assign n310 = x3 ^ ~x7;
  assign n311 = (~x5 | x6 | x0 | ~x2) & (~x0 | x2 | x5 | ~x6);
  assign n312 = ~x3 & x0 & x2;
  assign n313 = x7 & ~x5 & x6;
  assign n314 = ~x3 & x5;
  assign n315 = x0 ^ ~x2;
  assign n316 = x3 ? (x4 & (x5 | x6)) : (~x4 | ~x5 | (~x1 & ~x6));
  assign n317 = ~x0 & (n318 | n319 | (n272 & n320));
  assign n318 = ~x2 & ((x3 & (~x4 | ~x5)) | (x5 & x6 & ~x3 & x4));
  assign n319 = x6 & ~x5 & x4 & x2 & x3;
  assign n320 = ~x6 & x4 & x5;
  assign z004 = ~n347 | n337 | n333 | n322 | ~n323;
  assign n322 = ~x0 & x2 & (x1 ? (x4 & x5) : (~x4 & ~x5));
  assign n323 = ~n326 & n332 & (x5 | ~n324 | n325);
  assign n324 = x0 & x2;
  assign n325 = (x1 | ~x3 | ~x4 | ~x6) & (~x1 | x3 | x4 | x6);
  assign n326 = ~n331 & ((n328 & n330) | (n327 & n329));
  assign n327 = x5 & x6;
  assign n328 = ~x5 & ~x6;
  assign n329 = ~x0 & x4;
  assign n330 = x0 & ~x4;
  assign n331 = x1 & x2;
  assign n332 = (~x0 | ~x4 | (x1 & x2) | ~x5) & (x4 | x5 | x0 | ~x1);
  assign n333 = ~x2 & (n334 | (x0 & n273 & n276));
  assign n334 = n336 & (x1 ? n284 : n335);
  assign n335 = ~x4 & ~x5;
  assign n336 = ~x6 & ~x0 & x3;
  assign n337 = (n338 | (n344 & n345)) & n346;
  assign n338 = n343 & ((n340 & n342) | (n339 & n341));
  assign n339 = ~x2 & ~x3;
  assign n340 = x2 & x3;
  assign n341 = x4 & x7;
  assign n342 = ~x4 & ~x7;
  assign n343 = x0 & x6;
  assign n344 = ~x3 & ~x0 & ~x2;
  assign n345 = x7 & ~x4 & ~x6;
  assign n346 = ~x1 & ~x5;
  assign n347 = ~n349 & (x2 | n348);
  assign n348 = (x0 | x1 | x4 | (~x5 ^ x6)) & (~x0 | ~x1 | ~x4 | x5 | ~x6);
  assign n349 = ~n350 & ((~x1 & ~n351) | (n295 & n352));
  assign n350 = ~x4 ^ ~x7;
  assign n351 = (~x0 | x5 | ~x6 | (x2 ^ ~x3)) & (x0 | ~x2 | ~x5 | x6);
  assign n352 = ~x6 & ~x3 & x5;
  assign z005 = ~n355 | ~n360 | ~n370 | (~x1 & ~n354);
  assign n354 = (x0 | ((x3 | ~x5 | ~x6) & (x5 | x6 | x2 | ~x3))) & (~x5 | x6 | ~x0 | x3);
  assign n355 = (n357 | n358) & (~n328 | ~n356 | ~n359);
  assign n356 = ~x3 & x4;
  assign n357 = x1 ? (x3 | x4) : (~x3 | ~x4);
  assign n358 = x0 ? ((~x5 | x6) & (~x2 | x5 | ~x6)) : (~x5 | ~x6);
  assign n359 = ~x2 & ~x0 & ~x1;
  assign n360 = ~n365 & (~x5 | (~n361 & n362));
  assign n361 = ~x0 & x6 & (x1 ? (~x3 & x4) : (x3 & ~x4));
  assign n362 = x6 | (x3 ? (x4 | ~n363) : (~x4 | ~n364));
  assign n363 = x0 & ~x1;
  assign n364 = ~x2 & x0 & x1;
  assign n365 = n367 & (n368 | (~x5 & n366 & ~n369));
  assign n366 = ~x2 & ~x4;
  assign n367 = ~x0 & ~x6;
  assign n368 = (~x5 ^ x7) & (x1 ? (~x2 & ~x3) : x2);
  assign n369 = x1 ? (~x3 | x7) : (x3 | ~x7);
  assign n370 = (~x1 | n371) & (~x0 | x1 | ~x6 | n372);
  assign n371 = (~x5 | ((x0 | (~x3 & (~x2 | x6))) & (x2 | ~x3 | x6))) & (~x0 | x2 | x5 | ~x6);
  assign n372 = (x7 & (x5 | (~x2 & ~x3 & ~x4))) | (~x5 & ~x7) | (x2 & x3 & x4);
  assign z006 = ~n375 | n386 | (x1 ? ~n390 : ~n374);
  assign n374 = x0 ? ((~x2 | ~x3 | ~x6 | ~x7) & (x6 | x7 | x2 | x3)) : (x2 ? ((x6 | ~x7) & (~x3 | ~x6 | x7)) : (~x6 | (x3 & ~x7)));
  assign n375 = ~n376 & (x4 ? n381 : (~n324 | n385));
  assign n376 = n366 & (n378 | (~x7 & ~n377 & n380));
  assign n377 = x5 ^ ~x6;
  assign n378 = ~n379 & n363 & ~x3 & x7;
  assign n379 = ~x5 ^ ~x6;
  assign n380 = x3 & ~x0 & x1;
  assign n381 = (~n383 | n384) & (~x3 | ~n295 | ~n382);
  assign n382 = ~x6 & ~x7;
  assign n383 = x6 & x0 & ~x1;
  assign n384 = x2 ? (~x3 | x7) : (x3 | ~x7);
  assign n385 = (~x1 | x3 | ~x6) & (x1 | ~x3 | x6 | x7);
  assign n386 = ~n388 & ((n308 & n387) | (~x1 & ~n389));
  assign n387 = ~x0 & x1;
  assign n388 = x2 ^ ~x3;
  assign n389 = x0 ? (x6 ^ x7) : (~x6 | x7);
  assign n390 = (x0 | x6 | (x2 ^ (x3 | ~x7))) & (x2 | ~x6 | (~x0 & (x3 | x7)));
  assign z007 = n392 | n396 | ~n402 | (~x3 & ~n401);
  assign n392 = ~x4 & ((n394 & n395) | (~x2 & ~n393));
  assign n393 = (x1 | x3 | (x0 ? (x5 ^ x7) : (~x5 | x7))) & (x0 | ~x1 | ~x3 | ~x5 | x7);
  assign n394 = x2 & x0 & ~x1;
  assign n395 = x7 & x3 & ~x5;
  assign n396 = ~x4 & (n397 | (n308 & n295 & n400));
  assign n397 = ~x1 & ((n280 & n344) | n398);
  assign n398 = x5 & n399 & (x2 ? (x3 & x7) : (~x3 & ~x7));
  assign n399 = x0 & ~x6;
  assign n400 = x3 & ~x5;
  assign n401 = (~x0 | ((~x4 | ~x7 | x1 | x2) & (~x1 | ~x2 | x4 | x7))) & (x0 | x1 | x2 | ~x4 | x7);
  assign n402 = n406 & n407 & (n405 | (~n403 & ~n404));
  assign n403 = ~x3 & x7;
  assign n404 = ~x7 & x3 & x4;
  assign n405 = x0 ? (x1 | ~x2) : (~x1 | x2);
  assign n406 = (x0 | ~x2 | (~x1 ^ x7)) & (~x0 | ~x1 | x2 | x7);
  assign n407 = (~n410 | ~n411) & (~x3 | ~n408 | n409);
  assign n408 = ~x1 & ~x2;
  assign n409 = ~x0 ^ ~x7;
  assign n410 = ~x3 & x2 & x0 & x1;
  assign n411 = ~x7 & ~x6 & x4 & ~x5;
  assign z008 = ~n416 | (~x1 & ((n413 & n411) | n414));
  assign n413 = x3 & ~x0 & x2;
  assign n414 = ~x4 & ((n294 & n344) | (x5 & ~n415));
  assign n415 = (x0 | x2 | x3 | ~x6 | x7) & (~x0 | ~x7 | (x2 ? (~x3 | ~x6) : (x3 | x6)));
  assign n416 = n419 & (~n408 | n417) & (~x3 | n418);
  assign n417 = (~x5 | ((~x0 | (x3 ? (~x4 | x6) : (x4 | ~x6))) & (x0 | x3 | x4 | x6))) & (x0 | x3 | x4 | x5 | ~x6);
  assign n418 = (x1 | (x0 ? (x2 ^ x4) : (~x2 | x4))) & (x2 | ~x4 | x0 | ~x1);
  assign n419 = ~n422 & (x3 | (n420 & n421)) & n427;
  assign n420 = x0 ? (~x1 | x2) : (x1 | ~x2);
  assign n421 = (~x2 | x4 | x0 | ~x1) & (~x0 | x1 | x2 | ~x4);
  assign n422 = n387 & ((n423 & n424) | (n425 & n426));
  assign n423 = ~x2 & x3;
  assign n424 = ~x4 & x5;
  assign n425 = x4 & ~x5;
  assign n426 = x2 & ~x3;
  assign n427 = (~n428 | ~n429) & (~n423 | ~n387 | ~n430);
  assign n428 = ~x2 & x0 & ~x1;
  assign n429 = ~x5 & x3 & x4;
  assign n430 = x7 & x6 & ~x4 & ~x5;
  assign z009 = ~n447 | ~n439 | ~n434 | n432 | n433;
  assign n432 = ~x4 & (x1 ? (x3 & (~x0 ^ ~x2)) : (x2 & ~x3));
  assign n433 = ~x1 & x4 & ((~x2 & ~x3) | (x0 & x2 & x3));
  assign n434 = ~n437 & (x2 | ~x5 | n435 | n436);
  assign n435 = x0 ? (x1 | ~x6) : (~x1 | x6);
  assign n436 = ~x3 ^ ~x4;
  assign n437 = n438 & n425 & (x0 ? (~x3 & ~x6) : (x3 & x6));
  assign n438 = ~x1 & x2;
  assign n439 = ~n440 & (x2 | n442);
  assign n440 = n441 & ((~x2 & x3 & ~x4 & ~x5) | (x2 & x4 & (x3 ^ ~x5)));
  assign n441 = ~x0 & ~x1;
  assign n442 = x5 ? (n444 | n445) : (~n443 | n446);
  assign n443 = x3 & ~x4;
  assign n444 = x0 ^ ~x6;
  assign n445 = (~x1 | ~x3 | ~x4 | x7) & (x1 | x3 | x4 | ~x7);
  assign n446 = (x0 | ~x1 | ~x6 | ~x7) & (~x0 | x1 | x6 | x7);
  assign n447 = x1 ? n448 : (~x2 | (~n449 & ~n452));
  assign n448 = (x0 | ~x5 | (x2 ? (x3 | ~x4) : (~x3 | x4))) & (x2 | x5 | (x3 ^ x4));
  assign n449 = n343 & (n451 | (n356 & n450));
  assign n450 = ~x5 & ~x7;
  assign n451 = x7 & x5 & x3 & ~x4;
  assign n452 = ~n453 & ~x6 & n329;
  assign n453 = x3 ? (x5 | ~x7) : (~x5 | x7);
  assign z010 = ~n471 | ~n462 | n455 | n459;
  assign n455 = x2 & ((n457 & n458) | (~x0 & ~n456));
  assign n456 = (x1 | ((x3 | ~x5 | (x4 ^ x6)) & (~x3 | ~x4 | x5 | ~x6))) & (~x3 | x6 | ((x4 | x5) & (~x1 | ~x4 | ~x5)));
  assign n457 = ~x3 & x0 & x1;
  assign n458 = ~x6 & ~x4 & ~x5;
  assign n459 = ~x2 & (x0 ? ~n461 : ~n460);
  assign n460 = (x1 | ~x3 | ~x4 | x5 | x6) & (~x1 | x3 | x4 | ~x5 | ~x6);
  assign n461 = x4 ? (x3 ? (~x5 | ~x6) : (x5 | x6)) : ((x1 | ~x6 | (~x3 ^ x5)) & (~x1 | ~x3 | ~x5 | x6));
  assign n462 = ~n463 & ~n466 & (x4 | n469 | n470);
  assign n463 = n329 & ((~x2 & n465) | (~x1 & x2 & n464));
  assign n464 = x3 & x5;
  assign n465 = ~x3 & ~x5;
  assign n466 = ~n467 & ((n278 & n387) | (x0 & ~n468));
  assign n467 = x3 ^ ~x5;
  assign n468 = x1 ? (x2 | x4) : (~x2 | ~x4);
  assign n469 = x2 ? (x3 | x5) : (~x3 | ~x5);
  assign n470 = x0 & x1;
  assign n471 = (~x3 & n472) | (~n479 & ~n482 & x3 & ~n477);
  assign n472 = (n474 | n475) & (~x5 | ~n473 | n476);
  assign n473 = ~x1 & ~x4;
  assign n474 = x0 ? (x5 | ~x6) : (~x5 | x6);
  assign n475 = (~x1 | ~x2 | x4 | x7) & (x1 | ~x4 | (~x2 ^ ~x7));
  assign n476 = (~x0 | x2 | x6 | ~x7) & (x0 | ~x6 | (~x2 ^ x7));
  assign n477 = ~n478 & ((n363 & n458) | (n387 & n301));
  assign n478 = x2 ^ ~x7;
  assign n479 = ~n481 & (x2 ? (~x5 & n441) : (x5 & n480));
  assign n480 = x0 & x1;
  assign n481 = x4 ? (x6 | ~x7) : (~x6 | x7);
  assign n482 = ~n485 & ((n483 & n363) | (n387 & n484));
  assign n483 = x2 & x5;
  assign n484 = ~x2 & ~x5;
  assign n485 = x4 ? (x6 | x7) : (~x6 | ~x7);
  assign z011 = ~n491 | (~n487 & (~n489 | (x1 & ~n488)));
  assign n487 = ~x3 ^ ~x7;
  assign n488 = (x2 | ((~x0 | ~x5 | (~x4 ^ x6)) & (x0 | x4 | x5 | ~x6))) & (x0 | ~x2 | ~x4 | ~x5 | ~x6);
  assign n489 = (~n273 | ~n300) & (n379 | n490);
  assign n490 = (x2 | ~x4 | x0 | ~x1) & (~x0 | x1 | ~x2 | x4);
  assign n491 = ~n492 & n497 & n508 & (~n408 | n496);
  assign n492 = n493 & (x0 ? ~n495 : (n276 & n494));
  assign n493 = x2 & x7;
  assign n494 = x6 & ~x4 & x5;
  assign n495 = (~x1 | x3 | x4 | x5 | ~x6) & (x1 | ~x4 | (x3 ? (~x5 | x6) : (x5 | ~x6)));
  assign n496 = (x3 | (((x4 ^ x5) | (x0 ^ ~x6)) & (~x5 | ~x6 | ~x0 | x4))) & (x0 | ~x3 | x4 | ~x5 | x6);
  assign n497 = ~n500 & n502 & n505 & (n498 | n499);
  assign n498 = ~x3 ^ ~x5;
  assign n499 = (x0 | x4 | x6 | (x1 ^ ~x2)) & (~x0 | ~x1 | x2 | ~x4 | ~x6);
  assign n500 = n387 & n501 & (x3 ? (~x4 ^ ~x6) : (~x4 & ~x6));
  assign n501 = x2 & ~x5;
  assign n502 = (~x4 | ((x6 | n504) & (x0 | ~x6 | n503))) & (x4 | ~x6 | n504) & (~x0 | x6 | n503);
  assign n503 = (x3 | ~x5 | x1 | ~x2) & (~x1 | x2 | ~x3 | x5);
  assign n504 = (x3 | ~x5 | x0 | ~x1) & (~x0 | x1 | ~x3 | x5);
  assign n505 = (~x0 | ~x5 | n325) & (x5 | n506 | ~n507);
  assign n506 = ~x3 ^ ~x6;
  assign n507 = x4 & ~x0 & ~x1;
  assign n508 = ~n511 & (n509 | n510);
  assign n509 = (x5 | ((~x1 | x7 | (~x3 ^ ~x6)) & (x1 | ~x3 | x6 | ~x7))) & (x1 | ~x5 | x6 | (~x3 ^ x7));
  assign n510 = x0 ? (x2 | x4) : (~x2 | ~x4);
  assign n511 = ~n310 & ((n512 & n514) | (n408 & ~n513));
  assign n512 = ~x6 & ~x4 & x5;
  assign n513 = (~x4 | (x0 ? (x5 | ~x6) : (~x5 | x6))) & (x0 | x4 | (x5 ^ x6));
  assign n514 = x2 & ~x0 & x1;
  assign z012 = ~n529 | ~n536 | (x1 ? ~n516 : ~n523);
  assign n516 = x4 ? n520 : (~n518 & (x3 | n517));
  assign n517 = x0 ? ((~x5 | x6 | x7) & (~x6 | ~x7 | ~x2 | x5)) : ((~x2 | ~x5 | x6 | ~x7) & (x2 | x5 | (x6 ^ x7)));
  assign n518 = n519 & ((x5 & ~x7 & ~x0 & x2) | (~x2 & x7 & (x0 | ~x5)));
  assign n519 = x3 & x6;
  assign n520 = x5 ? n522 : (~n521 | ~n344);
  assign n521 = x6 & ~x7;
  assign n522 = x0 ? (x2 | ((x6 | ~x7) & (x3 | ~x6 | x7))) : (~x2 | ((x6 | x7) & (~x3 | ~x6 | ~x7)));
  assign n523 = x0 ? (~n528 & (~x4 | n527)) : n524;
  assign n524 = (~x5 | n525) & (~x2 | ~n526);
  assign n525 = (x2 | ~x3 | x7 | (x4 ^ x6)) & (~x7 | ((~x4 | x6) & (~x2 | x3 | x4 | ~x6)));
  assign n526 = ~x5 & x7 & ((~x4 & x6) | (x3 & x4 & ~x6));
  assign n527 = x2 ? (~x7 | (x3 ? (~x5 | x6) : (x5 | ~x6))) : (x6 | x7 | (x3 ^ ~x5));
  assign n528 = n335 & ((~x3 & x6 & ~x7) | (~x2 & ((x6 & ~x7) | (x3 & ~x6 & x7))));
  assign n529 = ~n530 & (n534 | n535) & (n379 | n533);
  assign n530 = ~x2 & (x1 ? ~n531 : ~n532);
  assign n531 = x0 ? (x5 | (x3 ? (x4 | x6) : (~x4 | ~x6))) : (~x5 | ((~x4 | x6) & (x3 | x4 | ~x6)));
  assign n532 = (x0 | ((~x4 | x5 | ~x6) & (~x5 | x6 | x3 | x4))) & (~x0 | ~x3 | ~x4 | ~x5 | ~x6);
  assign n533 = (~x0 | x3 | (x1 ? (~x2 | x4) : (x2 | ~x4))) & (x0 | x1 | ~x2 | ~x3 | x4);
  assign n534 = x4 ? (x5 | ~x6) : (~x5 | x6);
  assign n535 = x0 ? (x2 | (x1 ? (~x3 | x7) : ~x7)) : (~x2 | (x1 ? (~x3 | ~x7) : x7));
  assign n536 = ~n537 & (n379 | (x1 & n540) | (~x1 & n539));
  assign n537 = x2 & ((~x5 & ~n538) | (n363 & n512));
  assign n538 = (x0 | ((x4 | x6 | x1 | x3) & (~x1 | ((x4 | ~x6) & (~x3 | ~x4 | x6))))) & (~x0 | x1 | ~x3 | ~x4 | ~x6);
  assign n539 = x0 ? (~x2 | (~x4 ^ x7)) : (x2 | ((x4 | ~x7) & (x3 | ~x4 | x7)));
  assign n540 = (~x0 | x2 | x3 | x4 | ~x7) & (x0 | ((x2 | ((~x4 | ~x7) & (~x3 | x4 | x7))) & (x3 | ((~x4 | ~x7) & (~x2 | x4 | x7)))));
  assign z013 = ~n548 | (~n542 & (~n544 | (x1 & ~n543)));
  assign n542 = ~x6 ^ ~x7;
  assign n543 = (x0 | ~x2 | ~x3 | ~x4 | x5) & (x3 | ((x4 | (x0 ? (~x2 ^ x5) : (x2 | x5))) & (x0 | x2 | ~x4 | ~x5)));
  assign n544 = ~n545 & ~n546 & (~n359 | ~n547);
  assign n545 = ~x0 & ((~x1 & x2 & ~x5) | (x5 & (x1 ? (~x2 ^ ~x3) : (~x2 & ~x3))));
  assign n546 = x0 & ((~x2 & x3 & ~x5) | (~x1 & (~x2 ^ x5)));
  assign n547 = x5 & x3 & ~x4;
  assign n548 = ~n564 & n569 & (x3 ? n557 : n549);
  assign n549 = x1 ? (n554 & (x6 | n553)) : n550;
  assign n550 = x2 ? n552 : n551;
  assign n551 = (x0 | ~x4 | ~x5 | x6 | ~x7) & (~x0 | x4 | x5 | ~x6 | x7);
  assign n552 = x0 ? ((~x5 | ~x6 | x7) & (~x4 | x5 | x6 | ~x7)) : ((x5 | ~x6 | x7) & (x4 | ~x5 | x6 | ~x7));
  assign n553 = (x0 | x4 | ~x7 | (~x2 ^ ~x5)) & (~x0 | ~x2 | ~x4 | x5 | x7);
  assign n554 = (~x0 | x2 | x4 | n555) & (x0 | ~x4 | (x2 ? n555 : ~n556));
  assign n555 = x5 ? (x6 | ~x7) : (~x6 | x7);
  assign n556 = ~x7 & x5 & x6;
  assign n557 = ~n560 & ~n562 & (n558 | ~n559);
  assign n558 = (~x1 | x2 | x5 | ~x6 | x7) & (x1 | x6 | ~x7 | (x2 ^ x5));
  assign n559 = x0 & x4;
  assign n560 = ~n555 & ((n366 & n480) | (~x0 & ~n561));
  assign n561 = x1 ? (~x2 | ~x4) : (x2 | x4);
  assign n562 = ~n563 & ((n366 & n363) | (~x0 & ~n468));
  assign n563 = x5 ? (~x6 | x7) : (x6 | ~x7);
  assign n564 = ~n565 & (n568 | (~n566 & (n269 | n567)));
  assign n565 = x6 ^ ~x7;
  assign n566 = ~x0 ^ ~x5;
  assign n567 = x1 & (x2 ? (~x3 & ~x4) : (x3 & x4));
  assign n568 = n438 & (x0 ? (x3 & ~x5) : (x5 & (~x3 ^ ~x4)));
  assign n569 = n572 & (n570 | n571);
  assign n570 = ~x5 ^ ~x7;
  assign n571 = (x0 | ~x3 | (x1 ? (~x2 | x4) : (x2 | ~x4))) & (~x0 | ~x1 | x2 | x3 | ~x4);
  assign n572 = (~n363 | n573) & (x3 | n574 | ~n575);
  assign n573 = (~x2 | x3 | x4 | x5 | ~x7) & (x2 | ~x3 | ~x4 | ~x5 | x7);
  assign n574 = x4 ? (x5 | ~x7) : (~x5 | x7);
  assign n575 = ~x2 & ~x0 & x1;
  assign z014 = n610 | n603 | ~n596 | ~n577 | ~n586;
  assign n577 = n578 & (n584 | n585) & (n490 | n583);
  assign n578 = (n580 | n581) & (x3 | ~n579 | n582);
  assign n579 = ~x0 & ~x2;
  assign n580 = x3 ? (~x4 | x6) : (x4 | ~x6);
  assign n581 = (~x2 | x5 | x0 | ~x1) & (~x0 | x1 | x2 | ~x5);
  assign n582 = (x5 | ~x6 | x1 | ~x4) & (~x1 | x4 | ~x5 | x6);
  assign n583 = (x3 | ~x5 | ~x6 | ~x7) & (~x3 | x5 | x6 | x7);
  assign n584 = (x0 | x1 | ~x2 | x3) & (~x0 | ~x1 | x2 | ~x3);
  assign n585 = (~x4 | ~x5 | x6 | x7) & (x4 | x5 | ~x6 | ~x7);
  assign n586 = ~n589 & n591 & (~n587 | ~n588 | ~n394);
  assign n587 = ~x5 & x6;
  assign n588 = x3 & x4;
  assign n589 = n428 & n590;
  assign n590 = x6 & ~x3 & x4;
  assign n591 = (~n592 | ~n593) & (~n594 | ~n595);
  assign n592 = x3 & x2 & ~x0 & x1;
  assign n593 = x7 & x6 & x4 & ~x5;
  assign n594 = ~x3 & ~x2 & x0 & ~x1;
  assign n595 = ~x7 & ~x6 & ~x4 & x5;
  assign n596 = n597 & ~n600 & (n584 | n602);
  assign n597 = (n490 | n506) & (n598 | n599);
  assign n598 = x2 ? (x4 | ~x6) : (~x4 | x6);
  assign n599 = x0 ? (~x1 | x3) : (x1 | ~x3);
  assign n600 = n601 & (x3 ? (~x6 & n282) : (x6 & n408));
  assign n601 = ~x0 & ~x4;
  assign n602 = x4 ? (~x5 | ~x6) : (x5 | x6);
  assign n603 = ~n565 & (n604 | ~n608 | (~n510 & ~n607));
  assign n604 = ~n605 & ((n363 & n588) | (n387 & n606));
  assign n605 = ~x2 ^ ~x5;
  assign n606 = ~x3 & ~x4;
  assign n607 = x1 ^ ~x3;
  assign n608 = x0 | x1 | x2 | (~n443 & ~n609);
  assign n609 = x5 & ~x3 & x4;
  assign n610 = ~n542 & (~n611 | ~n615 | (~n584 & ~n614));
  assign n611 = (~n514 | ~n612) & (~n428 | ~n613);
  assign n612 = x5 & x3 & x4;
  assign n613 = ~x5 & ~x3 & ~x4;
  assign n614 = x4 ^ ~x5;
  assign n615 = (x0 | ~x1 | x2 | ~x3 | x4) & (~x0 | x1 | ~x2 | x3 | ~x4);
  assign z015 = n627 | ~n639 | (x0 ? ~n631 : ~n617);
  assign n617 = x5 ? (~n621 & ~n623) : (~n618 & ~n619);
  assign n618 = n606 & ((x1 & ~x2 & ~x6 & x7) | (~x1 & (x2 ? (~x6 ^ x7) : (x6 & ~x7))));
  assign n619 = x4 & n620 & (x2 ? (x6 & x7) : (~x6 ^ ~x7));
  assign n620 = x1 & x3;
  assign n621 = ~x1 & ((n426 & n622) | (n423 & n345));
  assign n622 = ~x7 & x4 & x6;
  assign n623 = n625 & ((n624 & n382) | (~x2 & n626));
  assign n624 = x2 & ~x4;
  assign n625 = x1 & ~x3;
  assign n626 = x4 & (~x6 ^ x7);
  assign n627 = x0 & ((~x1 & ~n630) | (n628 & n629));
  assign n628 = x3 & x1 & ~x2;
  assign n629 = x7 & x4 & ~x5;
  assign n630 = (x2 | ((~x3 | ~x4 | (~x5 ^ x7)) & (x5 | ~x7 | x3 | x4))) & (~x2 | ~x3 | x4 | ~x5 | x7);
  assign n631 = n636 & (x5 | (~n632 & (~n272 | ~n635)));
  assign n632 = x1 & ((n426 & n634) | (n423 & n633));
  assign n633 = x7 & ~x4 & x6;
  assign n634 = ~x7 & x4 & ~x6;
  assign n635 = ~x7 & ~x4 & ~x6;
  assign n636 = (n565 | n637) & (~x5 | ~n438 | n638);
  assign n637 = (~x1 | x2 | ~x3 | ~x4 | ~x5) & (x1 | x4 | (x2 ? (~x3 | x5) : (x3 | ~x5)));
  assign n638 = (~x3 | ~x4 | x6 | x7) & (x3 | x4 | ~x6 | ~x7);
  assign n639 = ~n640 & ~n644 & n646 & (n570 | n643);
  assign n640 = ~x0 & ((~x3 & ~n641) | (n423 & ~n642));
  assign n641 = (x1 | ~x2 | ~x7 | (x4 ^ ~x5)) & (x2 | x7 | ((x4 | ~x5) & (~x1 | ~x4 | x5)));
  assign n642 = (~x1 | ~x4 | ~x5 | x7) & (x1 | x4 | x5 | ~x7);
  assign n643 = (x0 | x3 | (x1 ? (~x2 | x4) : (x2 | ~x4))) & (~x3 | ((~x0 | (x1 ? (x2 | x4) : (~x2 | ~x4))) & (~x2 | ~x4 | x0 | ~x1)));
  assign n644 = ~n645 & ((~x1 & x4 & (x2 ^ ~x7)) | (~x4 & ((x1 & ~x2 & x7) | (x2 & ~x7))));
  assign n645 = x0 ^ ~x3;
  assign n646 = (~n514 | ~n649) & (~n647 | n648);
  assign n647 = x0 & ~x2;
  assign n648 = (x4 | ~x7 | x1 | ~x3) & (~x1 | x3 | ~x4 | x7);
  assign n649 = x7 & ~x3 & x4;
  assign z016 = ~n664 | ~n671 | (x1 ? ~n657 : ~n651);
  assign n651 = x2 ? n655 : (~n652 & (~n556 | ~n654));
  assign n652 = ~x5 & ((n285 & n345) | (x0 & ~n653));
  assign n653 = (~x6 | x7 | x3 | ~x4) & (~x3 | x4 | x6 | ~x7);
  assign n654 = ~x4 & ~x0 & ~x3;
  assign n655 = (x0 | (x3 ? (x4 | ~n280) : (~x4 | ~n656))) & (~x0 | ~x3 | ~x4 | ~n656);
  assign n656 = x7 & x5 & ~x6;
  assign n657 = (~x6 | n658) & (~x5 | x6 | n310 | ~n663);
  assign n658 = (~n659 | ~n660) & (~n661 | ~n662);
  assign n659 = ~x0 & x3;
  assign n660 = x4 & (x2 ? (~x5 & x7) : (x5 & ~x7));
  assign n661 = ~x3 & x0 & ~x2;
  assign n662 = ~x7 & ~x4 & ~x5;
  assign n663 = ~x4 & ~x0 & x2;
  assign n664 = n667 & (n485 | n666) & (x0 | n665);
  assign n665 = (~x3 | (x1 ? ((x4 | x5) & (~x2 | ~x4 | ~x5)) : (~x4 | x5))) & (x1 | x2 | x3 | ~x4 | ~x5);
  assign n666 = x0 ? ((x1 | ~x2 | x3 | ~x5) & (~x1 | x2 | ~x3 | x5)) : (x2 | (x1 ? (x3 | x5) : (~x3 | ~x5)));
  assign n667 = (n271 | ~n669) & (~x0 | (n670 & (n271 | n668)));
  assign n668 = x3 ? (x4 | ~x5) : (~x4 | x5);
  assign n669 = x5 & ~x4 & ~x0 & ~x3;
  assign n670 = (~x1 | ~x2 | x3 | x4 | x5) & (x1 | x2 | ~x3 | ~x4 | ~x5);
  assign n671 = x3 ? (~n680 & (x2 | n679)) : n672;
  assign n672 = ~n674 & n676 & (n673 | n675);
  assign n673 = x4 ? (x5 | x6) : (~x5 | ~x6);
  assign n674 = n579 & (x1 ? (x4 & n327) : (~x4 & ~n377));
  assign n675 = x0 ? (x1 | x2) : (~x1 | ~x2);
  assign n676 = (n677 | n678) & (~n394 | ~n458);
  assign n677 = ~x4 ^ ~x5;
  assign n678 = (~x0 | ~x1 | x2 | x6) & (x0 | x1 | ~x2 | ~x6);
  assign n679 = ((~x5 ^ x6) | (x0 ? (x1 | x4) : (~x1 | ~x4))) & (~x0 | ~x1 | ~x4 | ~x5 | ~x6) & (x0 | x1 | x4 | x5 | x6);
  assign n680 = n438 & ~n677 & (x0 ^ ~x6);
  assign z017 = ~n698 | (x5 ? ~n691 : ~n682);
  assign n682 = x1 ? n683 : (~n686 & (x3 | n690));
  assign n683 = x2 ? n684 : n685;
  assign n684 = (x0 | ~x3 | ~x4 | ~x6 | ~x7) & (~x0 | x3 | x4 | x6 | x7);
  assign n685 = x6 ? ((x3 | x4 | ~x7) & (~x0 | ((x4 | ~x7) & (x3 | ~x4 | x7)))) : ((x0 | ((x4 | x7) & (x3 | ~x4 | ~x7))) & (~x3 | ((~x0 | ~x4 | ~x7) & (x4 | x7))));
  assign n686 = ~n688 & (n689 | (~x0 & ~n687));
  assign n687 = x2 ? (~x3 | ~x6) : (x3 | x6);
  assign n688 = x4 ^ ~x7;
  assign n689 = ~x6 & x3 & x0 & ~x2;
  assign n690 = (x0 | ~x2 | ~x4 | ~x6 | x7) & (~x0 | x2 | (x4 ? (x6 ^ x7) : (~x6 | x7)));
  assign n691 = ~n692 & ~n695 & (n350 | n694);
  assign n692 = x3 & ((n428 & n622) | (~x0 & ~n693));
  assign n693 = (~x1 | ~x2 | x4 | x6 | ~x7) & (x1 | x2 | (x4 ? (~x6 ^ x7) : (~x6 | ~x7)));
  assign n694 = (x0 | ((x3 | x6 | x1 | ~x2) & (~x3 | ~x6 | ~x1 | x2))) & (~x0 | x1 | ~x2 | ~x3 | x6);
  assign n695 = ~x3 & ((~n688 & ~n696) | (x2 & ~n697));
  assign n696 = (~x0 | x1 | ~x2 | ~x6) & (x0 | (x1 ? (~x2 | x6) : (x2 | ~x6)));
  assign n697 = (~x0 | x1 | ~x4 | x6 | ~x7) & (~x1 | x4 | ~x6 | x7);
  assign n698 = ~n704 & (x5 | n699) & (n702 | n703);
  assign n699 = ~n701 & (~x3 | ~n700 | ~n359);
  assign n700 = x4 & ~x6;
  assign n701 = x2 & ((~x4 & ~x6 & ~x0 & x1) | (~x1 & ((x4 & ~x6) | (x0 & ~x4 & x6))));
  assign n702 = (x2 | ((~x3 | x5 | ~x6) & (~x0 | ((~x5 | ~x6) & (x3 | x5 | x6))))) & (x0 | ((x3 | x5 | ~x6) & (~x2 | ~x3 | ~x5 | x6)));
  assign n703 = ~x1 ^ ~x4;
  assign n704 = x5 & (x0 ? ~n705 : ~n706);
  assign n705 = (x1 | ~x2 | ~x3 | ~x4 | ~x6) & (x6 | (x1 ? ((x2 & x3) | x4) : (x2 | ~x4)));
  assign n706 = (~x4 | ((~x1 | x2 | x3 | ~x6) & (x1 | (x2 ? ~x6 : (x3 | x6))))) & (~x1 | x4 | (x2 ? (~x3 | ~x6) : x6));
  assign z018 = ~n715 | (~x1 & (n708 | n712));
  assign n708 = x4 & ((n709 & ~n711) | (x3 & ~n710));
  assign n709 = ~x3 & x6;
  assign n710 = (~x6 | ((~x0 | x7 | (x2 ^ x5)) & (x0 | x2 | ~x5 | ~x7))) & (x0 | x5 | x6 | (~x2 ^ ~x7));
  assign n711 = (~x5 | x7 | x0 | ~x2) & (~x0 | ~x7 | (x2 ^ x5));
  assign n712 = n713 & n714;
  assign n713 = x3 & x0 & ~x2;
  assign n714 = ~x7 & x6 & ~x4 & x5;
  assign n715 = ~n716 & ~n727 & n732 & (n542 | n721);
  assign n716 = n718 & (x5 ? (n717 & n720) : ~n719);
  assign n717 = x6 & x7;
  assign n718 = x1 & ~x4;
  assign n719 = (~x6 | (x0 ? (x2 ? (x3 | x7) : (~x3 | ~x7)) : (x2 ? (~x3 | x7) : (x3 | ~x7)))) & (x0 | x2 | ~x3 | x6 | ~x7);
  assign n720 = ~x3 & ~x0 & x2;
  assign n721 = ~n723 & ~n724 & n726 & (~x0 | n722);
  assign n722 = (~x1 | x2 | x3 | ~x4 | x5) & (x1 | ((~x4 | ~x5 | x2 | x3) & (~x2 | ~x3 | x5)));
  assign n723 = ~x3 & ((~x0 & x2 & x4 & ~x5) | (x0 & ~x4 & (x2 ^ ~x5)));
  assign n724 = ~x0 & ((n725 & n612) | (n438 & n613));
  assign n725 = x1 & ~x2;
  assign n726 = (x0 | (x2 ? (~x3 | x5) : (x3 | ~x5))) & (x2 | ~x3 | ~x5 | (~x0 & x4));
  assign n727 = x2 & (n729 | (~n555 & (n363 | n728)));
  assign n728 = ~x3 & ~x0 & x1;
  assign n729 = n730 & ((n521 & n620) | (~x1 & ~n731));
  assign n730 = ~x0 & x5;
  assign n731 = x3 ? (~x6 | x7) : (x6 | ~x7);
  assign n732 = ~n735 & (x2 | (x0 & n734) | (~x0 & n733));
  assign n733 = x3 ? ((x5 | ~x6 | x7) & (x6 | ~x7 | x1 | ~x5)) : ((x5 | x6 | ~x7) & (~x6 | x7 | ~x1 | ~x5));
  assign n734 = x5 ? (~x6 | x7 | (~x1 & x3)) : (x6 | ~x7 | (x1 & ~x3));
  assign n735 = ~n736 & (x0 ? (n294 & n625) : ~n737);
  assign n736 = x2 ^ ~x4;
  assign n737 = (~x1 | ~x3 | ~x5 | x6 | ~x7) & (x1 | x3 | x5 | ~x6 | x7);
  assign z019 = ~n747 | n739 | n743;
  assign n739 = ~x3 & ((n411 & n742) | (n740 & ~n741));
  assign n740 = ~x2 & x6;
  assign n741 = (x5 | ((x0 | x1 | x4 | x7) & (~x0 | ~x7 | (x1 ^ x4)))) & (x0 | ~x5 | (x1 ? (x4 | x7) : (~x4 | ~x7)));
  assign n742 = x2 & x0 & x1;
  assign n743 = ~n506 & ((~x0 & ~n745) | (n744 & ~n746));
  assign n744 = x0 & ~x7;
  assign n745 = (~x1 | ~x2 | x4 | x5 | x7) & (~x7 | (x1 ^ (x4 & (~x2 | x5))));
  assign n746 = (x1 & (x2 | (~x4 & ~x5))) | (x4 & (x2 ? x5 : ~x1));
  assign n747 = ~n748 & n752 & n758 & (n750 | n751);
  assign n748 = ~n749 & ~x6 & n340;
  assign n749 = (x1 | (x0 ? (~x7 | (x4 ^ ~x5)) : (~x5 | x7))) & (~x5 | x7 | x0 | ~x4);
  assign n750 = (x0 | ~x2 | ~x3 | x5 | x6) & (~x0 | x2 | x3 | ~x5 | ~x6);
  assign n751 = x1 ? (x4 | ~x7) : (~x4 | x7);
  assign n752 = n756 & (n753 | n755) & (~n441 | ~n754);
  assign n753 = x3 ? (~x5 | x6) : (x5 | ~x6);
  assign n754 = x4 & x5 & (x3 ^ ~x6);
  assign n755 = x0 ? (x1 | ~x4) : (~x1 | x4);
  assign n756 = (~n457 | ~n458) & (~n300 | ~n757);
  assign n757 = ~x6 & ~x5 & x3 & ~x4;
  assign n758 = ~n759 & ~n767 & n769 & (x2 | n763);
  assign n759 = ~n761 & ((n363 & n760) | (~x0 & n762));
  assign n760 = ~x4 & x7;
  assign n761 = x2 ? (x3 | ~x6) : (~x3 | x6);
  assign n762 = ~x7 & (x1 ^ ~x4);
  assign n763 = (~n764 | ~n765) & (~x6 | ~n480 | n766);
  assign n764 = ~x6 & x4 & ~x5;
  assign n765 = ~x3 & ~x0 & ~x1;
  assign n766 = x3 ? (x4 | x5) : (~x4 | ~x5);
  assign n767 = ~n768 & x4 & n725;
  assign n768 = (x0 | x3 | ~x6 | x7) & (~x0 | ~x3 | x6 | ~x7);
  assign n769 = (n675 | n772) & (n770 | n771);
  assign n770 = x1 ? (x4 | x6) : (~x4 | ~x6);
  assign n771 = (x0 | x2 | ~x3 | x5) & (~x0 | ~x2 | x3 | ~x5);
  assign n772 = (~x3 | ~x4 | x5 | x6) & (x3 | x4 | ~x5 | ~x6);
  assign z020 = ~n780 | (~x3 & ~n774) | (x4 & ~n777);
  assign n774 = ~n775 & (n581 | (~n635 & (~x4 | n565)));
  assign n775 = ~x0 & (x1 ? (n366 & n656) : ~n776);
  assign n776 = (x6 | ((x2 | ~x5 | (~x4 ^ ~x7)) & (~x2 | ~x4 | x5 | x7))) & (x2 | x4 | ~x6 | (x5 ^ x7));
  assign n777 = (x2 | n778) & (~x2 | ~x3 | x5 | n779);
  assign n778 = (~x5 | (x1 ? (x7 | (x0 & ~x3)) : (~x3 | ~x7))) & (~x0 | ~x1 | x5 | x7);
  assign n779 = (x1 | x7) & (x0 | ~x1 | ~x7);
  assign n780 = n781 & (n791 | n792) & (x4 | n785);
  assign n781 = (n605 | n783) & (~x3 | ~n782 | n784);
  assign n782 = ~x0 & x2;
  assign n783 = x1 ? ((x3 | x4 | ~x7) & (x0 | (~x4 ^ x7))) : (x4 ? ~x7 : (x7 | (~x0 & ~x3)));
  assign n784 = (~x1 | x4 | x5 | ~x6 | ~x7) & (x1 | x6 | (x4 ? (~x5 | x7) : (x5 | ~x7)));
  assign n785 = ~n787 & ~n788 & (~x3 | ~n295 | ~n786);
  assign n786 = x5 & x7;
  assign n787 = ~n310 & ~n581;
  assign n788 = ~n388 & ((n790 & n441) | (n789 & n480));
  assign n789 = ~x5 & x7;
  assign n790 = x5 & ~x7;
  assign n791 = x1 ? (x2 | ~x5) : (~x2 | x5);
  assign n792 = (x3 | ~x6 | (x4 ^ x7)) & (~x0 | x6 | (x3 ? (x4 | ~x7) : (~x4 | x7)));
  assign z021 = x1 ? (n801 | ~n804) : ~n794;
  assign n794 = x5 ? (x3 ? n795 : n796) : n797;
  assign n795 = (~x0 | (x2 & (x4 | ~x6 | ~x7))) & (x0 | ~x2 | ~x4 | x6 | x7) & (x2 | (x4 & ~x6 & ~x7));
  assign n796 = x2 ? ((~x6 & (x4 | ~x7)) | (~x0 & (~x6 | (x4 & ~x7)))) : ((x6 & (~x4 | x7)) | (x0 & (x6 | (~x4 & x7))));
  assign n797 = ~n798 & ~n799 & n800 & (~n633 | ~n713);
  assign n798 = ~x4 & ((x2 & ~x7 & (x3 ^ ~x6)) | (~x2 & ~x3 & ~x6 & x7));
  assign n799 = x2 & x4 & (x3 ^ ~x6);
  assign n800 = x2 ? (~x3 | x6) : (x3 | ~x6);
  assign n801 = ~x3 & ((x5 & ~n802) | (n328 & ~n803));
  assign n802 = (x0 | ~x4 | ~x6 | (~x2 ^ ~x7)) & (x4 | x6 | ((~x2 | ~x7) & (~x0 | x2 | x7)));
  assign n803 = x2 ? (x7 | (~x0 ^ ~x4)) : (x4 | ~x7);
  assign n804 = ~n806 & n808 & (~x6 | ~n443 | n805);
  assign n805 = (x0 | ~x2 | x5 | x7) & (x2 | ((x5 | ~x7) & (~x0 | ~x5 | x7)));
  assign n806 = ~x0 & ((x2 & n807) | (~n283 & ~n506));
  assign n807 = ~x6 & x3 & ~x5;
  assign n808 = (~x2 | x3 | x4 | ~x5 | ~x6) & (x2 | ((x3 | x5 | ~x6) & (~x5 | ((~x4 | x6) & (~x3 | (~x4 & x6))))));
  assign z022 = n815 | (x5 ? ~n818 : ~n810);
  assign n810 = x0 ? (x1 ? n811 : n812) : n813;
  assign n811 = (x4 | ((x2 | ~x3 | x6) & (~x6 | ~x7 | ~x2 | x3))) & (x6 | x7 | x3 | ~x4) & (x2 | (x3 ? (~x6 | (~x4 & x7)) : (~x4 | x6)));
  assign n812 = (~x4 | (~x3 ^ ~x6)) & (~x3 | ((~x6 | x7) & (x4 | x6 | ~x7)));
  assign n813 = (~x3 | ((x4 | n814) & (~x6 | ~n408))) & (~x4 | (~x3 ^ ~x6));
  assign n814 = x7 ? x6 : (~x6 | (~x1 & ~x2));
  assign n815 = ~n542 & (~n817 | (n606 & ~n816));
  assign n816 = (~x0 | (x1 ? (x2 | x5) : (~x2 | ~x5))) & (x0 | x1 | ~x2 | x5);
  assign n817 = (x0 | x1 | ~x3 | ~x4 | ~x5) & (x3 | x4 | (x0 ? (~x1 ^ ~x5) : (~x1 | x5)));
  assign n818 = ~n819 & ~n821 & n824 & (n565 | n823);
  assign n819 = ~n487 & ~n820;
  assign n820 = (~x0 | x1 | x2 | x4 | x6) & (x0 | ~x1 | ((~x4 | ~x6) & (~x2 | x4 | x6)));
  assign n821 = n387 & ((n339 & n700) | (x2 & ~n822));
  assign n822 = x3 ? (x4 | ~x6) : (~x4 | x6);
  assign n823 = (x0 | x1 | x3 | ~x4) & (~x0 | ~x3 | x4 | (x1 ^ ~x2));
  assign n824 = (~n428 | ~n825) & (n331 | n506 | n826);
  assign n825 = x6 & x3 & ~x4;
  assign n826 = ~x0 ^ ~x4;
  assign z023 = ~n830 | (~x2 & (n829 | (x3 & ~n828)));
  assign n828 = x0 ? ((~x1 | ~x4 | x5 | ~x7) & (~x5 | x7 | x1 | x4)) : ((x4 | ~x5 | ~x7) & (x1 | x7 | (x4 ^ x5)));
  assign n829 = n314 & ((x0 & ~x1 & ~x4 & ~x7) | (~x0 & ((~x4 & x7) | (~x1 & x4 & ~x7))));
  assign n830 = ~n831 & ~n835 & ~n840 & (n350 | n839);
  assign n831 = ~x7 & (n832 | (n387 & n834));
  assign n832 = ~x2 & ((n457 & n764) | (~x0 & ~n833));
  assign n833 = (x1 | x3 | x4 | x5 | ~x6) & (~x1 | ~x5 | (x4 ^ x6));
  assign n834 = x2 & x5 & (x4 ^ ~x6);
  assign n835 = ~n836 & (n838 | (x0 & ~n837));
  assign n836 = x4 ^ ~x6;
  assign n837 = (x1 | x2 | ~x5 | ~x7) & (~x1 | x5 | x7 | (x2 ^ ~x3));
  assign n838 = ~x0 & x7 & (x1 ? (x2 & x5) : (~x2 & ~x5));
  assign n839 = (x0 & x1 & (x2 | (x3 & ~x5))) | (~x1 & ~x2 & x5) | (~x0 & (x5 | (~x1 & ~x2)));
  assign n840 = n483 & ((n480 & n842) | (~x0 & n841));
  assign n841 = ~x1 & (~x4 ^ ~x7);
  assign n842 = ~x7 & ~x3 & ~x4;
  assign z024 = n850 | ~n852 | (x3 ? ~n849 : ~n844);
  assign n844 = x5 ? (~n480 | ~n848) : ((~n480 | ~n845) & ~n846);
  assign n845 = x6 & x2 & ~x4;
  assign n846 = ~n847 & ((n700 & n387) | (x0 & ~n770));
  assign n847 = ~x2 ^ ~x7;
  assign n848 = ~x6 & ~x7 & (~x2 ^ ~x4);
  assign n849 = x5 ? (~n382 | ~n364) : (n847 | n435);
  assign n850 = ~x2 & ((n441 & n851) | (n294 & n480));
  assign n851 = x6 & (~x5 ^ ~x7);
  assign n852 = n853 & (n435 | n855) & (~x6 | n854);
  assign n853 = (~x0 | x1 | x5 | x6) & (x0 | ~x5 | (~x1 ^ ~x6));
  assign n854 = (~x0 | ~x1 | x2 | x5) & (x0 | x1 | ~x2 | ~x5);
  assign n855 = x2 ? (x5 | x7) : (~x5 | ~x7);
  assign z025 = n858 | ~n861 | (~n860 & (~x0 | n857));
  assign n857 = x0 & x3;
  assign n858 = ~x3 & ((n359 & n634) | (x0 & ~n859));
  assign n859 = (~x1 | ~x6 | x7 | (x2 ^ ~x4)) & (x6 | (~x2 ^ ~x7) | (x1 ^ ~x4));
  assign n860 = (x1 | ~x2 | x6) & (x2 | (x1 ? (x6 ^ ~x7) : (~x6 | ~x7)));
  assign n861 = (~x3 | n864) & (~n606 | n862) & (x3 | n863);
  assign n862 = x5 ? (~n382 | ~n359) : (n847 | n435);
  assign n863 = (~x1 | ((x0 | ~x2 | ~x6) & (x6 | ~x7 | ~x0 | x2))) & (~x0 | x1 | (x2 ? (x6 | x7) : (~x6 | ~x7)));
  assign n864 = (x0 | ~x1 | ~x2 | ~x6) & (x6 | x7 | x1 | x2);
  assign z026 = ~n869 | (~x3 & (~n866 | (~x4 & ~n867)));
  assign n866 = (x0 | ~x1 | ~x2 | ~x4 | x7) & (~x0 | ((~x1 | x4 | (x2 ^ x7)) & (~x4 | ((x2 | ~x7) & (x1 | ~x2 | x7)))));
  assign n867 = (~n394 | ~n556) & (x6 | n847 | n868);
  assign n868 = x0 ? (x1 | ~x5) : (~x1 | x5);
  assign n869 = n871 & (~n606 | n870);
  assign n870 = (~x2 | ((x0 | ~x1 | ~x5 | x7) & (~x0 | x1 | x5 | ~x7))) & (~x0 | x1 | x2 | (x5 ^ x7));
  assign n871 = (x0 & (~x3 | (x1 & ~x7))) | (x2 & x7) | (~x7 & (~x2 | (x1 & ~x3)));
  assign z027 = x4 ? ~n873 : (~n880 | (~n878 & ~n879));
  assign n873 = x3 ? ((~n294 | ~n364) & n877) : n874;
  assign n874 = (~n359 | ~n875) & (~n742 | ~n876);
  assign n875 = x7 & x5 & x6;
  assign n876 = ~x7 & ~x5 & ~x6;
  assign n877 = x0 & x1 & (x2 | (~x5 & ~x6));
  assign n878 = ~x2 ^ ~x6;
  assign n879 = (~x0 | x1 | ~x3 | ~x5 | ~x7) & (x0 | ~x1 | x3 | x5 | x7);
  assign n880 = n883 & (n868 | n881) & (~n428 | ~n882);
  assign n881 = x2 ? (x3 | x6) : (~x3 | ~x6);
  assign n882 = ~x7 & ~x6 & ~x3 & x5;
  assign n883 = x3 ? (x0 | (x1 & ~x5)) : (~x0 | (~x1 & x5));
  assign z028 = ~n895 | (x0 ? ~n891 : (n885 | n888));
  assign n885 = x6 & ((n269 & n886) | (x7 & ~n887));
  assign n886 = ~x7 & ~x4 & x5;
  assign n887 = (x1 | x2 | ~x3 | ~x4 | ~x5) & (~x1 | ~x2 | x5 | (x3 ^ ~x4));
  assign n888 = n328 & ((n725 & n889) | (n438 & n890));
  assign n889 = x7 & x3 & ~x4;
  assign n890 = ~x7 & ~x3 & x4;
  assign n891 = x1 ? (x5 ? ~n892 : n894) : (~x5 | n893);
  assign n892 = ~x4 & x2 & ~x3;
  assign n893 = (~x2 | ~x3 | x4 | ~x6 | x7) & (x2 | x3 | ~x4 | x6 | ~x7);
  assign n894 = (~x4 | x6 | x7 | (x2 ^ ~x3)) & (~x2 | x3 | x4 | (~x6 & ~x7));
  assign n895 = ~n897 & n901 & n904 & (~n896 | ~n900);
  assign n896 = ~x5 & ~x4 & ~x0 & x1;
  assign n897 = ~x1 & ((n294 & n898) | (x5 & ~n899));
  assign n898 = x4 & ~x0 & x2;
  assign n899 = x0 ? ((~x2 | ~x4 | ~x6 | ~x7) & (x6 | x7 | x2 | x4)) : (x2 | ~x6 | (~x4 ^ x7));
  assign n900 = ~x7 & (x2 ^ ~x6);
  assign n901 = (n868 | n902) & (~n507 | n903);
  assign n902 = x2 ? (x4 | x6) : (~x4 | ~x6);
  assign n903 = x2 ? (x5 | ~x6) : (~x5 | x6);
  assign n904 = x0 ? (x4 | (x1 ? x2 : x5)) : (~x4 | ((~x5 | (~x1 & ~x2)) & (x1 | x2 | x5)));
  assign z029 = ~n917 | ~n925 | (x0 ? ~n911 : ~n906);
  assign n906 = x2 ? n907 : (~n909 & (~x5 | n908));
  assign n907 = (~x1 | x3 | x4 | ~n875) & (~x4 | ~n876 | x1 | ~x3);
  assign n908 = x1 ? (x4 | (x3 ? (~x6 | x7) : (x6 | ~x7))) : (~x4 | ~x6 | (~x3 ^ ~x7));
  assign n909 = n465 & ((n521 & n473) | (n308 & n910));
  assign n910 = x1 & x4;
  assign n911 = ~n912 & (x6 | ~n484 | n916);
  assign n912 = x5 & ((n913 & ~n914) | (n718 & ~n915));
  assign n913 = ~x1 & x4;
  assign n914 = (x6 | ~x7 | x2 | ~x3) & (~x2 | x3 | ~x6 | x7);
  assign n915 = (x2 | ~x3 | x6 | x7) & (~x2 | x3 | (~x6 & ~x7));
  assign n916 = (~x1 | ~x3 | ~x4 | x7) & (x1 | x4 | (~x3 ^ ~x7));
  assign n917 = ~n920 & (x3 ? (~n438 | n918) : n919);
  assign n918 = (x6 | ~x7 | x0 | ~x5) & (~x0 | ~x6 | (~x5 ^ x7));
  assign n919 = x0 ? ((x1 | ~x2 | x5 | ~x6) & (~x1 | x2 | ~x5 | x6)) : (~x5 | (x1 ? (x2 | ~x6) : (~x2 | x6)));
  assign n920 = ~x2 & (n922 | (x0 & n276 & n921));
  assign n921 = ~x7 & x5 & ~x6;
  assign n922 = n924 & ((n717 & n923) | (n382 & n625));
  assign n923 = ~x1 & x3;
  assign n924 = ~x0 & ~x5;
  assign n925 = n927 & (n444 | n926);
  assign n926 = x1 ? ((~x5 | ~x7 | x2 | ~x3) & (x5 | x7 | ~x2 | x3)) : (x2 | (x3 ? (~x5 | x7) : (x5 | ~x7)));
  assign n927 = ~n928 & ~n929 & (~n387 | ~n400 | n878);
  assign n928 = ~x1 & (x0 ? (x2 ? (x5 & ~x6) : (~x5 & x6)) : (x5 & (~x2 ^ x6)));
  assign n929 = x1 & ((x5 & x6 & x0 & ~x2) | (~x5 & ~x6 & ~x0 & x2));
  assign z030 = n937 | ~n939 | (~x0 & (n931 | ~n934));
  assign n931 = ~x3 & ((~x6 & ~n933) | (n932 & n280));
  assign n932 = x4 & ~x1 & ~x2;
  assign n933 = (x1 | x2 | x4 | x5 | ~x7) & (~x1 | ~x5 | (x2 ? (~x4 | ~x7) : (x4 | x7)));
  assign n934 = (~x7 | ((x6 | n935) & (~n923 | n936))) & (~x6 | x7 | n935);
  assign n935 = ((x4 & x5) | (x1 ? (~x2 | x3) : (x2 | ~x3))) & (x2 | ~x4 | ~x5 | (~x1 ^ ~x3));
  assign n936 = (~x5 | x6 | x2 | ~x4) & (~x2 | x4 | x5 | ~x6);
  assign n937 = ~x3 & ((n301 & n514) | (~x1 & ~n938));
  assign n938 = (x0 | x2 | x4 | ~x5 | x6) & (x5 | ((~x0 | (x2 ? (~x4 | x6) : (x4 | ~x6))) & (x0 | x2 | ~x4 | x6)));
  assign n939 = n942 & (n542 | (n941 & (x4 | n940)));
  assign n940 = (~x0 | x1 | x2 | x3 | ~x5) & (x0 | ((~x3 | ~x5 | x1 | ~x2) & (x3 | x5 | ~x1 | x2)));
  assign n941 = (x0 | x1 | ~x2 | ~x3 | ~x4) & (~x0 | (x1 ? (x2 ? (x3 | x4) : (~x3 | ~x4)) : (x2 | (~x3 ^ x4))));
  assign n942 = n945 & (~x0 | (~n944 & (~x1 | n943)));
  assign n943 = (x4 | ~n875 | x2 | ~x3) & (~x2 | x3 | ~x4 | ~n876);
  assign n944 = n438 & ~n565 & (x3 | n284);
  assign n945 = ~n947 & (~n423 | n946) & (x6 | n948);
  assign n946 = (~x0 | ~x1 | x4 | x5 | ~x6) & (x0 | ~x4 | (x1 ? (x5 | x6) : (~x5 | ~x6)));
  assign n947 = x6 & ((x0 & x1 & ~x2 & ~x3) | (~x0 & x2 & (x1 ^ ~x3)));
  assign n948 = x0 ? (x1 | (x2 ? (x3 | x4) : (~x3 | ~x4))) : (~x1 | x2 | (~x3 ^ x4));
  assign z031 = ~n950 | n959 | ~n963 | (n438 & ~n958);
  assign n950 = (n310 | n952) & (x2 | (n951 & n953));
  assign n951 = ((x4 ^ x7) | (x0 ? (x1 | ~x3) : (~x1 | x3))) & (x0 | ~x1 | ~x3 | x4 | ~x7) & (~x0 | x3 | (x1 ? (x4 | ~x7) : (~x4 | x7)));
  assign n952 = x0 ? (x1 ? (x2 | ~x4) : (~x2 | x4)) : (x1 | (x2 ^ x4));
  assign n953 = (n954 | n956) & (~n955 | n957);
  assign n954 = ~x1 ^ ~x3;
  assign n955 = ~x1 & ~x7;
  assign n956 = (~x5 | x7 | x0 | ~x4) & (~x0 | x4 | x5 | ~x7);
  assign n957 = (~x4 | x5 | x0 | ~x3) & (~x0 | x3 | x4 | ~x5);
  assign n958 = (x0 | ~x3 | x4 | ~x5 | x7) & (~x0 | x3 | ~x4 | (~x5 ^ x7));
  assign n959 = x2 & (n961 | (x4 & n625 & ~n960));
  assign n960 = (x0 | ~x5 | ~x6 | ~x7) & (~x0 | x5 | x6 | x7);
  assign n961 = n962 & n441 & x3 & ~x4;
  assign n962 = ~x5 & (~x6 ^ ~x7);
  assign n963 = x2 ? n964 : (~n965 & (x0 | n968));
  assign n964 = x1 ? ((x3 | x4 | x7) & (x0 | (x3 ^ x7))) : ((x0 | x3 | x4 | ~x7) & (~x4 | x7 | ~x0 | ~x3));
  assign n965 = ~n966 & ~n967;
  assign n966 = x3 ? (~x5 | ~x6) : (x5 | x6);
  assign n967 = (~x0 | ~x1 | x4 | x7) & (x0 | x1 | ~x4 | ~x7);
  assign n968 = (x1 | ~x4 | x7 | n753) & (~x1 | ~x7 | n772);
  assign z032 = n970 | ~n979 | (x1 & (n973 | n977));
  assign n970 = ~x3 & (x0 ? ~n972 : (n408 & n971));
  assign n971 = x6 & x4 & ~x5;
  assign n972 = (x1 | ~x2 | x4 | x5 | x6) & (x2 | ((~x5 | x6 | x1 | ~x4) & (~x1 | x5 | (~x4 ^ x6))));
  assign n973 = ~x0 & ((n974 & n875) | (~n975 & ~n976));
  assign n974 = ~x4 & ~x2 & ~x3;
  assign n975 = x4 ? (~x6 | ~x7) : (x6 | x7);
  assign n976 = x2 ? (x3 | ~x5) : (~x3 | x5);
  assign n977 = ~n978 & n647 & ~n498;
  assign n978 = x4 ? (~x6 | x7) : (x6 | ~x7);
  assign n979 = ~n980 & ~n985 & n988 & (x1 | n984);
  assign n980 = x3 & ((~x0 & ~n982) | (n981 & ~n983));
  assign n981 = x0 & x5;
  assign n982 = (~x1 | ~x2 | ~x4 | x5 | x6) & (x1 | ~x6 | (x2 ? (x4 | x5) : (~x4 | ~x5)));
  assign n983 = (x1 | ~x2 | x4 | x6) & (~x1 | x2 | (x4 ^ ~x6));
  assign n984 = ((~x0 ^ ~x2) | (x3 ? (x4 | x5) : (~x4 | ~x5))) & ((x3 ^ x5) | (x0 ? (x2 | ~x4) : (~x2 | x4)));
  assign n985 = n387 & (~n986 | ~n987);
  assign n986 = x2 ? (~x3 | x4) : (x3 | ~x4);
  assign n987 = (x2 | ~x3 | ~x4 | ~x5) & (~x2 | x3 | x4 | x5);
  assign n988 = (~n714 | ~n990) & (n989 | (~n300 & ~n647));
  assign n989 = x3 ? (~x4 | x5) : (x4 | ~x5);
  assign n990 = x3 & x2 & x0 & ~x1;
  assign z033 = n1002 | ~n1005 | (x5 ? ~n997 : ~n992);
  assign n992 = ~n993 & (~n300 | ~n996);
  assign n993 = ~x2 & (x0 ? ~n994 : ~n995);
  assign n994 = (x1 | ~x3 | x4 | ~x6 | x7) & (x3 | ((x6 | x7 | x1 | ~x4) & (~x1 | ~x7 | (x4 ^ x6))));
  assign n995 = (x1 | x3 | x4 | x6 | ~x7) & (~x3 | ((x6 | x7 | x1 | ~x4) & (~x1 | ~x7 | (x4 ^ x6))));
  assign n996 = ~x7 & x6 & ~x3 & ~x4;
  assign n997 = ~n999 & (n751 | (~n689 & (~n285 | n998)));
  assign n998 = x2 ^ ~x6;
  assign n999 = x6 & ((n364 & n1001) | (x2 & ~n1000));
  assign n1000 = (x1 | x4 | (x0 ? (x3 ^ x7) : (~x3 | x7))) & (x0 | ~x1 | ~x4 | (~x3 ^ x7));
  assign n1001 = x7 & x3 & x4;
  assign n1002 = ~x2 & (x0 ? ~n1003 : ~n1004);
  assign n1003 = x1 ? (x3 ? (x4 ? (x5 | x6) : (~x5 | ~x6)) : (x4 | (~x5 ^ x6))) : ((~x5 | ~x6 | x3 | ~x4) & (x5 | x6 | ~x3 | x4));
  assign n1004 = ((~x3 ^ ~x6) | (x1 ? (x4 | x5) : (~x4 | ~x5))) & (~x1 | ~x3 | x4 | ~x5 | x6) & (x1 | x3 | x5 | ~x6);
  assign n1005 = ~n1010 & ~n1013 & (~x2 | (~n1006 & n1007));
  assign n1006 = n285 & ((n328 & n473) | (x1 & ~n673));
  assign n1007 = (~n458 | ~n1008) & (n377 | n1009);
  assign n1008 = x3 & x0 & ~x1;
  assign n1009 = (~x0 | x1 | x3 | x4) & (x0 | ~x3 | (~x1 ^ ~x4));
  assign n1010 = ~n645 & (x1 ? ~n1012 : (x5 & ~n1011));
  assign n1011 = ~x2 ^ ~x4;
  assign n1012 = x2 ? (x4 | x5) : (~x4 | ~x5);
  assign n1013 = n425 & (n1014 | (~x1 & (n857 | n720)));
  assign n1014 = ~x3 & ~x2 & ~x0 & x1;
  assign z034 = n1017 | ~n1023 | ~n1032 | (~n1016 & ~n1031);
  assign n1016 = x1 ^ ~x4;
  assign n1017 = ~x2 & (n1018 | (n765 & n1022));
  assign n1018 = ~x5 & ((~n565 & ~n1020) | (n1019 & ~n1021));
  assign n1019 = ~x4 & ~x6;
  assign n1020 = (~x3 | x4 | x0 | ~x1) & (~x0 | x1 | x3 | ~x4);
  assign n1021 = (~x0 | ~x1 | x3 | ~x7) & (x0 | x1 | (x3 ^ ~x7));
  assign n1022 = x7 & x6 & x4 & x5;
  assign n1023 = ~n1027 & (n989 | n1026) & (n1024 | n1025);
  assign n1024 = x3 ? (x4 | x7) : (~x4 | ~x7);
  assign n1025 = (~x0 | ~x1 | x2 | x5 | ~x6) & (x0 | ~x2 | ~x5 | (~x1 ^ ~x6));
  assign n1026 = (x0 | x2 | ~x6 | (~x1 ^ ~x7)) & (~x0 | x1 | ~x2 | x6 | x7);
  assign n1027 = ~n688 & (n1030 | (~n1028 & ~n1029));
  assign n1028 = x0 ? (x2 | ~x3) : (~x2 | x3);
  assign n1029 = x1 ? (~x5 | x6) : (x5 | ~x6);
  assign n1030 = ~n645 & n438 & x5 & x6;
  assign n1031 = x2 ? ((x0 | (x3 ? x6 : (~x5 | ~x6))) & (x3 | x6 | (~x0 & x5))) : ((~x0 | ((~x5 | ~x6) & (~x3 | x5 | x6))) & (~x6 | ((~x3 | ~x5) & (x0 | x3 | x5))));
  assign n1032 = ~n1042 & ~n1040 & n1038 & ~n1033 & ~n1035;
  assign n1033 = ~n1034 & ~n903;
  assign n1034 = x0 ? (x1 | x4) : (~x1 | ~x4);
  assign n1035 = ~n1036 & (n1037 | (n624 & n441));
  assign n1036 = x3 ? (x5 | ~x6) : (~x5 | x6);
  assign n1037 = x4 & ~x2 & x0 & x1;
  assign n1038 = ~n1039 | ((~x3 | ~x4 | ~n394) & (x4 | ~n359));
  assign n1039 = x5 & ~x6;
  assign n1040 = ~n1041 & (x1 ? (~x3 & ~x7) : (x3 & x7));
  assign n1041 = (~x0 | ~x2 | x4 | ~x5 | ~x6) & (x0 | x2 | ~x4 | x5 | x6);
  assign n1042 = ~n1044 & (n1043 | (n588 & n786));
  assign n1043 = ~x7 & ~x5 & ~x3 & ~x4;
  assign n1044 = (x0 | ~x1 | ~x2 | ~x6) & (~x0 | x2 | (~x1 ^ ~x6));
  assign z035 = n1046 | ~n1049 | n1056 | (x2 & ~n1059);
  assign n1046 = ~x1 & (x2 ? ~n1047 : ~n1048);
  assign n1047 = (x0 | x3 | x4 | x5 | ~x7) & (~x0 | ~x3 | ~x4 | ~x5 | x7);
  assign n1048 = ((x0 ^ ~x3) | ((~x4 | x5 | ~x7) & (~x5 | x7))) & (x4 | ~x7 | (x0 ? (~x3 | x5) : (x3 | ~x5)));
  assign n1049 = n1053 & (x2 | (n1051 & (n1016 | n1050)));
  assign n1050 = (~x0 | ~x3 | ~x5 | x6 | ~x7) & (x0 | x3 | x5 | ~x6 | x7) & ((x0 ? (~x3 | x5) : (x3 | ~x5)) | (x6 ^ x7));
  assign n1051 = (x0 | x1 | x3 | ~n1052) & (~x0 | ~x1 | ~x3 | ~n593);
  assign n1052 = ~x4 & ~x7 & (~x5 ^ ~x6);
  assign n1053 = (n570 | n1054) & (~n725 | n1055);
  assign n1054 = (~x1 | ~x4 | (x0 ? (x2 | ~x3) : (~x2 | x3))) & (~x2 | (x1 & x4) | (x0 ^ ~x3));
  assign n1055 = (x0 | x3 | ~x4 | ~x5 | x7) & ((x0 ^ ~x3) | ((x5 | ~x7) & (x4 | ~x5 | x7)));
  assign n1056 = ~n379 & (n1058 | (~x1 & ~n1057));
  assign n1057 = (~x0 | ~x2 | ~x3 | ~x4 | ~x7) & (x4 | ((x2 | (x0 ? (~x3 ^ x7) : (~x3 | ~x7))) & (x0 | ~x2 | x3 | x7)));
  assign n1058 = x4 & n725 & (x0 ? (~x3 & ~x7) : (x3 ^ x7));
  assign n1059 = n1062 & (n310 | n1061) & (n542 | n1060);
  assign n1060 = (~x0 | x1 | ~x3 | x4 | ~x5) & (x0 | ((~x4 | x5 | x1 | x3) & (~x1 | (x3 ? (~x4 | ~x5) : (x4 | x5)))));
  assign n1061 = (~x0 | x1 | x4 | x5 | ~x6) & (x0 | ((~x1 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (x1 | ~x4 | ~x5 | x6)));
  assign n1062 = (~n430 | ~n1063) & (~n1039 | ~n1064 | ~n1065);
  assign n1063 = x3 & ~x0 & ~x1;
  assign n1064 = x0 & ~x3;
  assign n1065 = ~x7 & (~x1 ^ ~x4);
  assign z036 = n1067 | n1071 | ~n1076 | (~n350 & ~n1070);
  assign n1067 = x6 & ((~x7 & ~n1068) | (n760 & ~n1069));
  assign n1068 = (x2 | (((~x1 ^ x4) | (x0 ^ ~x3)) & (~x0 | ~x1 | ~x3 | ~x4))) & (~x4 | ((~x0 | x1 | ~x2 | ~x3) & (x0 | ~x1 | x3)));
  assign n1069 = x0 ? (~x1 | x3) : (x1 ? ~x3 : (x2 | x3));
  assign n1070 = (x0 | ~x1 | x2 | x3 | x6) & (x1 | (x0 ? (~x3 ^ x6) : ((~x3 | ~x6) & (~x2 | x3 | x6))));
  assign n1071 = ~x6 & (n1073 | n1075 | (~x2 & ~n1072));
  assign n1072 = (x0 | x1 | ~x3 | x4 | ~x7) & (~x0 | x7 | (x1 ? (x3 ^ ~x4) : (~x3 | ~x4)));
  assign n1073 = ~n954 & ((n647 & n760) | (~x0 & n1074));
  assign n1074 = x4 & ~x7;
  assign n1075 = ~x4 & ~x3 & x2 & ~x0 & x1;
  assign n1076 = x5 ? n1077 : (~n1083 & n1085);
  assign n1077 = n1080 & (x3 | (~n1079 & (x0 | n1078)));
  assign n1078 = (~x1 | x2 | x4 | x6 | ~x7) & (x1 | ~x2 | ~x4 | ~x6 | x7);
  assign n1079 = n324 & ((n382 & n718) | (~x1 & ~n485));
  assign n1080 = (n350 | n1081) & (~n923 | n1082);
  assign n1081 = (~x0 | ~x1 | x2 | ~x3 | ~x6) & (x0 | ((x3 | x6 | x1 | x2) & (~x1 | ~x2 | (~x3 ^ x6))));
  assign n1082 = x0 ? ((~x2 | x4 | x6 | ~x7) & (x2 | ~x4 | ~x6 | x7)) : (~x2 | (x4 ? (x6 | x7) : (~x6 | ~x7)));
  assign n1083 = x0 & ((n272 & n633) | (n700 & ~n1084));
  assign n1084 = (~x3 | x7 | x1 | ~x2) & (~x1 | (x2 ? (x3 | x7) : (~x3 | ~x7)));
  assign n1085 = x0 ? (x3 | n1086) : (x3 ? n1086 : (n847 | n1087));
  assign n1086 = (x1 | x4 | x6 | (~x2 ^ ~x7)) & (~x6 | ((~x1 | (x2 ? (x4 | x7) : (~x4 | ~x7))) & (x1 | ~x2 | ~x4 | x7)));
  assign n1087 = x1 ? (~x4 | x6) : (x4 | ~x6);
  assign z037 = n1095 | ~n1100 | (x3 ? ~n1097 : ~n1089);
  assign n1089 = x1 ? n1090 : (x0 ? n1094 : n1093);
  assign n1090 = (x7 | n1092) & (~n330 | n1091 | x6 | ~x7);
  assign n1091 = x2 ^ ~x5;
  assign n1092 = (x0 | ~x6 | (x2 ? (x4 | ~x5) : (~x4 | x5))) & (~x0 | ~x2 | ~x4 | x5 | x6);
  assign n1093 = (x2 | x4 | x5 | x6 | ~x7) & (~x2 | ~x4 | ~x5 | ~x6 | x7);
  assign n1094 = (~x2 | ~x4 | x5 | x6 | ~x7) & (x2 | ((~x4 | ~x5 | x6 | ~x7) & (~x6 | x7 | x4 | x5)));
  assign n1095 = ~n542 & (x3 ? (~n1091 & ~n1034) : ~n1096);
  assign n1096 = (x0 | x1 | ~x2 | x4 | ~x5) & (x2 | ((~x0 | ~x1 | ~x4 | ~x5) & (x0 | x5 | (~x1 ^ x4))));
  assign n1097 = (n1091 | n1098) & (~n366 | ~n521 | n1099);
  assign n1098 = (~x0 | x1 | ~x4 | ~x6 | x7) & (x0 | x6 | ~x7 | (x1 ^ ~x4));
  assign n1099 = x0 ? (~x1 | ~x5) : (x1 | x5);
  assign n1100 = ~n1101 & n1104 & (n688 | n1103);
  assign n1101 = ~x1 & ((n339 & n886) | (~n1024 & ~n1102));
  assign n1102 = x0 ? (x2 | x5) : (x2 ^ ~x5);
  assign n1103 = ((~x0 & ~x3) | (x1 ? (x2 | x5) : (~x2 | ~x5))) & (x0 | ~x1 | x3 | (~x2 ^ x5));
  assign n1104 = (n1105 | n1106) & (~n387 | ~n483 | n1107);
  assign n1105 = (x2 | ~x3 | ~x4 | ~x7) & (~x2 | x3 | x4 | x7);
  assign n1106 = (x1 | x5) & (~x0 | ~x1 | ~x5);
  assign n1107 = (~x4 | ~x7) & (~x3 | x4 | x7);
  assign z038 = n1109 | ~n1112 | n1126 | (n408 & ~n1129);
  assign n1109 = x1 & ((n296 & n413) | n1110);
  assign n1110 = x6 & ((n782 & ~n1111) | (x0 & ~n573));
  assign n1111 = (~x5 | x7 | x3 | ~x4) & (~x3 | x4 | x5 | ~x7);
  assign n1112 = n1118 & (x0 | (n1113 & n1115)) & n1123;
  assign n1113 = (~n301 | ~n628) & (~n1114 | ~n458);
  assign n1114 = ~x3 & ~x1 & x2;
  assign n1115 = (n534 | n1117) & (n836 | n1116);
  assign n1116 = (x1 | x2 | ~x3 | x5) & (~x1 | ~x2 | x3 | ~x5);
  assign n1117 = x1 ? (~x2 | ~x3) : (x2 | x3);
  assign n1118 = (n1119 | n1120) & (~n1121 | ~n1122);
  assign n1119 = x1 ? (x2 | x5) : (~x2 | ~x5);
  assign n1120 = x0 ? (x3 | x6) : (x3 ^ ~x6);
  assign n1121 = x6 & (~x2 ^ ~x5);
  assign n1122 = x3 & x0 & ~x1;
  assign n1123 = (n574 | n1124) & (n570 | n1016 | n1125);
  assign n1124 = (x0 | ~x1 | x2 | x3 | x6) & (x1 | ~x2 | (x0 ? (~x3 ^ x6) : (~x3 | ~x6)));
  assign n1125 = (x0 | ~x2 | x3 | x6) & (x2 | (x0 ? (x3 ^ ~x6) : (~x3 | ~x6)));
  assign n1126 = x0 & ((~x2 & ~n1128) | (n512 & n1127));
  assign n1127 = ~x3 & x1 & x2;
  assign n1128 = (~x1 | x3 | ~x4 | ~x5 | ~x6) & (x1 | ~x3 | x4 | x5 | x6) & ((x1 ? (~x3 | ~x5) : (x3 | x5)) | (~x4 ^ x6));
  assign n1129 = (~x0 | x3 | x4 | ~n294) & (x0 | (x3 ? (x4 | ~n294) : n585));
  assign z039 = n1134 | ~n1136 | ~n1140 | (x2 & ~n1131);
  assign n1131 = ~n1132 & (n565 | n1060) & (~n387 | n1133);
  assign n1132 = ~x1 & ~n481 & (x0 ? n400 : n314);
  assign n1133 = (~x3 | ~x4 | x5 | ~x6 | x7) & (x3 | x4 | ~x5 | x6 | ~x7);
  assign n1134 = ~n542 & (n1135 | (x5 & n910 & ~n1028));
  assign n1135 = ~n645 & ((~x4 & x5 & ~x1 & x2) | ((~x2 | ~x5) & (~x1 ^ ~x4)));
  assign n1136 = (x1 | n1137) & (~x1 | ~x4 | x6 | n1139);
  assign n1137 = (x0 | x3 | x4 | ~n1121) & (~x0 | ~x3 | n1138);
  assign n1138 = (~x2 | ~x4 | ~x5 | x6) & (x2 | x4 | x5 | ~x6);
  assign n1139 = (~x0 | x2 | ~x3 | x5) & (x0 | x3 | (~x2 ^ x5));
  assign n1140 = (n645 | n1141) & (x2 | (n1143 & (n645 | n1142)));
  assign n1141 = (~x6 | ((x1 | ~x2 | ~x4 | ~x5) & (~x1 | (x2 ? (x4 | ~x5) : (~x4 | x5))))) & (x1 | x4 | x6 | (~x2 ^ x5));
  assign n1142 = (x1 | x4 | x5 | x6 | ~x7) & (~x1 | ~x4 | ~x5 | ~x6 | x7);
  assign n1143 = ~n1144 & n1146 & (~x0 | ~n620 | ~n1145);
  assign n1144 = ~n565 & ~n1016 & (x0 ? n400 : n314);
  assign n1145 = x7 & ~x6 & ~x4 & x5;
  assign n1146 = (n481 | n1148) & (~n441 | ~n465 | ~n1147);
  assign n1147 = x6 & (~x4 ^ ~x7);
  assign n1148 = (~x0 | x1 | ~x3 | ~x5) & (x0 | ~x1 | x3 | x5);
  assign z041 = ~n1165 | n1159 | n1150 | n1157;
  assign n1150 = ~x0 & (n1152 | n1155 | (n1151 & ~n1156));
  assign n1151 = ~x2 & x7;
  assign n1152 = ~x7 & ((n408 & n1154) | (x2 & ~n1153));
  assign n1153 = (~x4 | ((~x1 | x6 | (~x3 ^ ~x5)) & (~x5 | ~x6 | x1 | ~x3))) & (x1 | x4 | x5 | (~x3 ^ x6));
  assign n1154 = ~x4 & x5 & (~x3 ^ ~x6);
  assign n1155 = ~n1036 & ((~x1 & x2 & x4 & x7) | (x1 & (x2 ? (~x4 & x7) : (x4 & ~x7))));
  assign n1156 = x1 ? ((x5 | x6 | x3 | ~x4) & (~x5 | ~x6 | ~x3 | x4)) : ((x5 | ~x6 | x3 | x4) & (~x3 | (x4 ? (~x5 | ~x6) : (x5 | x6))));
  assign n1157 = x2 & ((n457 & n512) | (~x0 & ~n1158));
  assign n1158 = (~x1 | (x3 ? (x4 ? (x5 | ~x6) : (~x5 | x6)) : (x6 | (x4 ^ x5)))) & (x1 | ~x3 | x4 | ~x5 | ~x6);
  assign n1159 = ~x2 & (n1160 | n1162 | (x0 & ~n1164));
  assign n1160 = n387 & (n1161 | (x3 & x6 & ~n677));
  assign n1161 = ~x6 & x5 & ~x3 & ~x4;
  assign n1162 = ~n1163 & ((~x0 & ~x1 & x4 & ~x5) | (x0 & (x1 ? (x4 & x5) : (~x4 & ~x5))));
  assign n1163 = x3 ^ ~x6;
  assign n1164 = (~x1 | ~x3 | x4 | ~x5 | ~x6) & (x1 | x3 | ~x4 | x5 | x6);
  assign n1165 = n1169 & (~x0 | (n1167 & (n1163 | n1166)));
  assign n1166 = (x2 | (x5 ^ x7) | (x1 ^ ~x4)) & (x1 | ~x2 | (x4 ? (x5 | ~x7) : (~x5 | x7)));
  assign n1167 = (~n269 | ~n270) & (n573 | ~n1168);
  assign n1168 = x1 & x6;
  assign n1169 = x1 ? n1171 : n1170;
  assign n1170 = ((~x0 ^ ~x2) | (x3 ? (x5 | ~x6) : (~x5 | x6))) & (x0 | ~x2 | x3 | x5 | x6) & (~x5 | ((~x0 | x2 | ~x3 | ~x6) & (x0 | ~x2 | (~x3 ^ x6))));
  assign n1171 = (~x0 | x2 | x3 | x5 | x6) & (x0 | ((~x5 | ~x6 | ~x2 | x3) & (x2 | x5 | (~x3 ^ x6))));
  assign z042 = n1189 | ~n1194 | (x2 ? ~n1173 : ~n1180);
  assign n1173 = (x5 & ~n1174 & ~n1175 & ~n1176) | (~x5 & n1178);
  assign n1174 = ~n565 & ((x0 & ~x1 & x3 & ~x4) | (~x0 & (x1 ? (~x3 ^ x4) : (~x3 & x4))));
  assign n1175 = n276 & ((n382 & n601) | (x0 & ~n485));
  assign n1176 = n635 & n1177;
  assign n1177 = x3 & ~x0 & x1;
  assign n1178 = (~x0 | x1 | ~x3 | n481) & (x0 | (x1 ? (x3 | n481) : (~x3 | ~n1179)));
  assign n1179 = ~x4 & (~x6 ^ ~x7);
  assign n1180 = x6 ? (n1186 & (x7 | n1181)) : (n1182 & (~x7 | n1181));
  assign n1181 = x0 ? ((~x1 | ~x3 | x4 | x5) & (x1 | (x3 ? ~x4 : (x4 | x5)))) : ((x1 | ~x3 | x4) & (~x1 | x3 | ~x4 | x5));
  assign n1182 = (~n765 | ~n1183) & (n1184 | n1185);
  assign n1183 = x7 & ~x4 & ~x5;
  assign n1184 = x1 ? (~x5 | ~x7) : (x5 | x7);
  assign n1185 = x0 ? (~x3 | x4) : (x3 | ~x4);
  assign n1186 = (~n1063 | ~n1187) & (x3 | n826 | n1188);
  assign n1187 = x7 & x4 & x5;
  assign n1188 = x1 ? (~x5 | x7) : (x5 | ~x7);
  assign n1189 = ~n542 & (n1190 | n1191 | n1192);
  assign n1190 = x4 & x3 & x2 & ~x0 & ~x1;
  assign n1191 = ~n1091 & ((x3 & ~x4 & ~x0 & x1) | (~x3 & (x0 ? (x1 ^ x4) : (~x1 & ~x4))));
  assign n1192 = n725 & ((n425 & n659) | (x0 & ~n1193));
  assign n1193 = x3 ? (~x4 | ~x5) : (x4 | x5);
  assign n1194 = n1197 & (~x2 | (~n1196 & (x0 | n1195)));
  assign n1195 = (x1 | x3 | ~x4 | x5 | ~x6) & (~x1 | ((~x3 | ~x6 | (x4 ^ ~x5)) & (x3 | ~x4 | ~x5 | x6)));
  assign n1196 = ~x4 & n1064 & (x1 ? (x5 & x6) : ~x6);
  assign n1197 = ~n1198 & (x2 | ((~n301 | ~n1177) & ~n1199));
  assign n1198 = ~n1163 & ((~x0 & n932) | (~n1119 & ~n826));
  assign n1199 = n363 & (x3 ? (~x4 & x6) : (~x6 & (~x4 ^ ~x5)));
  assign z043 = ~n1212 | ~n1210 | n1206 | n1201 | n1204;
  assign n1201 = ~x3 & (x5 ? ~n1202 : ~n1203);
  assign n1202 = ((x1 ^ x2) | (x0 ? (x4 | x7) : (~x4 ^ x7))) & (~x1 | x2 | x4 | (~x0 ^ ~x7));
  assign n1203 = (x0 | ~x1 | x2 | x4 | x7) & (~x0 | ((x4 | x7 | x1 | ~x2) & (~x1 | x2 | (~x4 ^ x7))));
  assign n1204 = x3 & ((~x5 & ~n1205) | (n300 & n1187));
  assign n1205 = (x0 | x1 | x2 | ~x4 | x7) & (~x7 | (((~x1 ^ x4) | (x0 ^ ~x2)) & (x0 | x1 | x2 | x4)));
  assign n1206 = x1 & (x7 ? (n1207 & ~n1209) : ~n1208);
  assign n1207 = ~x2 & x4;
  assign n1208 = (~n320 | ~n661) & (x4 | n315 | n966);
  assign n1209 = (~x0 | x3 | ~x5 | ~x6) & (x0 | x6 | (x3 ^ ~x5));
  assign n1210 = x5 ? ((~x7 | n1211) & (~x3 | x7 | n418)) : ((x7 | n1211) & (x3 | ~x7 | n418));
  assign n1211 = (~x4 | (x0 ^ ~x2) | (~x1 ^ ~x3)) & (~x3 | x4 | (x0 ? (x1 | ~x2) : (~x1 | x2)));
  assign n1212 = ~n1213 & (x1 | (~n1216 & ~n1218));
  assign n1213 = ~n688 & ((n579 & ~n1215) | (x2 & ~n1214));
  assign n1214 = x5 ? ((~x0 | x1 | x3 | ~x6) & (x0 | ~x1 | ~x3 | x6)) : (x0 ? (x1 ? (x3 | x6) : (~x3 | ~x6)) : (x1 ? (x3 | ~x6) : (~x3 | x6)));
  assign n1215 = (~x1 | x3 | ~x5 | ~x6) & (x1 | (x3 ? (~x5 | x6) : (x5 | ~x6)));
  assign n1216 = x0 & (x6 ? (n484 & ~n1024) : ~n1217);
  assign n1217 = (x2 | ~x3 | ~x4 | ~x5 | ~x7) & (~x2 | ((~x3 | ~x4 | x5 | ~x7) & (~x5 | x7 | x3 | x4)));
  assign n1218 = ~x0 & (x2 ? (n606 & n556) : ~n1219);
  assign n1219 = x3 ? ((~x4 | ~x5 | ~x6 | ~x7) & (x6 | x7 | x4 | x5)) : (x5 | (x4 ? (x6 | ~x7) : (~x6 | x7)));
  assign z044 = n1227 | n1232 | (x3 ? ~n1221 : ~n1238);
  assign n1221 = x0 ? n1224 : (x4 ? n1222 : n1223);
  assign n1222 = (~x1 | ~x2 | ~x5 | x6 | ~x7) & (x1 | x2 | x5 | ~x6 | x7) & ((~x5 ^ x7) | (x1 ? (x2 | ~x6) : (~x2 | x6)));
  assign n1223 = (x1 | x2 | ~x5 | ~x6 | ~x7) & (x5 | (~x2 ^ ~x6) | (x1 ^ ~x7));
  assign n1224 = x2 ? (x1 | (~n296 & ~n1226)) : n1225;
  assign n1225 = (x6 | (x1 ? (x4 ? (x5 | x7) : (~x5 | ~x7)) : (x4 | (~x5 ^ x7)))) & (~x4 | ~x5 | ~x6 | (x1 ^ ~x7));
  assign n1226 = ~x4 & x6 & (x5 ^ x7);
  assign n1227 = x1 & (n1229 | n1231 | (~x2 & ~n1228));
  assign n1228 = (~x3 | ~x4 | ~x5 | x6) & (x4 | ((~x0 | x3 | x5 | ~x6) & (x0 | (x3 ? ~x5 : (x5 | x6)))));
  assign n1229 = ~n379 & (n413 | (~x2 & ~n1230));
  assign n1230 = (~x0 | ~x3 | x4) & (x3 | ~x4);
  assign n1231 = n426 & ((n1039 & n330) | (~x0 & n587));
  assign n1232 = ~x1 & (n1234 | ~n1236 | (x0 & ~n1233));
  assign n1233 = (~x2 | x3 | ~x4 | ~x5 | ~x6) & (x2 | (x3 ? (x5 | (~x4 & ~x6)) : (~x5 | x6)));
  assign n1234 = ~n379 & ((n324 & n606) | (~x0 & ~n1235));
  assign n1235 = x2 ? (x3 | x4) : (~x3 | ~x4);
  assign n1236 = (~n340 | n534) & (x0 | (n1237 & (~n339 | n534)));
  assign n1237 = (~x2 | x3 | ~x4 | ~x5 | x6) & (x2 | ~x3 | x4 | x5 | ~x6);
  assign n1238 = n1240 & (~n430 | ~n742) & (n868 | n1239);
  assign n1239 = (x2 | x4 | ~x6 | x7) & (~x2 | ~x4 | x6 | ~x7);
  assign n1240 = ~n1242 & (n854 | n978) & (n585 | ~n1241);
  assign n1241 = ~x2 & ~x0 & ~x1;
  assign n1242 = ~n1243 & ((n425 & n363) | (n424 & n387));
  assign n1243 = x2 ? (x6 | x7) : (~x6 | ~x7);
  assign z045 = n1269 | n1264 | ~n1253 | n1245 | n1251;
  assign n1245 = ~x0 & (n1248 | (~x1 & (n1246 | n1247)));
  assign n1246 = x2 & ((n656 & n588) | (n280 & n606));
  assign n1247 = n366 & ((~x3 & x5 & ~x6 & ~x7) | (x7 & (x3 ? (~x5 ^ x6) : (~x5 & x6))));
  assign n1248 = x1 & (x7 ? (n465 & ~n1249) : ~n1250);
  assign n1249 = x2 ? (~x4 | x6) : (x4 | ~x6);
  assign n1250 = x2 ? (~x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))) : (x3 | ~x4 | (x5 ^ x6));
  assign n1251 = x6 & ((n364 & n609) | (~x0 & ~n1252));
  assign n1252 = (~x2 | ~x3 | x4 | ~x5) & (x3 | ((~x1 | ~x2 | x4 | x5) & (x1 | x2 | (~x4 ^ x5))));
  assign n1253 = n1258 & (n1255 | n1257) & (n1254 | n1256);
  assign n1254 = ~x4 ^ ~x6;
  assign n1255 = ~x1 ^ ~x5;
  assign n1256 = (x0 | ~x1 | x2 | x3 | x5) & (x1 | ((~x0 | (x2 ? (~x3 | x5) : (x3 | ~x5))) & (~x3 | ~x5 | x0 | x2)));
  assign n1257 = (~x0 | x2 | ~x3 | ~x4 | x6) & (x3 | ((x0 | ~x2 | ~x4 | x6) & (~x0 | x4 | (~x2 ^ ~x6))));
  assign n1258 = x0 ? (~n1260 & n1261) : (~n725 | ~n1259);
  assign n1259 = ~x6 & x5 & x3 & ~x4;
  assign n1260 = ~n1163 & n424 & x7 & n408;
  assign n1261 = (n481 | n503) & (n1262 | n1263);
  assign n1262 = x3 ? (~x6 | ~x7) : (x6 | x7);
  assign n1263 = (~x1 | x2 | ~x4 | ~x5) & (x1 | ~x2 | x4 | x5);
  assign n1264 = ~n542 & ((n428 & n1265) | n1266 | n1267);
  assign n1265 = ~x5 & ~x3 & x4;
  assign n1266 = n730 & (x1 ? (~x2 & ~n436) : (x2 & n356));
  assign n1267 = ~n736 & (n1268 | (~x0 & n400));
  assign n1268 = x0 & (x1 ? (~x3 & ~x5) : (x3 & x5));
  assign n1269 = ~n565 & ((n428 & n1270) | n1271 | n1272);
  assign n1270 = ~x5 & x3 & ~x4;
  assign n1271 = n730 & ((~x1 & ~x2 & ~x3 & x4) | (x2 & ((~x3 & ~x4) | (x1 & x3 & x4))));
  assign n1272 = ~n468 & (x0 ? (~x3 ^ x5) : (x3 & ~x5));
  assign z046 = n1277 | ~n1281 | ~n1288 | (~n1274 & ~n1275);
  assign n1274 = ~x0 ^ ~x3;
  assign n1275 = (x7 | n1276) & (x1 | ~n624 | ~n313);
  assign n1276 = (x1 | ~x2 | x4 | x5 | x6) & (x2 | ((~x5 | ~x6 | x1 | x4) & (~x1 | ~x4 | (~x5 ^ x6))));
  assign n1277 = ~n444 & ((~n1278 & ~n1279) | (~x2 & ~n1280));
  assign n1278 = x1 ? (x3 | x5) : (~x3 | ~x5);
  assign n1279 = x2 ? (~x4 | x7) : (x4 | ~x7);
  assign n1280 = (~x1 | x3 | ~x4 | ~x5 | ~x7) & (x1 | ~x3 | x4 | x5 | x7);
  assign n1281 = ~n1283 & ~n1285 & n1287 & (n570 | n1282);
  assign n1282 = (~x3 | ((~x2 | ~x4 | x0 | ~x1) & (~x0 | (x1 ? (x2 | x4) : ~x4)))) & (x0 | x3 | (~x1 ^ x4));
  assign n1283 = ~n574 & (n1284 | (~n271 & n1064));
  assign n1284 = x3 & x2 & ~x0 & ~x1;
  assign n1285 = ~n1286 & ((n725 & n1074) | (n438 & n760));
  assign n1286 = (~x0 | x3 | ~x5 | ~x6) & (x0 | ~x3 | x5 | x6);
  assign n1287 = (n675 | n1111) & (~n789 | ~n295 | ~n588);
  assign n1288 = n1290 & n1294 & (~n473 | n1289);
  assign n1289 = x0 ? ((~x2 | ~x3 | ~x5 | ~x7) & (x5 | x7 | x2 | x3)) : ((x2 | (x3 ? (~x5 | x7) : (x5 | ~x7))) & (~x5 | ~x7 | ~x2 | x3));
  assign n1290 = (n574 | n1293) & (n1291 | n1292);
  assign n1291 = x5 ^ ~x7;
  assign n1292 = (~x0 | ~x1 | ~x2 | x3 | x4) & (x0 | x2 | ~x3 | (~x1 ^ x4));
  assign n1293 = (~x0 | x1 | x2 | x3 | x6) & (x0 | ~x1 | ~x2 | (x3 ^ x6));
  assign n1294 = (n1296 | n1297) & (~x7 | ~n1295 | n1298);
  assign n1295 = ~x1 & x5;
  assign n1296 = (~x1 | x2 | ~x3 | ~x7) & (x1 | ~x2 | x3 | x7);
  assign n1297 = (~x5 | x6 | x0 | ~x4) & (~x0 | ~x6 | (x4 ^ x5));
  assign n1298 = (~x0 | x2 | x3 | x4 | ~x6) & (x0 | x6 | (x2 ? (~x3 | ~x4) : (x3 | x4)));
  assign z047 = ~n1311 | ~n1317 | (x2 ? ~n1305 : ~n1300);
  assign n1300 = x0 ? n1301 : (~n1304 & (x3 | n1303));
  assign n1301 = (x7 | n1302) & (~x1 | ~n526);
  assign n1302 = (x3 | x4 | (x1 ? (~x5 | x6) : (x5 | ~x6))) & (x1 | ~x4 | ((x5 | x6) & (~x3 | ~x5 | ~x6)));
  assign n1303 = (x1 | ~x4 | ~x5 | ~x6 | x7) & (x5 | ((x6 | x7 | x1 | ~x4) & (~x7 | (x1 ? (~x4 ^ x6) : (x4 | x6)))));
  assign n1304 = n588 & ((x6 & ~x7 & ~x1 & x5) | (x1 & x7 & (~x5 ^ x6)));
  assign n1305 = ~n1309 & (x0 | (~n1307 & (x4 | n1306)));
  assign n1306 = (x1 | ~x3 | x5 | ~x6 | ~x7) & (~x5 | (x1 ? ((x6 | ~x7) & (x3 | ~x6 | x7)) : (x6 | x7)));
  assign n1307 = n588 & ((n521 & n346) | (x1 & ~n1308));
  assign n1308 = x5 ? (x6 | x7) : (~x6 | ~x7);
  assign n1309 = ~n1310 & x5 & n363;
  assign n1310 = (~x3 | x4 | x6 | x7) & (~x4 | ((x6 | ~x7) & (x3 | ~x6 | x7)));
  assign n1311 = ~n1313 & (n379 | n1312) & (~n1207 | n1316);
  assign n1312 = (~x0 | x2 | x3 | (~x1 ^ ~x4)) & (~x2 | ((x1 | ~x3 | ~x4) & (x0 | (x1 ? (~x3 | x4) : ~x4))));
  assign n1313 = ~x4 & ((n359 & n1314) | (~n1029 & ~n1315));
  assign n1314 = x6 & ~x3 & ~x5;
  assign n1315 = (~x0 | ~x2 | x3) & (x2 | ~x3);
  assign n1316 = x1 ? (~x6 | (x0 ? ~x3 : x5)) : (x6 | ((~x3 | ~x5) & (x0 | (~x3 & ~x5))));
  assign n1317 = (n1091 | n1319) & (n1318 | (~n1320 & ~n1321));
  assign n1318 = x1 ^ ~x7;
  assign n1319 = (x1 | ((x0 | x3 | x4 | ~x6) & (~x0 | (x3 ? (x4 | ~x6) : (~x4 | x6))))) & (x0 | ~x1 | x3 | (x4 ^ x6));
  assign n1320 = ~x3 & (x4 ? ~n311 : (n324 & ~n379));
  assign n1321 = ~x4 & n423 & ((~x5 & ~x6) | (~x0 & x5 & x6));
  assign z048 = ~n1332 | (~n565 & ~n1329) | (~x0 & ~n1323);
  assign n1323 = x1 ? n1324 : (n1328 & (x6 | n1327));
  assign n1324 = x3 ? n1325 : n1326;
  assign n1325 = (x2 | ~x4 | ~x5 | x6 | ~x7) & (~x2 | x4 | x5 | ~x6 | x7);
  assign n1326 = x5 ? (x2 ? (~x7 | (x4 & x6)) : (x7 | (x4 & ~x6))) : (x2 ? (x7 | (~x4 & ~x6)) : (x6 | ~x7));
  assign n1327 = (x2 | ~x7 | (x3 ? (x4 | ~x5) : (~x4 | x5))) & (~x2 | x3 | x4 | x5 | x7);
  assign n1328 = x2 ? (x3 ? (~x4 | n563) : n555) : (x3 ? (~x4 | n555) : (x4 | n563));
  assign n1329 = (x4 | n1330) & (~x3 | ~x4 | n605 | n1331);
  assign n1330 = x0 ? (x3 | ((~x2 | x5) & (~x1 | x2 | ~x5))) : (~x3 | (x2 ^ x5));
  assign n1331 = x0 ^ ~x1;
  assign n1332 = ~n1337 & (n542 | (n1334 & (x2 | n1333)));
  assign n1333 = x0 ? ((x1 | ~x3 | x4 | ~x5) & (~x1 | x3 | ~x4 | x5)) : (x3 | x4 | (~x1 ^ x5));
  assign n1334 = ~n1335 & ~n1336 & (~n438 | ~n425 | n1274);
  assign n1335 = ~x2 & ((~x4 & ~x5 & x0 & ~x3) | (x5 & ((x3 & x4) | (~x0 & (x3 | x4)))));
  assign n1336 = x2 & ((~x4 & x5 & x0 & ~x3) | (~x0 & x3 & ~x5));
  assign n1337 = x0 & ((~x2 & ~n1338) | (n438 & ~n1339));
  assign n1338 = (x1 & (x4 ? n563 : ~x3)) | (n563 & n1308) | (~x1 & (x4 ? x3 : n563));
  assign n1339 = x4 ? ((x5 | ~x6 | x7) & (x3 | ~x5 | ~x7)) : ((~x5 | x6 | ~x7) & (~x3 | x5 | x7));
  assign z049 = ~n1355 | (x3 ? ~n1341 : (n1346 | n1351));
  assign n1341 = ~n1344 & (n565 | n1343) & (n605 | n1342);
  assign n1342 = (x0 | ~x1 | x4 | x6 | ~x7) & (~x4 | ((~x0 | x1 | x6 | ~x7) & (x0 | ((~x6 | ~x7) & (x1 | x6 | x7)))));
  assign n1343 = (~x1 | ((~x0 | x2 | ~x4) & (x4 | x5 | x0 | ~x2))) & (~x0 | x1 | ((~x2 | ~x4 | x5) & (x4 | (x2 & ~x5))));
  assign n1344 = ~x0 & ((n932 & n921) | (~n542 & ~n1345));
  assign n1345 = (~x1 | x2 | ~x4 | ~x5) & (x1 | (x2 ? (~x4 | x5) : (x4 | ~x5)));
  assign n1346 = ~x5 & (n1348 | n1350 | (x4 & ~n1347));
  assign n1347 = (x6 | x7 | ~x0 | ~x2) & (x0 | ((x1 | ((x6 | ~x7) & (~x2 | ~x6 | x7))) & (x2 | ((x6 | ~x7) & (~x1 | ~x6 | x7)))));
  assign n1348 = ~n1349 & (x1 ? (~x4 & ~x6) : x6);
  assign n1349 = x0 ? (~x2 | ~x7) : (x2 | x7);
  assign n1350 = ~n542 & ((x2 & ~x4 & ~x0 & x1) | (x0 & ~x2 & (x1 ^ ~x4)));
  assign n1351 = x5 & (~n1353 | (x7 & ~n1352));
  assign n1352 = (~x1 | ((x0 | ~x4 | x6) & (x4 | ~x6 | ~x0 | x2))) & (x0 | x6 | ((~x2 | ~x4) & (x1 | x2 | x4)));
  assign n1353 = (n389 | n1354) & (~n782 | ~n622);
  assign n1354 = x1 ? (x2 | ~x4) : x4;
  assign n1355 = n1356 & (x1 ? n1360 : n1359);
  assign n1356 = x1 ? n1358 : n1357;
  assign n1357 = (x0 | ~x2 | ~x3 | x4 | x6) & (~x0 | x2 | x3 | ~x4 | ~x6);
  assign n1358 = (x0 | ~x2 | ~x3 | ~x4 | x6) & (x2 | x4 | (x0 ? (x3 ^ x6) : (x3 | ~x6)));
  assign n1359 = x0 ? ((~x3 | n936) & (~x2 | x3 | n602)) : ((x2 | ~x3 | n602) & (x3 | n936));
  assign n1360 = (~n312 | ~n512) & (x0 | n614 | n761);
  assign z050 = n1362 | n1365 | ~n1373 | (~x3 & ~n1368);
  assign n1362 = ~x4 & (x2 ? ~n1364 : ~n1363);
  assign n1363 = (~x7 | ((~x0 | ~x1 | x3 | x5) & (x0 | ~x3 | (~x1 ^ ~x5)))) & (x1 | ~x5 | x7 | (x0 & ~x3));
  assign n1364 = (x1 | ((x0 | x3 | x5 | ~x7) & (~x0 | ((~x3 | x5 | ~x7) & (~x5 | x7))))) & (x0 | ~x1 | ((x5 | x7) & (x3 | ~x5 | ~x7)));
  assign n1365 = x3 & ((~n836 & ~n1366) | (n382 & ~n1367));
  assign n1366 = (~x0 | x1 | x2 | x5 | x7) & (x0 | ~x1 | ~x7 | (x2 ^ x5));
  assign n1367 = (~x0 | x1 | ~x2 | ~x4 | ~x5) & (x0 | ((~x4 | ~x5 | x1 | x2) & (~x1 | x4 | (x2 ^ x5))));
  assign n1368 = (~n1369 | n1372) & (n1371 | (~n1370 & ~n1179));
  assign n1369 = x1 & ~x7;
  assign n1370 = x7 & x4 & x6;
  assign n1371 = x0 ? (x1 ? (x2 | ~x5) : (~x2 | x5)) : (x1 | (x2 ^ x5));
  assign n1372 = (~x2 | ((x5 | x6 | ~x0 | x4) & (~x5 | ~x6 | x0 | ~x4))) & (x0 | x2 | x5 | (x4 ^ x6));
  assign n1373 = n1376 & (x3 | n1374) & (~x4 | n1375);
  assign n1374 = (~x0 | x1 | x2 | ~x4 | ~x7) & (x4 | ((~x0 | (x1 ? (~x2 | ~x7) : (x2 | x7))) & (x0 | ~x1 | x2 | ~x7)));
  assign n1375 = (x0 | ~x1 | (x2 ? (x5 | ~x7) : (~x5 | x7))) & (x1 | (x5 ^ x7) | (~x0 ^ ~x2));
  assign n1376 = (~x4 | x7 | n420) & (~x3 | ~x7 | (x4 ? ~n428 : n420));
  assign z051 = n1378 | ~n1384 | n1388 | (~x5 & ~n1387);
  assign n1378 = x1 & (n1380 | n1382 | (~n506 & ~n1379));
  assign n1379 = (~x0 | x2 | x4 | x5 | ~x7) & (x0 | ~x5 | (x2 ? (~x4 | x7) : (x4 | ~x7)));
  assign n1380 = ~n1381 & (x0 ? n314 : n400);
  assign n1381 = (~x6 | x7 | x2 | ~x4) & (~x2 | x4 | x6 | ~x7);
  assign n1382 = n1383 & ((n382 & n924) | (x0 & n327));
  assign n1383 = ~x4 & x2 & ~x3;
  assign n1384 = x5 ? n1385 : (x6 | n1386);
  assign n1385 = (x0 & (x2 | (x1 & ~x3 & x6))) | (x1 & x2 & (~x3 | x6)) | (~x1 & ((~x2 & x3 & ~x6) | (~x0 & ~x3 & x6))) | (~x0 & ~x2 & (x3 | ~x6));
  assign n1386 = ((x2 ^ x7) | (x0 ? (x1 | ~x3) : (~x1 | x3))) & (x0 | x1 | x2 | ~x7) & (~x0 | ~x1 | ~x2 | x3 | x7);
  assign n1387 = x6 ? (x0 ? (x1 ? (x2 | x3) : (~x2 | ~x3)) : ((x1 | x2 | ~x3) & (~x2 | (~x1 & x3)))) : ((x2 | ~x3 | x0 | ~x1) & (~x0 | x1 | ~x2 | x3));
  assign n1388 = ~x1 & (n1391 | n1392 | (~x4 & ~n1389));
  assign n1389 = x0 ? (~x2 | n583) : (x2 ? (x5 | ~n1390) : n583);
  assign n1390 = x7 & (x3 ^ ~x6);
  assign n1391 = ~n753 & ((n579 & n1074) | (x0 & ~n1279));
  assign n1392 = n285 & n1074 & (x2 ? n327 : n328);
  assign z052 = n1394 | ~n1400 | ~n1404 | (n327 & ~n1399);
  assign n1394 = ~x6 & ((n300 & n1043) | n1395 | n1397);
  assign n1395 = ~x2 & ((n765 & n1183) | (x3 & ~n1396));
  assign n1396 = (x0 | ~x1 | ~x4 | ~x5 | ~x7) & (~x0 | ((x5 | x7 | x1 | ~x4) & (~x5 | ~x7 | ~x1 | x4)));
  assign n1397 = ~n1398 & (x1 ? n450 : n786);
  assign n1398 = (~x3 | x4 | x0 | ~x2) & (x3 | (x0 ? (~x2 ^ ~x4) : (x2 | ~x4)));
  assign n1399 = x1 ? ((~x3 | ~x4 | ~x0 | x2) & (x3 | x4 | x0 | ~x2)) : (x0 ? (x2 ? (~x3 | x4) : (x3 | ~x4)) : (~x3 | (x2 ^ x4)));
  assign n1400 = n1401 & (n565 | (n611 & (n420 | n766)));
  assign n1401 = (n766 | n1403) & (n987 | n1402);
  assign n1402 = x0 ? (x1 | x6) : (~x1 | ~x6);
  assign n1403 = (~x0 | x1 | ~x2 | ~x6) & (x0 | x2 | (~x1 ^ x6));
  assign n1404 = n1406 & (n565 | n614 | n1405);
  assign n1405 = (~x0 | x1 | ~x2 | x3) & (x0 | x2 | (~x1 ^ ~x3));
  assign n1406 = (n614 | n1408) & (n542 | n1407);
  assign n1407 = ((x2 ^ x4) | (x0 ? (x1 | ~x3) : (~x1 | x3))) & (~x0 | ~x1 | ~x2 | x3 | x4) & (x0 | x1 | x2 | ~x3 | ~x4);
  assign n1408 = (~x0 | x1 | x2 | x3 | ~x6) & (x0 | ~x1 | ~x2 | ~x3 | x6) & ((x0 ? (~x1 | x2) : (x1 | ~x2)) | (x3 ^ x6));
  assign z053 = n1410 | n1413 | ~n1419 | (x0 & ~n1418);
  assign n1410 = ~x2 & (x0 ? ~n1411 : ~n1412);
  assign n1411 = x1 ? ((x3 | (x4 ? (~x5 ^ x7) : (~x5 | ~x7))) & (x5 | x7 | ~x3 | x4)) : ((~x3 | ~x4 | ~x5 | ~x7) & (x5 | x7 | x3 | x4));
  assign n1412 = (~x1 | x3 | ~x4 | ~x5 | ~x7) & ((~x1 ^ ~x3) | (x4 ? (x5 | x7) : (~x5 ^ x7)));
  assign n1413 = ~n542 & (n724 | n1415 | (x0 & ~n1414));
  assign n1414 = (~x1 | x2 | ~x3 | x4 | ~x5) & (x1 | ~x4 | (x2 ? (x3 | ~x5) : (~x3 | x5)));
  assign n1415 = ~n1417 & (n1416 | (~x0 & ~n986));
  assign n1416 = ~x4 & ~x3 & x0 & ~x2;
  assign n1417 = x1 ^ ~x5;
  assign n1418 = x1 ? ((~x4 | ~x7 | x2 | ~x3) & (x4 | x7 | ~x2 | x3)) : ((~x4 | ~x7 | x2 | x3) & (~x3 | (x2 ? (~x4 ^ x7) : (x4 | x7))));
  assign n1419 = ~n1420 & (x0 | n1426) & (~x2 | n1421);
  assign n1420 = n410 & n411;
  assign n1421 = ~n1423 & ~n1425 & (~x0 | ~n276 | ~n1422);
  assign n1422 = ~x7 & x4 & ~x5;
  assign n1423 = n601 & ((n620 & n786) | (~x1 & ~n1424));
  assign n1424 = x3 ? (x5 | x7) : (~x5 | ~x7);
  assign n1425 = ~n1291 & ((n363 & n606) | (n329 & ~n954));
  assign n1426 = (x1 | ~x2 | ~x3 | ~x4 | ~x7) & (~x1 | x2 | x3 | x4 | x7) & ((x1 ? (~x2 | x3) : (x2 | ~x3)) | (~x4 ^ x7));
  assign z054 = ~n1438 | ~n1441 | (x6 ? ~n1428 : ~n1429);
  assign n1428 = ~n724 & ~n1415 & (~x0 | n1414);
  assign n1429 = n1432 & (x3 | (x2 & n1431) | (~x2 & n1430));
  assign n1430 = (~x0 | ~x1 | x4 | ~x5 | ~x7) & (x0 | x1 | ~x4 | x5 | x7);
  assign n1431 = (x7 | ((x0 | ~x1 | ~x4 | ~x5) & (~x0 | (x1 ? (x4 | ~x5) : (~x4 | x5))))) & (x0 | x4 | ~x7 | (~x1 ^ x5));
  assign n1432 = (n350 | n1433) & (~x3 | (~n1434 & ~n1437));
  assign n1433 = x0 ? (x2 | (x1 ? (~x3 | x5) : (x3 ^ x5))) : ((~x1 | x2 | x3 | ~x5) & (x1 | ~x2 | ~x3 | x5));
  assign n1434 = ~n1436 & ~x1 & ~n1435;
  assign n1435 = x4 ? (~x5 | x7) : (x5 | ~x7);
  assign n1436 = ~x0 ^ ~x2;
  assign n1437 = n387 & ((n624 & n786) | (n1207 & n450));
  assign n1438 = ~n1439 & ~n1440 & (~n387 | n1011 | n498);
  assign n1439 = ~n1012 & ((x1 & ~x3 & ~x7) | (x0 & (x1 ? ~x3 : (x3 & ~x7))));
  assign n1440 = ~x1 & ((n647 & n1270) | (n782 & n609));
  assign n1441 = ~n1442 & (x7 | ((~n428 | ~n1265) & ~n1443));
  assign n1442 = ~n989 & ((x0 & (x1 ? (~x2 & ~x7) : x2)) | (~x1 & (x2 ? ~x7 : ~x0)));
  assign n1443 = ~x4 & n659 & (x1 ? n483 : n484);
  assign z055 = n1445 | ~n1448 | ~n1455 | (~n1308 & ~n1399);
  assign n1445 = x0 & (n1446 | (~x1 & ~n1447));
  assign n1446 = ~n998 & ((n335 & n625) | (~x1 & ~n989));
  assign n1447 = (~x2 | x3 | ~x4 | ~x5 | ~x6) & (x2 | ~x3 | x4 | x5 | x6);
  assign n1448 = ~n1449 & ~n1450 & ~n1454 & (~n363 | n1452);
  assign n1449 = ~n822 & ((~x0 & x2 & (x1 ^ x5)) | (x0 & x1 & ~x2 & x5));
  assign n1450 = ~n1451 & ((n339 & n480) | (n782 & ~n954));
  assign n1451 = (x4 | ~x5 | ~x6 | ~x7) & (~x4 | x5 | x6 | x7);
  assign n1452 = (~n892 | ~n876) & (~n1453 | ~n875);
  assign n1453 = x4 & ~x2 & x3;
  assign n1454 = n575 & ((n356 & n875) | (n443 & n876));
  assign n1455 = ~n1460 & (n565 | (~n1456 & n1457));
  assign n1456 = n438 & ((~x0 & x3 & ~x4 & ~x5) | (x0 & x4 & (x3 ^ ~x5)));
  assign n1457 = x0 ? (x4 | n1459) : ((~n725 | ~n1458) & (~x4 | n1459));
  assign n1458 = x5 & ~x3 & ~x4;
  assign n1459 = x1 ? (x2 ? (x3 | ~x5) : (~x3 | x5)) : (x2 | (x3 ^ x5));
  assign n1460 = ~x0 & (x2 ? ~n1461 : ~n1462);
  assign n1461 = (x1 | x3 | x4 | x5 | ~x6) & (~x1 | ~x3 | ~x4 | ~x5 | x6);
  assign n1462 = (x1 | ~x3 | ~x4 | x5 | x6) & ((x4 ^ x6) | (x1 ? (~x3 ^ ~x5) : (x3 | ~x5)));
  assign z056 = ~n1467 | (~n542 & ~n1464);
  assign n1464 = n1466 & (n421 | n498) & (x0 | ~n1465);
  assign n1465 = ~x2 & ((x4 & x5 & x1 & ~x3) | (~x4 & ~x5 & ~x1 & x3));
  assign n1466 = (n420 | n989) & (~n394 | ~n1270);
  assign n1467 = n1470 & n1474 & n1475 & (n1468 | n1469);
  assign n1468 = x0 ? (x1 | ~x3) : (~x1 | x3);
  assign n1469 = (x2 | ~x4 | x5 | ~x6 | x7) & (~x2 | x4 | ~x5 | x6 | ~x7);
  assign n1470 = n1472 & (n420 | n1111) & (~n1145 | ~n1471);
  assign n1471 = x3 & ~x2 & ~x0 & ~x1;
  assign n1472 = (~n428 | ~n1473) & (~n790 | ~n588 | ~n514);
  assign n1473 = x7 & ~x5 & ~x3 & ~x4;
  assign n1474 = (n570 | n1407) & (n574 | n1405);
  assign n1475 = (n481 | n1477) & (n1405 | (~n270 & ~n1476));
  assign n1476 = ~x7 & x6 & x4 & x5;
  assign n1477 = (~x0 | x1 | x2 | x3 | ~x5) & (x0 | ~x1 | ~x2 | ~x3 | x5) & ((x0 ? (~x1 | x2) : (x1 | ~x2)) | (x3 ^ x5));
  assign z057 = ~n1496 | (x3 ? (n1479 | n1482) : ~n1487);
  assign n1479 = ~x2 & (x0 ? ~n1480 : ~n1481);
  assign n1480 = x1 ? ((~x6 | ~x7 | x4 | x5) & (x7 | (x4 ? (x5 ^ x6) : (~x5 | x6)))) : ((~x4 | ~x5 | x6 | ~x7) & (~x6 | x7 | x4 | x5));
  assign n1481 = (~x1 | ~x4 | ~x5 | x6 | x7) & ((~x1 ^ ~x7) | (x4 ? (x5 | ~x6) : (x5 ^ x6)));
  assign n1482 = x2 & ((n280 & n1483) | n1484 | n1485);
  assign n1483 = x4 & x0 & ~x1;
  assign n1484 = n601 & (x1 ? (x5 & n308) : ~n1308);
  assign n1485 = ~n379 & ((n363 & n342) | (n329 & ~n1486));
  assign n1486 = ~x1 ^ ~x7;
  assign n1487 = ~n1488 & ~n1492 & (n1254 | n1491);
  assign n1488 = ~x0 & (x2 ? ~n1489 : ~n1490);
  assign n1489 = (~x1 | x4 | ~x5 | ~x6 | x7) & (x1 | ~x4 | x5 | x6 | ~x7);
  assign n1490 = x1 ? ((~x4 | ~x5 | x6 | ~x7) & (~x6 | x7 | x4 | x5)) : (~x5 | (x4 ? (x6 | x7) : (~x6 | ~x7)));
  assign n1491 = x1 ? ((~x5 | ~x7 | ~x0 | x2) & (x5 | x7 | x0 | ~x2)) : (x0 ? (x2 ? (x5 | ~x7) : (~x5 | x7)) : (~x7 | (x2 ^ x5)));
  assign n1492 = x0 & ((~n485 & n1493) | (n1494 & ~n1495));
  assign n1493 = ~x1 & (~x2 ^ x5);
  assign n1494 = x1 & ~x5;
  assign n1495 = (x6 | ~x7 | x2 | ~x4) & (~x2 | x7 | (x4 ^ ~x6));
  assign n1496 = ~n1497 & n1501 & (~n782 | n1500);
  assign n1497 = ~x2 & ((n1498 & n1177) | (x7 & ~n1499));
  assign n1498 = ~x7 & ~x4 & x6;
  assign n1499 = (x0 | ~x1 | x3 | x4 | ~x6) & (x1 | ((~x0 | (x3 ? (x4 | ~x6) : (~x4 | x6))) & (~x4 | ~x6 | x0 | ~x3)));
  assign n1500 = (x1 | x3 | x4 | x6 | x7) & (~x1 | ((~x3 | x7 | (x4 ^ x6)) & (x6 | ~x7 | x3 | x4)));
  assign n1501 = (n952 | n1502) & (n1503 | n1504);
  assign n1502 = x3 ? (x6 | ~x7) : (~x6 | x7);
  assign n1503 = x2 ? (~x6 | ~x7) : (x6 | x7);
  assign n1504 = (x3 | ~x4 | x0 | ~x1) & (~x0 | (x1 ? (x3 | x4) : (~x3 | ~x4)));
  assign z058 = ~n1518 | ~n1512 | n1509 | n1413 | n1506;
  assign n1506 = ~n1291 & (x0 ? ~n1507 : ~n1508);
  assign n1507 = x1 ? ((~x2 | x3 | x4 | ~x6) & (x2 | ~x3 | ~x4 | x6)) : ((~x4 | x6 | x2 | x3) & (~x3 | (x2 ? (x4 ^ x6) : (x4 | ~x6))));
  assign n1508 = (~x1 | x2 | x3 | x4 | ~x6) & (x1 | ~x2 | ~x3 | ~x4 | x6) & ((x1 ? (~x2 | x3) : (x2 | ~x3)) | (x4 ^ x6));
  assign n1509 = ~n677 & ((~x0 & ~n1510) | (n647 & ~n1511));
  assign n1510 = (~x1 | x2 | x3 | x6 | ~x7) & (x1 | ~x2 | ~x3 | ~x6 | x7);
  assign n1511 = (~x1 | ~x3 | ~x6 | x7) & (x1 | (x3 ? (x6 | ~x7) : (~x6 | x7)));
  assign n1512 = ~n1513 & ~n1515 & (~n606 | ~n359 | ~n786);
  assign n1513 = ~x0 & ((n269 & n1514) | (~n954 & ~n1469));
  assign n1514 = ~x7 & x6 & ~x4 & ~x5;
  assign n1515 = ~n1517 & (n990 | (~x0 & ~n1516));
  assign n1516 = x1 ? (~x2 | x3) : (x2 | ~x3);
  assign n1517 = (~x6 | x7 | x4 | ~x5) & (~x4 | x5 | x6 | ~x7);
  assign n1518 = (n570 | n1520) & (~n1064 | (~n1519 & ~n1521));
  assign n1519 = n656 & x1 & n366;
  assign n1520 = (x3 | ((x0 | x1 | ~x2 | ~x4) & (~x0 | (x1 ? (x2 | ~x4) : (~x2 | x4))))) & (x0 | ~x1 | ~x3 | (x2 ^ x4));
  assign n1521 = n501 & ((x6 & ~x7 & ~x1 & x4) | (x1 & ~x6 & (x4 ^ x7)));
  assign z059 = n1530 | ~n1533 | (x1 ? ~n1526 : ~n1523);
  assign n1523 = x0 ? n1452 : (x2 ? n1525 : n1524);
  assign n1524 = (~x7 | ((x3 | x4 | x5 | x6) & (~x6 | (x3 ? (x4 ^ x5) : (~x4 | x5))))) & (x6 | x7 | (x3 ? x5 : (x4 | ~x5)));
  assign n1525 = x3 ? (x5 | ((~x6 | ~x7) & (~x4 | x6 | x7))) : (~x5 | ((x6 | x7) & (x4 | ~x6 | ~x7)));
  assign n1526 = ~n1528 & (n1451 | n1527);
  assign n1527 = x0 ? (x2 | x3) : (~x2 | ~x3);
  assign n1528 = ~x0 & ((~x2 & ~n1529) | (n892 & n876));
  assign n1529 = x3 ? ((x6 | x7 | x4 | ~x5) & (~x6 | ~x7 | ~x4 | x5)) : ((x6 | x7 | x4 | x5) & (~x5 | ((~x6 | ~x7) & (~x4 | x6 | x7))));
  assign n1530 = ~n565 & (n1456 | n1532 | (~x2 & ~n1531));
  assign n1531 = (x1 | (x3 ^ x5) | (x0 ^ ~x4)) & (x0 | x4 | ((x3 | ~x5) & (~x1 | (x3 & ~x5))));
  assign n1532 = ~n976 & (x0 ? (x1 & ~x4) : x4);
  assign n1533 = n1538 & (n1308 | n1537) & (x0 | n1534);
  assign n1534 = (~x1 | x2 | x5 | n1535) & (x1 | (x2 ? n1536 : (~x5 | n1535)));
  assign n1535 = x3 ? (x4 | x6) : (~x4 | ~x6);
  assign n1536 = (x3 | ~x4 | x5 | x6) & (~x3 | ~x5 | (~x4 ^ x6));
  assign n1537 = (~x1 | ((~x3 | ~x4 | ~x0 | x2) & (x3 | x4 | x0 | ~x2))) & (~x0 | x1 | (x2 ? (~x3 | x4) : (x3 | ~x4)));
  assign n1538 = ~n1540 & (n998 | n1542) & (~n363 | n1539);
  assign n1539 = (x2 | ~x3 | x4 | x5 | x6) & (~x2 | x3 | ~x5 | (x4 ^ x6));
  assign n1540 = ~n1541 & (x0 ? (~x2 & x5) : (x2 & ~x5));
  assign n1541 = (x1 | x3 | x4 | ~x6) & (~x1 | (x3 ? (x4 | ~x6) : (~x4 | x6)));
  assign n1542 = (x0 | ~x1 | ~x3 | ~x4 | ~x5) & (~x0 | x5 | (x1 ? (x3 | x4) : (~x3 | ~x4)));
  assign z060 = ~n1552 | ~n1559 | (x3 ? ~n1549 : ~n1544);
  assign n1544 = x2 ? n1547 : (~n1546 & (x5 | n1545));
  assign n1545 = (x0 | x1 | x4 | ~x6 | x7) & (~x0 | ((x6 | x7 | x1 | ~x4) & (~x1 | (x4 ? (x6 | ~x7) : (~x6 | x7)))));
  assign n1546 = n730 & ((n308 & n718) | (~x1 & ~n975));
  assign n1547 = (~n1179 | n1548) & (x0 | ~n313 | ~n910);
  assign n1548 = x0 ? (x1 | x5) : (~x1 | ~x5);
  assign n1549 = ~n1550 & (~n329 | n1551);
  assign n1550 = ~x4 & ((n313 & n428) | (n514 & n921));
  assign n1551 = (~x5 | ((~x1 | ~x2 | ~x6 | ~x7) & (x1 | ((~x6 | x7) & (x2 | x6 | ~x7))))) & (~x1 | ~x2 | x5 | (~x6 ^ x7));
  assign n1552 = x2 ? n1557 : (n1554 & (x1 | n1553));
  assign n1553 = (x0 | ~x3 | (x4 ? (x5 | ~x7) : (~x5 | x7))) & (x3 | ((~x5 | ~x7 | x0 | x4) & (~x0 | ((x5 | ~x7) & (x4 | ~x5 | x7)))));
  assign n1554 = (n1111 | n1556) & (~n1555 | ~n1177);
  assign n1555 = ~x7 & x4 & x5;
  assign n1556 = ~x0 ^ ~x1;
  assign n1557 = (~x0 | x1 | x3 | n574) & (x0 | (x1 ? n1558 : (~x3 | n574)));
  assign n1558 = (~x3 | ~x4 | ~x5 | x7) & (x3 | x4 | x5 | ~x7);
  assign n1559 = ~n1560 & ~n1563 & (n570 | n1562);
  assign n1560 = ~n542 & (x3 ? ~n1561 : (n284 & n300));
  assign n1561 = (x0 | ~x1 | x2 | x4 | ~x5) & (~x0 | x5 | (x1 ? (x2 | ~x4) : (~x2 | x4)));
  assign n1562 = (~x4 | (x0 ? (x1 | ~x3) : (~x1 | x3))) & (~x0 | ((~x1 | ~x2 | x3 | x4) & (x1 | x2 | ~x3))) & (x0 | ~x2 | x4 | (~x1 ^ ~x3));
  assign n1563 = ~n566 & ((~x1 & ~n1564) | (n725 & ~n1565));
  assign n1564 = (~x2 | ~x3 | x4 | x6 | ~x7) & (~x4 | ((x3 | ~x6 | x7) & (x2 | x6 | (~x3 ^ x7))));
  assign n1565 = x3 ? (x4 ? (x6 | ~x7) : (~x6 | x7)) : (x4 | (x6 ^ x7));
  assign z061 = n1579 | ~n1582 | (x1 ? ~n1573 : ~n1567);
  assign n1567 = x0 ? n1568 : (x2 ? n1572 : n1571);
  assign n1568 = x2 ? n1569 : n1570;
  assign n1569 = (x3 | ((x4 | ~x5 | ~x6) & (x7 | (x4 ? (x5 ^ ~x6) : (x5 | x6))))) & (~x3 | ~x4 | x5 | x6 | ~x7) & (x4 | ~x5 | ~x6 | x7);
  assign n1570 = (x3 | ((~x4 | ~x5 | x6 | ~x7) & (~x6 | x7 | x4 | x5))) & (x6 | ~x7 | x4 | x5) & (~x3 | ((~x6 | ~x7 | x4 | ~x5) & (~x4 | (x5 ? (x6 | x7) : (~x6 | ~x7)))));
  assign n1571 = x3 ? ((~x4 | ~x5 | x6 | ~x7) & (~x6 | x7 | x4 | x5)) : ((~x6 | ~x7 | x4 | x5) & (x7 | (x4 ? (x5 ^ x6) : (~x5 | x6))));
  assign n1572 = (~x3 | x4 | ~x5 | ~x6 | ~x7) & ((x3 ^ ~x7) | (x4 ? (x5 ^ ~x6) : (x5 | x6)));
  assign n1573 = n1576 & (n478 | n1575) & (n1254 | n1574);
  assign n1574 = (x0 | ~x2 | x3 | ~x5 | ~x7) & (x2 | ((~x0 | ~x5 | (~x3 ^ x7)) & (x5 | x7 | x0 | x3)));
  assign n1575 = x0 ? (x3 | x5 | (~x4 ^ x6)) : (~x3 | ~x5 | (x4 ^ x6));
  assign n1576 = ~n1577 & (x7 | n998 | ~n669);
  assign n1577 = ~x5 & ((~n485 & ~n1028) | (n659 & ~n1578));
  assign n1578 = (x6 | ~x7 | x2 | ~x4) & (~x2 | x4 | ~x6 | x7);
  assign n1579 = ~x1 & (x7 ? ~n1580 : (n278 & ~n1581));
  assign n1580 = (x0 | x2 | x3 | ~x4 | x6) & (~x3 | ((x0 | x2 | x4 | ~x6) & (~x0 | ~x2 | (x4 ^ x6))));
  assign n1581 = x0 ? (~x3 | ~x6) : (x3 | x6);
  assign n1582 = ~n1584 & n1585 & (n310 | n1583);
  assign n1583 = (x0 | x1 | ~x2 | x4 | ~x6) & ((~x2 ^ x6) | (x0 ? (x1 | x4) : (~x1 | ~x4)));
  assign n1584 = ~n1502 & (n1037 | (n782 & ~n703));
  assign n1585 = (~n295 | ~n1586) & (n645 | n1016 | n1503);
  assign n1586 = x7 & ~x6 & ~x3 & ~x4;
  assign z062 = ~n1592 | ~n1605 | (x2 & ~n1588);
  assign n1588 = ~n1590 & (x1 | ((~n921 | ~n1589) & ~n1591));
  assign n1589 = x4 & ~x0 & ~x3;
  assign n1590 = ~n310 & ((n363 & n458) | (n387 & n301));
  assign n1591 = n760 & ((~x0 & ~x3 & ~x5 & x6) | (x0 & x5 & (x3 ^ x6)));
  assign n1592 = ~n1593 & n1595 & ~n1601 & (n673 | n1604);
  assign n1593 = ~n565 & ((n514 & n1265) | (~x2 & ~n1594));
  assign n1594 = (x0 | ~x1 | x3 | ~x4 | ~x5) & (x4 | ((~x0 | (x1 ? (~x3 | x5) : (x3 | ~x5))) & (x0 | x1 | x3 | x5)));
  assign n1595 = n1598 & (~x0 | ((~n1183 | ~n1127) & ~n1596));
  assign n1596 = ~x1 & ~n1597 & (x2 ? (~x5 & x7) : (~x5 ^ x7));
  assign n1597 = x3 ^ ~x4;
  assign n1598 = x0 ? n1600 : n1599;
  assign n1599 = ((~x2 ^ ~x7) | (x1 ? (~x3 | x5) : (x3 | ~x5))) & (x3 | x5 | (x1 ? (x2 | ~x7) : (~x2 | x7)));
  assign n1600 = (x1 | ~x2 | x3 | ~x5 | x7) & (~x1 | x2 | (x3 ? (~x5 | x7) : (x5 ^ x7)));
  assign n1601 = ~x0 & ((~n1597 & ~n1602) | (x5 & ~n1603));
  assign n1602 = (~x1 | ~x2 | ~x5 | x7) & (x1 | x2 | x5 | ~x7);
  assign n1603 = (~x2 | ((~x4 | x7 | x1 | ~x3) & (x4 | ~x7 | ~x1 | x3))) & (~x1 | x2 | (x3 ? (~x4 | ~x7) : (x4 | x7)));
  assign n1604 = (~x0 | ~x1 | ~x2 | x3 | x7) & (~x3 | (x0 ? (x1 ? (x2 | ~x7) : (~x2 | x7)) : (x1 | (x2 ^ x7))));
  assign n1605 = ~n1606 & (x2 | (~n1608 & (~n1122 | ~n1611)));
  assign n1606 = ~n377 & (x3 ? ~n1607 : (n342 & n514));
  assign n1607 = (x0 | ~x1 | x2 | x4 | ~x7) & (x1 | ((x4 | x7 | x0 | ~x2) & (~x4 | (x0 ? (x2 ^ x7) : (x2 | ~x7)))));
  assign n1608 = ~x3 & (x0 ? ~n1610 : ~n1609);
  assign n1609 = (~x1 | ~x4 | x5 | x6 | x7) & (x1 | x4 | ~x5 | ~x6 | ~x7);
  assign n1610 = (~x1 | ~x4 | ~x5 | x6 | x7) & (x1 | x5 | ((~x6 | ~x7) & (x4 | x6 | x7)));
  assign n1611 = x5 & (x4 ? (x6 & x7) : (~x6 & ~x7));
  assign z063 = ~n1627 | n1623 | n1619 | n1613 | n1616;
  assign n1613 = ~x0 & (x1 ? ~n1614 : ~n1615);
  assign n1614 = x2 ? ((x3 | ~x4 | x5 | ~x6) & (~x3 | x4 | ~x5 | x6)) : (x3 ? (~x4 | x6) : (x4 ? (~x5 | ~x6) : (x5 | x6)));
  assign n1615 = (~x6 | ((~x2 | ~x3 | x4 | ~x5) & (x2 | x5 | (x3 ^ x4)))) & (x3 | x6 | (x2 ? (x4 ^ ~x5) : (~x4 | ~x5)));
  assign n1616 = x0 & (x2 ? ~n1618 : ~n1617);
  assign n1617 = (~x3 | ~x4 | ~x5 | (x1 ^ ~x6)) & (x4 | (x1 ? (x3 ? (x5 | ~x6) : (~x5 | x6)) : (x3 ? (x5 | x6) : ~x6)));
  assign n1618 = (~x1 | x3 | x4 | x5 | x6) & (x1 | ((x5 | x6 | x3 | ~x4) & (~x3 | ~x6 | (x4 ^ ~x5))));
  assign n1619 = ~n565 & (n1621 | ~n1622 | (x2 & ~n1620));
  assign n1620 = (~x0 | ~x1 | x3 | x4 | ~x5) & (x1 | (x3 ? (x4 | x5) : (~x4 | ~x5)));
  assign n1621 = ~x0 & ((x3 & ~x4 & ~x1 & ~x2) | (x1 & x2 & (~x3 ^ x4)));
  assign n1622 = x2 | ((~n356 | ~n480) & (n614 | n1468));
  assign n1623 = ~x2 & (n1624 | n1625 | (~n755 & ~n1626));
  assign n1624 = ~n1597 & ((n480 & n875) | (n441 & n876));
  assign n1625 = ~n542 & ~n954 & (x0 ? n425 : n424);
  assign n1626 = (~x3 | x5 | ~x6 | ~x7) & (x3 | ~x5 | x6 | x7);
  assign n1627 = ~n1628 & (x3 | n1631) & (~n659 | n1632);
  assign n1628 = n438 & (~n1630 | (~n542 & ~n1629));
  assign n1629 = (~x0 | ~x3 | ~x4 | ~x5) & (x0 | x3 | x4 | x5);
  assign n1630 = (x0 | ~x3 | ~x4 | x6 | x7) & (~x0 | x3 | x4 | ~x6 | ~x7);
  assign n1631 = (~n514 | ~n875) & (x7 | ~n399 | n1119);
  assign n1632 = (~x1 | ~x2 | x5 | x6 | x7) & (x1 | ~x6 | ~x7 | (x2 ^ ~x5));
  assign z064 = ~n1643 | (x1 ? ~n1639 : ~n1634);
  assign n1634 = x4 ? n1637 : (x7 ? n1636 : n1635);
  assign n1635 = (~x2 | ((x5 | ~x6 | x0 | ~x3) & (~x0 | (x3 ? (~x5 | ~x6) : (x5 | x6))))) & (x0 | x2 | x5 | (~x3 ^ x6));
  assign n1636 = (~x0 | x2 | x3 | ~x5 | ~x6) & (x0 | ~x3 | x6 | (~x2 ^ x5));
  assign n1637 = (~x7 | n1638) & (~x6 | x7 | ~n339 | n566);
  assign n1638 = (x0 | ~x2 | x3 | x5 | ~x6) & (x6 | ((x0 | ~x2 | ~x3 | ~x5) & (x2 | (x0 ? (x3 ^ ~x5) : (x3 | x5)))));
  assign n1639 = x0 ? (x3 | n1642) : n1640;
  assign n1640 = (x7 | n1641) & (~n624 | n467 | x6 | ~x7);
  assign n1641 = (x2 | ~x3 | ~x4 | x5 | ~x6) & (x3 | ~x5 | (x2 ? (~x4 ^ x6) : (x4 | x6)));
  assign n1642 = (~x2 | x4 | x5 | ~x6 | ~x7) & (x2 | ((~x6 | x7 | x4 | x5) & (x6 | (x4 ? (x5 ^ x7) : (x5 | ~x7)))));
  assign n1643 = n1647 & (n688 | n1646) & (~x0 | n1644);
  assign n1644 = (~x5 | n1645) & (x4 | x5 | x7 | n1516);
  assign n1645 = (x1 | ((~x2 | ~x3 | ~x4 | ~x7) & (x4 | x7 | x2 | x3))) & (~x2 | x3 | x4 | ~x7) & (~x1 | x2 | ~x3 | ~x4 | x7);
  assign n1646 = (x1 | ((x0 | x2 | ~x3 | x5) & (~x0 | (x2 ? x5 : (~x3 | ~x5))))) & (x0 | (x2 ? (x3 | x5) : (~x5 | (~x1 & x3))));
  assign n1647 = ~n1648 & n1651 & (n350 | n1650);
  assign n1648 = ~n542 & (x5 ? ~n1649 : (n380 & ~n1011));
  assign n1649 = (x0 | x1 | x2 | ~x3 | ~x4) & (~x0 | ((x1 | ~x2 | x3 | ~x4) & (~x1 | x2 | ~x3 | x4)));
  assign n1650 = (x0 | ~x1 | x2 | x3 | x5) & ((~x1 ^ ~x3) | (x0 ? (x2 | x5) : (~x2 | ~x5)));
  assign n1651 = (n574 | n1652) & (~n356 | ~n786 | ~n514);
  assign n1652 = (~x0 | ~x1 | x2 | x3) & (x0 | x1 | ~x2 | ~x3);
  assign z065 = ~n1660 | (~x0 & (n1654 | n1657));
  assign n1654 = ~x7 & (x5 ? (~n1011 & ~n1655) : ~n1656);
  assign n1655 = x1 ? (x3 | x6) : (~x3 | ~x6);
  assign n1656 = (x1 | ~x2 | x3 | ~x4 | ~x6) & (~x3 | ((~x1 | (x2 ? (x4 | ~x6) : (~x4 | x6))) & (x1 | x2 | x4 | x6)));
  assign n1657 = x7 & ((n1658 & n971) | (~x2 & ~n1659));
  assign n1658 = x3 & ~x1 & x2;
  assign n1659 = (x1 | ~x3 | ~x4 | x5 | ~x6) & (x3 | (x5 ^ x6) | (~x1 ^ ~x4));
  assign n1660 = ~n1661 & n1666 & n1671 & (n379 | n1665);
  assign n1661 = x0 & ((~x2 & ~n1662) | (n438 & ~n1664));
  assign n1662 = (n1655 | n1663) & (~x6 | ~n314 | ~n762);
  assign n1663 = x4 ? (x5 | x7) : (~x5 | ~x7);
  assign n1664 = (x3 | ~x4 | x5 | ~x6 | ~x7) & (~x5 | ((x3 | x4 | x6 | ~x7) & (~x3 | (x4 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n1665 = x0 ? ((~x3 | ~x4 | x1 | x2) & (~x1 | x3 | x4)) : ((x1 | x3 | ~x4) & (~x3 | (x1 ? (x2 ^ x4) : (~x2 | x4))));
  assign n1666 = ~n1667 & (x0 | (n1669 & (~x1 | n1668)));
  assign n1667 = ~n534 & ((x2 & ~x3 & ~x0 & x1) | (x0 & ~x2 & (x1 ^ ~x3)));
  assign n1668 = (~x2 | ~x3 | x4 | x5 | x6) & (x2 | ~x4 | ~x6 | (~x3 ^ ~x5));
  assign n1669 = (n331 | n1670) & (~n272 | ~n512);
  assign n1670 = (~x3 | ~x4 | ~x5 | x6) & (x3 | x4 | x5 | ~x6);
  assign n1671 = ~n1672 & ((~x1 & ~n1019) | n1674 | (x1 & n836));
  assign n1672 = x0 & (x1 ? (n339 & n320) : ~n1673);
  assign n1673 = (~x3 | x4 | x5 | ~x6) & (x3 | ~x4 | ~x5 | x6) & (~x2 | ((~x5 | ~x6 | x3 | x4) & (~x3 | ~x4 | x5)));
  assign n1674 = (x0 | ~x2 | ~x3 | ~x5 | ~x7) & (x5 | ((~x0 | (x2 ? (x3 | x7) : (~x3 | ~x7))) & (x0 | ~x2 | x3 | ~x7)));
  assign z066 = ~n1688 | (x7 ? (n1682 | ~n1684) : ~n1676);
  assign n1676 = ~n1677 & n1680 & (n388 | n1679);
  assign n1677 = x0 & ((n1114 & n494) | (n423 & ~n1678));
  assign n1678 = (x1 | x4 | x5 | x6) & (~x5 | (x1 ? (~x4 ^ ~x6) : (~x4 | x6)));
  assign n1679 = (x0 | ~x1 | ~x4 | ~x5 | ~x6) & (x5 | ((~x0 | ~x1 | (~x4 ^ x6)) & (x1 | ((~x4 | ~x6) & (x0 | x4 | x6)))));
  assign n1680 = (~n295 | ~n1259) & (n1417 | n1681);
  assign n1681 = (~x4 | x6 | x2 | x3) & (x0 | ((~x2 | x3 | x4 | ~x6) & (x2 | ~x4 | x6)));
  assign n1682 = ~n1548 & (x2 ? (x3 & ~n1254) : n1683);
  assign n1683 = ~x4 & x6;
  assign n1684 = ~n1685 & n1686 & (~n339 | n1254 | n1417);
  assign n1685 = ~x4 & ((n300 & n807) | (n740 & ~n1099));
  assign n1686 = (~n1658 | ~n320) & (~n514 | ~n1687);
  assign n1687 = ~x6 & ~x5 & x3 & x4;
  assign n1688 = ~n1689 & (n1254 | n1693) & (~n408 | n481);
  assign n1689 = x2 & (n1690 | n1691 | (~x0 & ~n1692));
  assign n1690 = n330 & ((n308 & n625) | (~x1 & ~n1262));
  assign n1691 = ~n836 & ((n363 & n403) | (~x0 & ~n369));
  assign n1692 = (~x1 | x3 | ~x4 | x6 | x7) & (x1 | ~x3 | x4 | ~x6 | ~x7);
  assign n1693 = (~x1 | x2 | (x3 ^ x7)) & (~x2 | ((x0 | ~x1 | x3 | ~x7) & (x1 | ~x3 | x7)));
  assign z067 = ~n1696 | ~n1701 | ~n1705 | (~n975 & ~n1695);
  assign n1695 = (~x0 | x1 | ~x2 | x3 | ~x5) & (x0 | ((x2 | ~x3 | x5) & (~x1 | ~x2 | x3 | ~x5)));
  assign n1696 = n1698 & (n377 | ((~n364 | ~n889) & ~n1697));
  assign n1697 = ~n470 & ((n426 & n1074) | (n423 & n760));
  assign n1698 = ~n1700 & (x0 | n1699) & (n570 | n1235);
  assign n1699 = (~x2 | ~x3 | ~x5 | x7) & (x2 | x3 | x5 | ~x7);
  assign n1700 = x7 & ~x5 & ~x3 & x0 & ~x2;
  assign n1701 = ~n1703 & (n379 | (~n1702 & (~n364 | ~n890)));
  assign n1702 = ~n470 & ((n340 & n760) | (n339 & n1074));
  assign n1703 = n342 & ((n514 & n1704) | (n399 & ~n1116));
  assign n1704 = x6 & x3 & ~x5;
  assign n1705 = n1709 & (~n1706 | ~n1708) & (~n857 | n1707);
  assign n1706 = ~x3 & ~x0 & ~x1;
  assign n1707 = (~x1 | x2 | x4 | x5 | x7) & (x1 | ~x2 | ((~x4 | x5 | ~x7) & (~x5 | x7)));
  assign n1708 = x4 & x5 & x7 & (x2 ^ ~x6);
  assign n1709 = (n481 | n1711) & (x0 | n1710);
  assign n1710 = (x1 | x2 | x3 | ~n886) & (~x1 | ~x2 | ~x3 | ~n629);
  assign n1711 = (x0 | x1 | ~x2 | ~x3 | x5) & (x2 | x3 | ~x5 | (~x0 & ~x1));
  assign z068 = (x3 | ~n1713) & (n1722 | n1724 | ~x3 | ~n1718);
  assign n1713 = ~n1714 & ~n1715 & n1716 & (x1 | n551);
  assign n1714 = ~x0 & ((~x4 & ~x5 & x6) | (x1 & x4 & x5 & ~x6));
  assign n1715 = ~n542 & ((~x0 & x4 & ~x5) | (~x4 & x5 & (x0 | n387)));
  assign n1716 = (n1717 | n485) & (~n320 | (~n363 & ~n364));
  assign n1717 = x0 ? x5 : (x1 | ~x5);
  assign n1718 = ~n1719 & ~n1721 & (n602 | (x0 & ~n428));
  assign n1719 = ~n565 & ~n1720;
  assign n1720 = (~x4 & ~x5 & (~x0 | (~x1 & ~x2))) | (x4 & x5) | (x0 & x1 & x2);
  assign n1721 = n559 & ~n271 & x5 & x6;
  assign n1722 = ~x1 & (~n1723 | (x0 & n624 & n876));
  assign n1723 = (~x0 | ~x4 | x5 | ~x6 | ~x7) & (x0 | x4 | ~x5 | x6 | x7);
  assign n1724 = n1494 & ((n782 & n1370) | (n647 & ~n975));
  assign z069 = ~n1730 | (~x7 & ~n836 & ~n1729) | (x7 & ~n1726);
  assign n1726 = x0 ? (x5 | n1728) : n1727;
  assign n1727 = (x1 | x2 | x3 | ~n512) & (~x1 | ~x2 | ~x3 | ~n971);
  assign n1728 = (~x4 & x6) | (x4 & ~x6) | (x1 & x2 & (x3 | x6));
  assign n1729 = x0 ? (x5 | (x1 ^ (~x2 | ~x3))) : (x1 | ~x5);
  assign n1730 = (n1731 | ~n1734) & (x5 | n1733) & (~x5 | n1732);
  assign n1731 = x1 ? (x4 | ~x5) : (~x4 | x5);
  assign n1732 = (~x7 & (x4 | (~x0 & ~x1))) | (~x4 & x7) | (x0 & x1 & x2);
  assign n1733 = (~x4 | x7 | x1 | x2) & (x0 | (~x4 ^ x7));
  assign n1734 = ~x7 & ~x3 & x0 & x2;
  assign z070 = ~n1736 | n1744 | (~x1 & ~n1742);
  assign n1736 = ~n1738 & ~n1739 & n1740 & (x1 | n1737);
  assign n1737 = x0 ? (~x6 | ((x5 | ~x7) & (x2 | ~x5 | x7))) : (~x2 | x6 | (x5 ^ x7));
  assign n1738 = x5 & ((~x6 & (x1 ? (~x0 | ~x2) : x0)) | (~x0 & (~x1 | ~x2) & x6));
  assign n1739 = ~n614 & n340 & n387 & x6 & x7;
  assign n1740 = ~n1741 & (~n514 | (~n556 & (~n717 | ~n314)));
  assign n1741 = x6 & ~x5 & ~x2 & x0 & x1;
  assign n1742 = (x7 | n1743) & (~n579 | n498 | x6 | ~x7);
  assign n1743 = (x0 | x2 | ~x3 | x5 | x6) & (~x0 | ~x2 | ~x6 | (x3 ^ ~x5));
  assign n1744 = ~x3 & ((n273 & n1747) | (~x6 & ~n1745));
  assign n1745 = (~x4 | n570 | ~n1241) & (~x1 | x4 | n1746);
  assign n1746 = (~x0 | ~x2 | ~x5) & (x0 | x2 | x5 | x7);
  assign n1747 = x2 & x0 & x1;
  assign z071 = n1749 | ~n1754 | (x1 & (~n1762 | ~n1763));
  assign n1749 = ~x0 & (n1751 | (n1295 & ~n565 & ~n1750));
  assign n1750 = ~x4 & ~x2 & ~x3;
  assign n1751 = ~x5 & (x7 ? ~n1753 : (n1752 & ~n1750));
  assign n1752 = ~x1 & x6;
  assign n1753 = x1 ? ((~x2 | ~x3 | ~x4 | ~x6) & (x4 | x6 | x2 | x3)) : (x6 | (~x2 & ~x3));
  assign n1754 = ~n1756 & ~n1758 & n1760 & (~n990 | ~n1755);
  assign n1755 = ~x7 & ~x6 & ~x4 & ~x5;
  assign n1756 = ~n542 & ((n514 & n612) | (n363 & ~n1757));
  assign n1757 = x2 & x3;
  assign n1758 = ~n1759 & ~x6 & n387;
  assign n1759 = (~x2 | ~x3 | ~x4 | x5) & (x2 | x3 | x4 | ~x5);
  assign n1760 = x1 | (x0 ? (~x2 | ~n519) : (x2 | ~n1761));
  assign n1761 = x6 & ~x3 & ~x4;
  assign n1762 = x0 ? (x2 | ~x6) : (x6 | (x2 ^ ~x3));
  assign n1763 = (~x0 | ~x2 | x3 | x4 | ~x6) & (x0 | x6 | (x2 ? (~x3 | x4) : (x3 | ~x4)));
  assign z072 = ~n1770 | (~x5 & (x4 ? ~n1767 : ~n1765));
  assign n1765 = (n565 | (~n990 & ~n1014)) & (~n359 | ~n1766);
  assign n1766 = ~x7 & ~x3 & x6;
  assign n1767 = x0 ? (~n282 | ~n1768) : n1769;
  assign n1768 = ~x7 & ~x3 & ~x6;
  assign n1769 = (x1 | x2 | x3 | ~x6 | ~x7) & (~x1 | ~x2 | ~x3 | (x6 ^ x7));
  assign n1770 = ~n1771 & ~n1774 & n1775 & (x7 | n1773);
  assign n1771 = ~x0 & ((n269 & n1422) | (x5 & ~n1772));
  assign n1772 = (~x1 | ~x2 | ~x3 | ~x4 | ~x7) & (x2 | x3 | ((x4 | x7) & (x1 | ~x4 | ~x7)));
  assign n1773 = (x0 | ~x1 | x2 | x3 | ~x4) & (~x2 | ((x0 | ~x1 | ~x3 | x4) & (~x0 | (x1 ? (x3 | x4) : (~x3 | ~x4)))));
  assign n1774 = ~x0 & ((x3 & x7 & ~x1 & ~x2) | (x1 & ~x7 & (~x2 ^ ~x3)));
  assign n1775 = n1776 & ~n1777 & (~n790 | ~n443 | ~n394);
  assign n1776 = (x0 | x1 | ~x2 | ~x7) & (~x0 | x2 | (~x1 ^ x7));
  assign n1777 = x7 & ~x3 & x2 & x0 & ~x1;
  assign z073 = n1781 | ~n1783 | (x0 ? ~n1780 : ~n1779);
  assign n1779 = (x1 | ((x2 | ~x4 | ~x5) & (x4 | x5 | ~x2 | x3))) & (~x1 | ~x2 | ~x3 | ~x4 | ~x5) & (x2 | ((~x1 | (~x4 ^ x5)) & (x3 | ~x4 | ~x5) & (~x3 | (x4 & x5))));
  assign n1780 = (x1 & (x3 | (x4 & x5))) | (x2 & (~x3 | (~x4 & ~x5))) | (~x2 & x3 & (x4 | x5));
  assign n1781 = ~x3 & ((n320 & n364) | (n601 & ~n1782));
  assign n1782 = (~x5 | x6 | x1 | ~x2) & (~x1 | x2 | x5 | ~x6);
  assign n1783 = (~x3 | ~n1033) & (x3 | ~x6 | ~n441 | n1784);
  assign n1784 = (x5 | ~x7 | x2 | ~x4) & (~x2 | x4 | ~x5 | x7);
  assign z074 = ~n1788 | ~n1793 | (x2 ? ~n1786 : ~n1787);
  assign n1786 = (x0 | x1 | ~x3 | x4 | x5) & ((x3 ^ x5) | (x0 ? (x1 | x4) : (~x1 | ~x4)));
  assign n1787 = (~x0 | ~x1 | ~x3 | ~x4 | x5) & (x0 | x3 | ~x5 | (~x1 ^ x4));
  assign n1788 = (~x6 | n1789) & (~n441 | n1791);
  assign n1789 = x3 ? (n1091 | n1034) : (~n725 | n1790);
  assign n1790 = x0 ? (~x4 | ~x5) : (x4 | x5);
  assign n1791 = x5 ? (~n717 | ~n892) : (~n1207 | n1792);
  assign n1792 = x3 ? (x6 | x7) : (~x6 | ~x7);
  assign n1793 = x0 ? ((~x1 | x2 | ~x3 | x4) & (x1 | ((~x3 | ~x4) & (x2 | x3 | x4)))) : ((~x3 | x4 | x1 | x2) & (x3 | (x1 ? (~x2 ^ x4) : (~x2 | ~x4))));
  assign z075 = n1795 | ~n1800 | n1810 | (~n1091 & ~n1809);
  assign n1795 = ~x4 & (n1796 | (n387 & n519 & n1799));
  assign n1796 = ~x3 & (x5 ? (n782 & ~n1798) : ~n1797);
  assign n1797 = (x0 | x1 | x2 | x6 | ~x7) & (~x0 | x7 | (x1 ? (~x2 | ~x6) : (x2 | x6)));
  assign n1798 = x1 ? (x6 | x7) : (~x6 | ~x7);
  assign n1799 = ~x7 & (~x2 ^ ~x5);
  assign n1800 = ~n1802 & ~n1804 & n1805 & (x0 | n1801);
  assign n1801 = (~x1 | x2 | x4 | (~x3 ^ x5)) & (~x2 | ((x4 | x5 | ~x1 | x3) & (x1 | (x3 ? (x4 | ~x5) : (~x4 | x5)))));
  assign n1802 = ~n1163 & ((n359 & n629) | (n744 & ~n1803));
  assign n1803 = (~x1 | x2 | x4 | ~x5) & (x1 | ~x4 | (~x2 ^ x5));
  assign n1804 = x4 & ((~x0 & x5 & (~x1 ^ x2)) | (x0 & ~x1 & ~x2 & ~x5));
  assign n1805 = n1806 & ~n1807 & (~n329 | ~n450 | n1808);
  assign n1806 = (~n364 | ~n612) & (~n330 | n1119);
  assign n1807 = ~n467 & n441 & ~x6 & n278;
  assign n1808 = (x1 | ~x2 | ~x3 | ~x6) & (~x1 | x2 | x3 | x6);
  assign n1809 = (~x1 | ((x4 | x6 | ~x0 | x3) & (x0 | ~x3 | (x4 ^ x6)))) & (~x0 | x1 | (x3 ? (x4 | ~x6) : (~x4 | x6)));
  assign n1810 = ~x2 & ((n458 & n1063) | (x6 & ~n1811));
  assign n1811 = (~x0 | ~x1 | x3 | ~x4 | ~x5) & (x0 | x5 | ((x3 | x4) & (x1 | ~x3 | ~x4)));
  assign z076 = n1813 | ~n1818 | ~n1822 | (~n1291 & ~n1816);
  assign n1813 = x1 & ((x5 & ~n1814) | (n924 & ~n1815));
  assign n1814 = (x0 | x2 | ~x3 | ~x4 | ~x6) & (x6 | (x0 ? (x2 ? (x3 | x4) : (~x3 | ~x4)) : (x3 | (~x2 ^ ~x4))));
  assign n1815 = (x4 | ~x6 | x2 | ~x3) & (~x2 | (x3 ? (~x4 | ~x6) : (x4 | x6)));
  assign n1816 = (~x0 | x3 | ~n408 | ~n1019) & (x0 | n1817);
  assign n1817 = (x1 | ~x2 | ~x3 | ~x4 | ~x6) & (~x1 | ((~x2 | ~x3 | x4 | ~x6) & (~x4 | x6 | x2 | x3)));
  assign n1818 = (~x1 | n1821) & (x1 | n1820) & (n1597 | n1819);
  assign n1819 = (x0 | x1 | ~x2 | ~x5 | ~x6) & (~x0 | x2 | (x1 ? (~x5 | ~x6) : (x5 | x6)));
  assign n1820 = ((~x0 ^ ~x2) | (x3 ? (x5 | ~x6) : (~x5 | x6))) & ((x3 ^ x5) | (x0 ? (x2 | ~x6) : (~x2 | x6)));
  assign n1821 = (~x0 | x2 | x3 | x5 | x6) & (x0 | (~x2 ^ ~x5) | (~x3 ^ x6));
  assign n1822 = x0 ? (n1827 & (n1163 | n1826)) : n1823;
  assign n1823 = x1 ? (n881 | n1663) : (~n1824 & ~n1825);
  assign n1824 = n892 & n875;
  assign n1825 = ~n1163 & ((n624 & n450) | (~x2 & ~n574));
  assign n1826 = (x1 | ~x2 | (x4 ? (x5 | ~x7) : (~x5 | x7))) & (x2 | ((~x5 | ~x7 | x1 | ~x4) & (~x1 | x4 | (x5 ^ x7))));
  assign n1827 = (~n272 | ~n411) & (n573 | ~n1168);
  assign z077 = ~n1833 | (x0 & (n1829 | (n438 & ~n1832)));
  assign n1829 = ~x2 & (x5 ? ~n1830 : ~n1831);
  assign n1830 = x1 ? ((~x3 | x4 | x6 | ~x7) & (x3 | ~x4 | ~x6 | x7)) : ((~x3 | ~x4 | (~x6 ^ x7)) & (x6 | ~x7 | x3 | x4));
  assign n1831 = (x1 | ~x3 | x4 | x6 | x7) & ((~x6 ^ x7) | (x1 ? (~x3 | x4) : (x3 ^ x4)));
  assign n1832 = (~x3 | ~x4 | x5 | (~x6 ^ x7)) & (~x5 | ((x6 | x7 | x3 | ~x4) & (x4 | (x3 ? (~x6 ^ x7) : (~x6 | ~x7)))));
  assign n1833 = n1843 & (n542 | n1840) & (x0 | n1834);
  assign n1834 = ~n1835 & ~n1836 & ~n1838 & (~x6 | n1839);
  assign n1835 = ~n1516 & ((x4 & ~x5 & ~x6 & x7) | (~x4 & ((x6 & ~x7) | (x5 & ~x6 & x7))));
  assign n1836 = n1837 & ((n1369 & ~n1193) | (n276 & n1183));
  assign n1837 = ~x2 & ~x6;
  assign n1838 = ~n565 & (x1 ? (~x2 & n356) : (x2 & n1270));
  assign n1839 = (~n1658 | ~n629) & (~x5 | n954 | n1279);
  assign n1840 = ~n1842 & (x2 ? n1841 : (~n606 | ~n480));
  assign n1841 = (x0 | x1 | ~x3 | ~x4 | ~x5) & (~x0 | x3 | x5 | (~x1 ^ x4));
  assign n1842 = ~n954 & ((x0 & ~x2 & x4 & x5) | (~x0 & (x2 ? ~x4 : (x4 & ~x5))));
  assign n1843 = ~n1844 & n1847 & (n1163 | n1846);
  assign n1844 = ~x1 & ((~x4 & ~n1845) | (n764 & n661));
  assign n1845 = x0 ? (x5 | (x2 ? (x3 | x6) : (~x3 | ~x6))) : (~x5 | x6 | (x2 ^ x3));
  assign n1846 = (x0 | ~x1 | x2 | x4) & (~x4 | (x0 ? (x1 ? (x2 | x5) : (~x2 | ~x5)) : (x1 | (~x2 ^ x5))));
  assign n1847 = (n1034 | n1848) & (~n327 | ~n606 | ~n742);
  assign n1848 = (x2 | ~x3 | ~x5 | ~x6) & (~x2 | (x3 ? (x5 | ~x6) : (~x5 | x6)));
  assign z078 = ~n1865 | n1860 | n1857 | n1850 | n1854;
  assign n1850 = x1 & (n712 | n1852 | (~n1851 & ~n1527));
  assign n1851 = (~x4 | ~x5 | ~x6 | ~x7) & (x4 | x5 | x6 | x7);
  assign n1852 = ~x0 & ((~x6 & ~n1853) | (n280 & n974));
  assign n1853 = (x2 | ~x3 | x4 | ~x5 | x7) & (~x4 | ((x2 | x3 | ~x5 | ~x7) & (~x2 | (x3 ? (~x5 | x7) : (x5 | ~x7)))));
  assign n1854 = ~x4 & ((n441 & ~n1856) | (x0 & ~n1855));
  assign n1855 = (x5 | ~x7 | x2 | x3) & (x7 | ((x1 | ~x3 | (~x2 ^ x5)) & (~x1 | ~x2 | x3 | ~x5)));
  assign n1856 = x2 ? ((x5 | ~x7) & (~x3 | ~x5 | x7)) : (~x3 | (x5 ^ x7));
  assign n1857 = ~n688 & (x1 ? ~n1859 : ~n1858);
  assign n1858 = x0 ? ((x5 | x6 | x2 | ~x3) & (~x5 | ~x6 | ~x2 | x3)) : ((x2 | ~x3 | x5 | ~x6) & (~x2 | x3 | ~x5 | x6));
  assign n1859 = (x0 | x2 | ~x3 | ~x5 | ~x6) & (x3 | x5 | (x0 ? (~x2 | x6) : (~x2 ^ ~x6)));
  assign n1860 = ~x1 & (x6 ? ~n1862 : (~n1436 & ~n1861));
  assign n1861 = (x3 | x4 | ~x5 | x7) & (~x3 | ~x4 | x5 | ~x7);
  assign n1862 = x3 ? (x5 | n1864) : ((~n579 | ~n1863) & (~x5 | n1864));
  assign n1863 = ~x4 & (~x5 ^ x7);
  assign n1864 = (x0 | ~x2 | ~x4 | ~x7) & (~x0 | x2 | x4 | x7);
  assign n1865 = ~n1869 & (n467 | n1868) & (~x4 | n1866);
  assign n1866 = (x1 | n1867) & (x2 | ~n789 | x0 | ~x1);
  assign n1867 = (~x2 | ((~x0 | (x3 ? (~x5 | x7) : (x5 | ~x7))) & (x5 | x7 | x0 | ~x3))) & (x0 | x2 | ((~x5 | x7) & (x3 | x5 | ~x7)));
  assign n1868 = (~x0 | x1 | x2 | ~x4 | ~x7) & (~x1 | ((x4 | x7 | x0 | x2) & ((~x4 ^ x7) | (x0 ^ ~x2))));
  assign n1869 = ~n1870 & (x0 ? ((~x2 & x4) | (~x1 & x2 & ~x4)) : (x2 & (x1 ^ x4)));
  assign n1870 = x3 ? (~x5 | ~x7) : (x5 | x7);
  assign z079 = ~n1883 | (x0 ? ~n1872 : ~n1877);
  assign n1872 = ~n1875 & (~x6 | (x1 & n1874) | (~x1 & n1873));
  assign n1873 = (x2 | x3 | ~x4 | ~x5 | x7) & (~x2 | ((x5 | x7 | x3 | x4) & (~x3 | (x4 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n1874 = (~x2 | x3 | x4 | x5 | ~x7) & (x2 | ~x4 | (x3 ? (~x5 | x7) : (x5 ^ x7)));
  assign n1875 = n1837 & ((n718 & n1876) | (~n1318 & ~n989));
  assign n1876 = x7 & (x3 ^ ~x5);
  assign n1877 = x7 ? (x5 ? n1878 : n1879) : n1880;
  assign n1878 = (~x1 | x2 | ~x3 | ~x4 | x6) & (x1 | ~x2 | x3 | x4 | ~x6);
  assign n1879 = x4 ? ((~x3 | ~x6 | x1 | ~x2) & (~x1 | x2 | x3 | x6)) : (x1 ? (~x2 | (~x3 ^ x6)) : (x2 | (x3 ^ x6)));
  assign n1880 = (~x2 | ~x6 | n1881) & (x6 | (n1882 & (x2 | n1881)));
  assign n1881 = (x1 | ~x3 | ~x4 | ~x5) & (~x1 | (x3 ? (~x4 | x5) : (x4 | ~x5)));
  assign n1882 = (~x1 | ~x2 | x3 | ~x4 | ~x5) & (x1 | x5 | (x2 ? (~x3 | x4) : (x3 | ~x4)));
  assign n1883 = n1886 & (n836 | n1885) & (n498 | n1884);
  assign n1884 = (x6 | ((x1 | ~x2) & (~x0 | (x1 ? (x2 | ~x4) : x4)))) & (~x1 | x2 | x4 | ~x6) & (x0 | (x1 ? (~x4 | ~x6) : (~x2 | x4)));
  assign n1885 = (x0 | ~x1 | ~x2 | ~x3 | x5) & (x3 | ~x5 | x1 | x2);
  assign n1886 = ~n1887 & ~n1888 & (~x5 | n1535 | ~n1241);
  assign n1887 = ~n976 & (~n770 | (n1683 & n363));
  assign n1888 = ~n1889 & ((n356 & n786) | (n443 & n450));
  assign n1889 = (x2 | ~x6 | x0 | ~x1) & (~x0 | x1 | ~x2 | x6);
  assign z080 = n1908 | n1904 | n1902 | ~n1891 | n1899;
  assign n1891 = n1894 & (n350 | n1893) & (n565 | n1892);
  assign n1892 = x2 ? (~n387 | n766) : (n1274 | n1731);
  assign n1893 = (x0 | x1 | ~x3 | n903) & (~x0 | x3 | n1782);
  assign n1894 = n1898 & (x2 | (n1895 & (n1896 | n1897)));
  assign n1895 = (~x0 | x3 | ~x4 | x5 | x6) & (x0 | ~x3 | x4 | ~x5 | ~x6) & ((~x0 ^ ~x3) | (x4 ? (~x5 | x6) : (x5 | ~x6)));
  assign n1896 = x0 ? (x3 | x4) : (~x3 | ~x4);
  assign n1897 = x1 ? (x6 | ~x7) : (~x6 | x7);
  assign n1898 = (~n594 | ~n1145) & (~n521 | ~n356 | ~n394);
  assign n1899 = ~n542 & (n1900 | n1901 | (n579 & n1270));
  assign n1900 = ~x3 & ((~x0 & x2 & ~x4 & x5) | (x0 & (x2 ? (~x4 & ~x5) : (x4 & x5))));
  assign n1901 = x4 & n340 & (x0 ? (~x1 & ~x5) : (x1 ^ x5));
  assign n1902 = ~n379 & (x4 ? ~n1903 : (~n847 & n1122));
  assign n1903 = (~x0 | ~x1 | x2 | ~x3 | ~x7) & (x0 | x3 | (x1 ? (x2 | ~x7) : (~x2 | x7)));
  assign n1904 = x2 & ((n764 & n1063) | n1905 | n1906);
  assign n1905 = ~n1254 & ((x0 & ~x1 & x3 & x5) | (~x0 & ((x1 & x3 & x5) | (~x3 & ~x5))));
  assign n1906 = n424 & (n1907 | (x0 & n709));
  assign n1907 = ~x6 & x3 & ~x0 & ~x1;
  assign n1908 = ~x0 & (n1910 | (n620 & n1074 & ~n1909));
  assign n1909 = x2 ? (~x5 | x6) : (x5 | ~x6);
  assign n1910 = ~x4 & (x1 ? (n426 & n313) : ~n1911);
  assign n1911 = (x2 | x3 | ~x5 | ~x6 | x7) & (~x2 | ~x3 | x5 | x6 | ~x7);
  assign z081 = ~n1913 | n1925 | ~n1928 | (x1 & ~n1922);
  assign n1913 = ~n1914 & ~n1917 & (n310 | n1916);
  assign n1914 = ~x0 & (x6 ? (n588 & ~n1188) : ~n1915);
  assign n1915 = x1 ? ((~x3 | x4 | x5 | ~x7) & (x3 | ~x4 | ~x5 | x7)) : (x3 | (x4 ? (x5 | ~x7) : (~x5 | x7)));
  assign n1916 = (x0 | ~x1 | x4 | ~x5) & (~x0 | ((~x4 | ~x5 | x1 | ~x2) & (~x1 | x2 | (x4 ^ x5))));
  assign n1917 = ~x1 & (n1919 | n1920 | (~x2 & ~n1918));
  assign n1918 = (~x0 | ~x3 | x4 | ~x5 | x7) & (x0 | ((~x3 | x4 | x5 | ~x7) & (x3 | ~x4 | ~x5 | x7)));
  assign n1919 = ~n570 & ((n647 & n356) | (~x0 & ~n1235));
  assign n1920 = n426 & ((n1921 & ~n688) | (n790 & n329));
  assign n1921 = x0 & ~x5;
  assign n1922 = (~x7 | n1923) & (x5 | x7 | ~n285 | n1924);
  assign n1923 = (~x0 | x2 | ~x3 | x4 | ~x5) & (x0 | ~x4 | ((~x3 | x5) & (~x2 | x3 | ~x5)));
  assign n1924 = ~x2 & x4;
  assign n1925 = x6 & ((n514 & n1473) | n1926);
  assign n1926 = ~x2 & ((~n570 & ~n1927) | (n886 & n1063));
  assign n1927 = (~x0 | ~x1 | ~x3 | ~x4) & (x0 | x1 | x3 | x4);
  assign n1928 = ~n1929 & (n1291 | n1931) & (~x0 | n1932);
  assign n1929 = ~n1163 & (n1930 | (~n271 & n329 & ~n570));
  assign n1930 = x0 & ((~n271 & ~n574) | (n408 & n1183));
  assign n1931 = (~x0 | ((~x3 | ~x4 | x1 | x2) & (~x1 | ~x2 | x3 | x4))) & (x0 | x1 | ~x2 | ~x3 | x4);
  assign n1932 = (n570 | ~n473 | n506) & (~n1933 | ~n876);
  assign n1933 = x4 & x1 & ~x3;
  assign z082 = n1947 | ~n1949 | (x3 ? ~n1935 : ~n1940);
  assign n1935 = ~n1936 & ~n1938;
  assign n1936 = ~x2 & (x1 ? (~n542 & ~n1790) : ~n1937);
  assign n1937 = x0 ? ((~x6 | ~x7 | x4 | ~x5) & (x6 | x7 | ~x4 | x5)) : (x4 ? (x5 ? (x6 | x7) : (~x6 | ~x7)) : (x5 ? (x6 | ~x7) : (~x6 | x7)));
  assign n1938 = x2 & (x0 ? (n313 & n913) : ~n1939);
  assign n1939 = (x1 | ~x4 | ~x5 | ~x6 | ~x7) & (x4 | ((~x6 | x7 | x1 | ~x5) & (~x1 | (x5 ? (x6 | x7) : (~x6 | ~x7)))));
  assign n1940 = x1 ? n1943 : (x4 ? n1941 : n1942);
  assign n1941 = (~x6 | (x0 ? (x2 ? (x5 | ~x7) : (~x5 | x7)) : (~x7 | (x2 ^ x5)))) & (~x2 | x6 | x7 | (x0 ^ ~x5));
  assign n1942 = (~x0 | x2 | ~x5 | ~x6 | ~x7) & (x6 | ((~x5 | ~x7 | x0 | ~x2) & (~x0 | (x2 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n1943 = ~n1946 & (n605 | n1945) & (~n579 | ~n1944);
  assign n1944 = ~x4 & ~x7 & (~x5 ^ x6);
  assign n1945 = (x6 | ~x7 | x0 | ~x4) & (~x0 | x4 | ~x6 | x7);
  assign n1946 = ~n688 & ((n587 & n782) | (n647 & n1039));
  assign n1947 = ~n565 & (x3 ? ~n1948 : (n335 & n359));
  assign n1948 = x0 ? (x4 | (x1 ? (x2 | ~x5) : (~x2 | x5))) : (~x1 | ~x4 | (x2 ^ x5));
  assign n1949 = n1954 & (x6 ? (~n473 | n1953) : n1950);
  assign n1950 = ~n1952 & (~x2 | n1951);
  assign n1951 = (x0 | ~x1 | ~x3 | ~x4 | x5) & (~x0 | ((x1 | ~x4 | ~x5) & (x4 | x5 | ~x1 | x3)));
  assign n1952 = n408 & ((~x0 & x3 & ~x4 & ~x5) | (x4 & ((~x3 & x5) | (x0 & (~x3 | x5)))));
  assign n1953 = (~x0 & (x3 | ~x5)) | (x0 & ~x2 & x5) | (x2 & x3 & ~x5);
  assign n1954 = (n998 | n1956) & (n1254 | n1955);
  assign n1955 = (x0 | x1 | ~x2 | x5) & (~x1 | (x0 ? (x2 | x5) : (~x5 | (x2 & x3))));
  assign n1956 = (~x0 | ~x1 | x3 | x4 | ~x5) & (x0 | ((x1 | ~x3 | x4 | ~x5) & (~x1 | x3 | ~x4 | x5)));
  assign z083 = n1958 | ~n1968 | (~n570 & ~n1961);
  assign n1958 = x3 & ((n364 & n430) | n1959);
  assign n1959 = ~x1 & (x4 ? (n647 & ~n563) : ~n1960);
  assign n1960 = (x0 | x2 | ~x5 | ~x6 | x7) & (x6 | ((x0 | (x2 ? (~x5 | x7) : (x5 | ~x7))) & (~x0 | ~x2 | x5 | ~x7)));
  assign n1961 = ~n1963 & ~n1965 & n1966 & (x2 | n1962);
  assign n1962 = x0 ? ((~x4 | ~x6 | x1 | ~x3) & (~x1 | x3 | x6)) : (x4 | (x1 ? (x3 | ~x6) : (~x3 | x6)));
  assign n1963 = n782 & (x1 ? (x3 & n1019) : (x3 ? n1964 : n1019));
  assign n1964 = x4 & x6;
  assign n1965 = ~x1 & (x0 ? (~x2 & ~x3) : (x2 & (x3 ^ x4)));
  assign n1966 = ~n1967 & (n1516 | (x0 ? (x4 | ~x6) : (~x4 | x6)));
  assign n1967 = x1 & x3 & (x0 ? ~x2 : (x2 & x4));
  assign n1968 = ~n1969 & ~n1972 & n1976 & (n1291 | n1971);
  assign n1969 = ~x3 & ((n296 & n428) | (~n1291 & ~n1970));
  assign n1970 = (x0 | x1 | x2 | x4 | x6) & (~x0 | ~x6 | (x1 ? (x2 | x4) : (~x2 | ~x4)));
  assign n1971 = (x1 | ((x0 | x2 | x3 | ~x6) & (~x0 | ~x2 | (x3 ^ x6)))) & (x0 | ~x1 | (x2 ^ (~x3 & x6)));
  assign n1972 = x4 & ((n359 & n1973) | (~n1974 & ~n1975));
  assign n1973 = ~x6 & ~x3 & ~x5;
  assign n1974 = x0 ^ ~x5;
  assign n1975 = (~x3 | x6 | x1 | ~x2) & (~x1 | x2 | x3 | ~x6);
  assign n1976 = (n566 | ~n1383 | n1977) & (~x3 | n1978);
  assign n1977 = x1 ^ ~x6;
  assign n1978 = (~n428 | ~n921) & (~n1979 | (~x1 ^ ~x2));
  assign n1979 = x7 & x6 & ~x0 & ~x5;
  assign z084 = ~n1990 | n1988 | n1987 | n1981 | ~n1983;
  assign n1981 = ~n565 & (x1 ? ~n1982 : n892);
  assign n1982 = (~x4 | ~x5 | x2 | x3) & (~x3 | ((x0 | ~x2 | (~x4 ^ x5)) & (x4 | x5 | ~x0 | x2)));
  assign n1983 = n1985 & (x3 | n1984);
  assign n1984 = x1 ? (x6 | ((x2 | x4) & (x0 | ~x2 | ~x4))) : (~x6 | (x2 ^ x4));
  assign n1985 = (~n1986 | ~n764) & (x4 | ~n923 | n903);
  assign n1986 = ~x3 & x1 & ~x2;
  assign n1987 = n423 & (x1 ? (x6 & (x0 ^ ~x4)) : (x4 & ~x6));
  assign n1988 = x3 & (n1989 | (n284 & ~n998 & ~n779));
  assign n1989 = ~n1486 & n579 & ~x6 & n335;
  assign n1990 = ~n1993 & (n1991 | ~n1992) & (~n620 | n1996);
  assign n1991 = (~x0 | ((~x6 | ~x7 | x1 | x2) & (~x1 | ~x2 | x6 | x7))) & (~x1 | x2 | ~x6 | x7);
  assign n1992 = ~x5 & ~x3 & x4;
  assign n1993 = ~n542 & ((~x3 & ~n1994) | (n923 & ~n1995));
  assign n1994 = x1 ? (~x2 | x4) : (x2 | ~x4 | (x0 & ~x5));
  assign n1995 = (~x0 | x2 | x4 | x5) & (~x2 | (x4 ^ ~x5));
  assign n1996 = (~x0 | x2 | x4 | ~x5 | ~x6) & (x0 | ((x2 | ~x4 | x5 | ~x6) & (~x2 | (x4 ? (~x5 | ~x6) : (x5 | x6)))));
  assign z085 = n1998 | ~n2002 | ~n2009 | (x2 & ~n2001);
  assign n1998 = ~x7 & ((~n470 & n1999) | (~x5 & ~n2000));
  assign n1999 = x5 & ~x4 & x2 & x3;
  assign n2000 = x3 ? ((x2 | x4) & (x0 | ~x2 | ~x4)) : ((~x0 | x1 | ~x2 | x4) & (x0 | (x1 ? (~x2 | x4) : (x2 | ~x4))));
  assign n2001 = (x7 | ((~x0 | (x1 ? (x3 | x4) : (~x3 | ~x4))) & (x0 | x1 | x3 | x4))) & (x3 | ~x4 | ~x7 | (x0 & x1));
  assign n2002 = n2005 & (n998 | ((~n1183 | ~n1063) & ~n2003));
  assign n2003 = n1074 & (~n2004 | (n387 & n465));
  assign n2004 = x0 ? (x3 | x5) : (~x3 | ~x5);
  assign n2005 = ~n2008 & (~n423 | ~n2007) & (x2 | ~n2006);
  assign n2006 = x7 & ~x3 & ~x4;
  assign n2007 = x7 & ~x4 & x5;
  assign n2008 = ~n453 & ((~n736 & ~n1331) | (n1207 & ~n1556));
  assign n2009 = ~n2011 & (x0 | ((~x3 | ~n1708) & ~n2010));
  assign n2010 = ~x5 & ((n1114 & n634) | (n628 & n633));
  assign n2011 = ~n2012 & n284 & n857;
  assign n2012 = (x1 | ~x6 | (~x2 ^ ~x7)) & (x2 | x6 | ~x7);
  assign z086 = n2014 | n2018 | ~n2023 | (~x1 & ~n2020);
  assign n2014 = ~x3 & (x5 ? (n559 & ~n2017) : ~n2015);
  assign n2015 = (x0 | n2016) & (~n1037 | (~x6 & ~x7));
  assign n2016 = (x1 | x6 | x7 | (x2 ^ ~x4)) & (~x1 | ~x2 | x4 | ~x6 | ~x7);
  assign n2017 = (~x6 | x7 | x1 | ~x2) & (~x1 | x2 | (x6 & x7));
  assign n2018 = n423 & ((n556 & n1483) | (x1 & ~n2019));
  assign n2019 = (x4 | ((~x0 | ~x5) & (~x6 | ~x7 | x0 | x5))) & (~x0 | ((~x5 | ~x6 | ~x7) & (x6 | x7 | ~x4 | x5)));
  assign n2020 = (~x4 | n2021) & (x0 | x4 | x5 | n2022);
  assign n2021 = (x6 | ~x7 | x3 | x5) & (~x3 | ((x5 | x6 | x7) & (~x6 | ~x7 | ~x0 | ~x5)));
  assign n2022 = x3 ? (~x6 | ~x7) : (x6 ^ ~x7);
  assign n2023 = (~x4 | n2027) & (n2024 | ~n2025) & (x4 | n2026);
  assign n2024 = (~x3 | ~x4 | x6 | x7) & (x3 | (x4 ? (x6 | ~x7) : (~x6 | x7)));
  assign n2025 = ~x5 & ~x0 & x1;
  assign n2026 = x3 ? (~x5 | (x0 & x1)) : (x5 | (~x0 & (~x1 | x6)));
  assign n2027 = (~x5 | ~x6 | x0 | ~x3) & (x3 | (x0 & x1) | (~x5 ^ x6));
  assign z087 = ~n2034 | (~n350 & ~n2032) | (~x3 & ~n2029);
  assign n2029 = ~n2030 & (~n329 | n331 | x7 | ~n587);
  assign n2030 = ~x4 & ((n441 & n313) | (x1 & ~n2031));
  assign n2031 = (x0 | x2 | x5 | ~x6 | ~x7) & (~x0 | ~x2 | x7 | (x5 ^ x6));
  assign n2032 = ~n2033 & (~n807 | ~n359) & (~n328 | n675);
  assign n2033 = (~x1 ^ ~x2) & ((~x5 & ~x6) | (x0 & x5 & x6));
  assign n2034 = ~n2040 & ~n2039 & n2037 & ~n2035 & ~n2036;
  assign n2035 = ~n315 & (x1 ? ~n534 : (x5 & ~n1254));
  assign n2036 = n425 & n579 & (x1 ? (x3 & x6) : (~x3 & ~x6));
  assign n2037 = x0 ? (~x2 | (x1 ? ~n1161 : ~n2038)) : (x2 | ~n2038);
  assign n2038 = ~x6 & ~x4 & x5;
  assign n2039 = n1964 & (~n1548 | (~x2 & x5 & n441));
  assign n2040 = n587 & n659 & (n841 | (n725 & n760));
  assign z088 = ~n2047 | (~x3 & ~n2043) | (~x1 & ~n2042);
  assign n2042 = (x0 | ((x5 | ~x7) & (~x2 | ~x5 | x7))) & (~x6 | x7 | ((~x0 | ~x2 | x5) & (x2 | ~x5)));
  assign n2043 = (~n2045 | ~n1747) & (x6 | (~n2044 & (~n2046 | ~n1747)));
  assign n2044 = ~x7 & x4 & ~x2 & ~x0 & ~x1;
  assign n2045 = ~x4 & x6 & (x5 ^ ~x7);
  assign n2046 = ~x4 & (~x5 ^ ~x7);
  assign n2047 = n2050 & (~x1 | n2048) & (~n579 | n2049);
  assign n2048 = (~x0 | x2 | x5 | ~x6 | x7) & (x0 | ((~x5 | ~x6 | x7) & (x2 | (x5 ? x7 : (x6 | ~x7)))));
  assign n2049 = (x1 | ~x3 | ~x5 | x6 | x7) & (~x1 | ~x6 | ~x7 | (x3 ^ x5));
  assign n2050 = (n2051 | n2052) & (~n423 | ~n387 | ~n430);
  assign n2051 = x5 ? (x6 ^ x7) : (x6 | ~x7);
  assign n2052 = x0 ^ (~x1 | ~x2);
  assign z089 = ~n2056 | ~n2057 | ~n2058 | (n579 & ~n2054);
  assign n2054 = (x4 | n2055) & (x1 | x3 | ~x4 | ~n876);
  assign n2055 = (x1 | x3 | ~x5 | x6 | x7) & (~x1 | ~x3 | ~x7 | (x5 ^ ~x6));
  assign n2056 = (~x0 | x6 | (x1 ^ ~x2)) & ~n1420 & (x0 | x1 | ~x2 | ~x6);
  assign n2057 = ~x6 | ~n579 | (n607 & (x4 | n369));
  assign n2058 = (n565 | n2060) & (x3 | n2059);
  assign n2059 = (~x0 | ~x1 | ~x2 | x4 | x6) & (x0 | x1 | x2 | ~x4 | ~x6);
  assign n2060 = x0 ? (x1 | x2) : (~x1 | (~x2 & (~x3 | ~x4)));
  assign z090 = n2062 | n2065 | ~n2066 | (n579 & ~n2064);
  assign n2062 = n408 & ((n280 & n654) | (x4 & ~n2063));
  assign n2063 = (~x0 | ~x3 | ~x5 | ~x6 | ~x7) & (x0 | x3 | x5 | (x6 ^ x7));
  assign n2064 = (x1 | x3 | ~x4 | ~x5 | ~x7) & (x4 | ((~x1 | ~x3 | (~x5 ^ x7)) & (x1 | x3 | ~x5 | x7)));
  assign n2065 = x1 & ((n324 & n2006) | (n579 & n404));
  assign n2066 = (x2 | ((~x0 | (~x1 ^ ~x7)) & (~x1 | x3 | ~x7))) & (x1 | ~x2 | ~x7) & (x0 | (x1 ? (~x2 | x7) : (~x3 | ~x7)));
  assign z091 = n2068 | ~n2071 | n2079 | (~x2 & ~n2078);
  assign n2068 = x4 & (n2069 | (n300 & n717 & n314));
  assign n2069 = n744 & ((n282 & n1973) | (n408 & n2070));
  assign n2070 = x6 & x3 & x5;
  assign n2071 = n2075 & ~n2074 & ~n2073 & ~n2072 & ~n1284;
  assign n2072 = n514 & n612;
  assign n2073 = x0 & ((x3 & ~x4 & ~x1 & ~x2) | (x1 & ~x3 & (x2 ^ x4)));
  assign n2074 = ~x2 & (x0 ? (x1 ^ ~x3) : (x1 & ~x3));
  assign n2075 = (~n359 | ~n2077) & (~n270 | ~n2076);
  assign n2076 = ~x3 & ~x2 & ~x0 & ~x1;
  assign n2077 = x6 & ~x5 & ~x3 & ~x4;
  assign n2078 = x0 ? ((~x1 | x3 | x4 | ~x5) & (x1 | ~x3 | ~x4 | x5)) : (x4 | (x1 ? (~x3 | x5) : (x3 | ~x5)));
  assign n2079 = x4 & (n2080 | (x3 & n1039 & n428));
  assign n2080 = n924 & (x3 ? (x6 & n282) : (~x6 & n408));
  assign z092 = ~n2086 | (~x1 & (~n2082 | n2083 | n2084));
  assign n2082 = x2 ? ((x0 | x3 | ~x4 | x5) & (x4 | ~x5 | ~x0 | ~x3)) : ((x0 | x3 | x4 | ~x5) & (~x4 | (x0 ? (~x3 ^ x5) : (~x3 | ~x5))));
  assign n2083 = n857 & ~n936;
  assign n2084 = n285 & ((n278 & n1039) | (~x2 & n2085));
  assign n2085 = ~x5 & (~x4 ^ ~x6);
  assign n2086 = ~n2093 & ~n2092 & n2089 & ~n2087 & ~n2088;
  assign n2087 = ~x0 & ((~x3 & ~x4 & ~x1 & x2) | (x1 & ((~x3 & x4) | (x2 & x3 & ~x4))));
  assign n2088 = x0 & (x1 ? (x2 ? (~x3 & ~x4) : (x3 & x4)) : (x3 & (~x2 ^ x4)));
  assign n2089 = (~n2025 | n2091) & (x4 | ~n725 | n2090);
  assign n2090 = x0 ? (x3 | x5) : (x3 ^ ~x5);
  assign n2091 = (~x2 | ~x3 | ~x4 | x6) & (x2 | x3 | x4 | ~x6);
  assign n2092 = ~n1028 & n327 & ~n751;
  assign n2093 = ~n2094 & ~x6 & n465;
  assign n2094 = (x0 | x1 | x2 | x4 | ~x7) & (~x0 | ~x1 | ~x2 | ~x4 | x7);
  assign z093 = ~n2098 | (~x2 & (x0 ? ~n2096 : ~n2097));
  assign n2096 = (~x1 | x3 | ~x4 | ~x5 | ~x6) & ((x1 ^ ~x4) | (x5 & (~x3 | x6)));
  assign n2097 = (x5 | (~x3 & x6) | (x1 ^ ~x4)) & (x1 | x4 | (~x5 & (x3 | ~x6)));
  assign n2098 = ~n2099 & ~n2105 & ~n2108 & (x3 | n2101);
  assign n2099 = n519 & ((n359 & n1183) | (x0 & ~n2100));
  assign n2100 = (~x1 | x2 | x4 | ~x5 | x7) & (x1 | ~x4 | (x2 ? (x5 | ~x7) : (~x5 | x7)));
  assign n2101 = (x5 | n2102) & (~x5 | ~x6 | ~n782 | ~n1065);
  assign n2102 = (~x0 | n2104) & (x0 | x2 | ~x7 | n2103);
  assign n2103 = x1 ? (~x4 | ~x6) : (x4 | x6);
  assign n2104 = (~x1 | ~x2 | ~x4 | x6 | x7) & (x1 | x2 | x4 | ~x6 | ~x7);
  assign n2105 = ~n1034 & (n2106 | (x3 & ~n2107));
  assign n2106 = x5 & ~x2 & ~x3;
  assign n2107 = x2 ? (x5 | x6) : (~x5 | ~x6);
  assign n2108 = x2 & (~n2110 | (x5 & n285 & ~n2109));
  assign n2109 = x1 ? (x4 | x6) : (x4 ^ ~x6);
  assign n2110 = (x0 & x3 & (~x4 | ~x5)) | (~x1 & ~x4) | (x1 & x4) | (~x0 & ~x3 & x5);
  assign z094 = n2112 | ~n2118 | (x2 ? ~n2116 : ~n2117);
  assign n2112 = x0 & ((~x7 & ~n2113) | (n270 & n272));
  assign n2113 = ~n2115 & (~x1 | ((~n426 | ~n764) & ~n2114));
  assign n2114 = x6 & x5 & ~x4 & ~x2 & x3;
  assign n2115 = n1752 & ((n425 & n340) | (~x2 & ~n1193));
  assign n2116 = (x0 | ~x5 | (x3 ^ x6)) & (x1 | ((x0 | x3 | x5 | ~x6) & (~x0 | (x3 ? (x5 | x6) : (~x5 | ~x6)))));
  assign n2117 = x5 ? ((x0 | x1 | x3 | ~x6) & (~x0 | ~x3 | x6)) : (((x0 ^ ~x1) | (x3 ^ x6)) & (x0 | x1 | ~x3 | x6) & (~x0 | ~x1 | x3 | ~x6));
  assign n2118 = n2119 & (n506 | n2124) & (~n709 | n2125);
  assign n2119 = ~n2121 & ~n2122 & (x4 | ~n441 | n2120);
  assign n2120 = (~x2 | x3 | x5 | x6 | ~x7) & (x2 | ((x3 | ~x5 | x6 | ~x7) & (~x3 | x5 | ~x6 | x7)));
  assign n2121 = n336 & ((x2 & (x1 ? (x4 & ~x5) : (~x4 & x5))) | (x1 & ~x2 & (~x4 ^ x5)));
  assign n2122 = ~n2123 & ((n308 & n1064) | (~x0 & ~n1502));
  assign n2123 = (x1 | ~x2 | ~x4 | ~x5) & (~x1 | (x2 ? (x4 | ~x5) : (~x4 | x5)));
  assign n2124 = (x0 | x1 | x2 | ~x4 | x5) & (~x0 | ((x1 | ~x2 | x4 | ~x5) & (~x1 | x2 | (x4 ^ x5))));
  assign n2125 = x0 ? ((~x1 | ~x2 | x4 | ~x5) & (~x4 | x5 | x1 | x2)) : (~x1 | (x2 ? (x4 ^ x5) : (x4 | ~x5)));
  assign z095 = n2127 | n2134 | n2141 | (~n602 & ~n2145);
  assign n2127 = x1 & (~n2130 | (~x0 & ~n2128));
  assign n2128 = x4 ? n2129 : (x2 | (~n882 & ~n1704));
  assign n2129 = x2 ? ((~x6 | ~x7 | x3 | x5) & (~x3 | ~x5 | x6 | x7)) : ((~x5 | x6 | ~x7) & (~x6 | x7 | x3 | x5));
  assign n2130 = ~n2133 & (~n413 | ~n2131) & (~n647 | n2132);
  assign n2131 = x7 & x4 & ~x6;
  assign n2132 = (~x3 | ~x4 | x5 | ~x6 | ~x7) & (x3 | ((~x4 | ~x5 | x6 | ~x7) & (x4 | x5 | ~x6)));
  assign n2133 = ~n645 & ((n624 & n717) | (n1207 & n382));
  assign n2134 = ~x1 & (n2135 | (x5 & (n2138 | ~n2139)));
  assign n2135 = ~x5 & ((n1683 & ~n2137) | (x4 & ~n2136));
  assign n2136 = (x0 | x2 | x3 | x6 | ~x7) & (~x0 | ~x2 | ~x3 | ~x6 | x7);
  assign n2137 = x0 ? ((~x2 & ~x3 & x7) | (x3 & (x2 | ~x7))) : ((~x3 & ~x7) | (~x2 & x3 & x7));
  assign n2138 = n700 & (x0 ? ((x3 & x7) | (x2 & ~x3 & ~x7)) : (~x3 & (x2 ^ ~x7)));
  assign n2139 = (x4 | n2140) & (n384 | (x0 ? (x4 | x6) : (x4 ^ ~x6)));
  assign n2140 = (~x0 | ~x2 | x3 | ~x6 | x7) & (x0 | x2 | ~x3 | x6 | ~x7);
  assign n2141 = ~n614 & (n2143 | n2144 | (~x6 & ~n2142));
  assign n2142 = (~x0 | x1 | ~x2 | ~x3 | ~x7) & (x0 | x2 | x3 | (~x1 ^ ~x7));
  assign n2143 = ~n1028 & ((x1 & x6 & ~x7) | (~x6 & (~x1 | x7)));
  assign n2144 = ~n645 & ((x1 & x2 & ~x6 & ~x7) | (x6 & ((~x2 & x7) | (~x1 & (~x2 | x7)))));
  assign n2145 = (~x1 | (x0 ? (x2 | ~x3) : x3)) & (x3 | x7 | x0 | ~x2) & (x1 | ((~x3 | ~x7 | (x0 & ~x2)) & (~x0 | (~x3 ^ x7))));
  assign z096 = n2147 | ~n2151 | n2159 | (~x0 & ~n2156);
  assign n2147 = x1 & ((n344 & n1145) | n2148 | n2150);
  assign n2148 = x4 & ((n313 & n713) | (n285 & ~n2149));
  assign n2149 = (~x2 | x5 | ~x6 | ~x7) & (x2 | ~x5 | (x6 ^ x7));
  assign n2150 = ~n1091 & ~n645 & (n634 | n1179);
  assign n2151 = ~n2153 & n2154 & (n1016 | n2152);
  assign n2152 = (x2 | x5 | ~x7) & (~x5 | x7 | ((~x0 | x2 | ~x3) & (~x2 | (x0 & x3))));
  assign n2153 = n340 & ((n387 & n341) | (x0 & n841));
  assign n2154 = (~n428 | ~n842) & (n570 | n2155);
  assign n2155 = x2 ? (x3 | ((x1 | x4) & (x0 | ~x1 | ~x4))) : ((~x1 | ~x3 | ~x4) & (~x0 | (x1 ? ~x4 : (~x3 | x4))));
  assign n2156 = (x3 | n2157) & (x1 | ~x3 | x4 | n2158);
  assign n2157 = (x1 | x2 | x4 | ~x5 | x7) & (~x1 | x5 | (x2 ? (x4 | ~x7) : (~x4 | x7)));
  assign n2158 = x2 ? (~x5 | ~x7) : (x5 | x7);
  assign n2159 = ~x1 & (n2160 | (~x6 & ~n1091 & ~n1024));
  assign n2160 = x6 & (~n2161 | (~n688 & ~n1091 & ~n645));
  assign n2161 = (x0 | x2 | x3 | ~n662) & (~x0 | ~x2 | ~x3 | ~n1187);
  assign z097 = n2163 | n2166 | ~n2171 | (n725 & ~n2169);
  assign n2163 = ~n1163 & ((~x0 & ~n2164) | (n330 & ~n2165));
  assign n2164 = (x7 | ((x1 | ~x2 | ~x4 | ~x5) & (~x1 | (x2 ? (x4 | ~x5) : (~x4 | x5))))) & (~x4 | ~x7 | ((~x2 | x5) & (x1 | x2 | ~x5)));
  assign n2165 = (x2 | x5 | x7) & (x1 | (x2 ? (x5 ^ ~x7) : (~x5 | ~x7)));
  assign n2166 = ~x2 & (x5 ? (n910 & ~n2168) : ~n2167);
  assign n2167 = (x0 | x1 | x3 | x4 | ~x6) & (x6 | ((x0 | ~x3 | (~x1 ^ x4)) & (x3 | ((~x1 | ~x4) & (~x0 | x1 | x4)))));
  assign n2168 = (~x0 | ~x3 | x6) & (x3 | ~x6);
  assign n2169 = (~x0 | x5 | ~n717 | ~n588) & (~x5 | n2170);
  assign n2170 = (x0 | x3 | x4 | ~x6 | ~x7) & (~x4 | ((x0 | ~x3 | x6 | ~x7) & (~x0 | (x3 ? (~x6 | x7) : (x6 | ~x7)))));
  assign n2171 = ~n2175 & ~n2176 & n2178 & (x1 | n2172);
  assign n2172 = (~x2 | n2173) & (x0 | x2 | x4 | n2174);
  assign n2173 = (x0 | x3 | x4 | ~n876) & (~x0 | ~x3 | ~x4 | ~n875);
  assign n2174 = (~x3 | x5 | ~x6 | x7) & (x3 | x6 | (~x5 ^ x7));
  assign n2175 = ~n1848 & (~x0 ^ (~x1 & ~x4));
  assign n2176 = ~n2177 & (x2 ? (~x5 ^ ~x6) : (~x5 ^ x6));
  assign n2177 = (x0 | x1 | ~x3 | x4) & (~x0 | x3 | (~x1 ^ x4));
  assign n2178 = (~x1 | x2 | x4 | n2179) & (x1 | (x2 ? n2180 : (~x4 | n2179)));
  assign n2179 = x0 ? (~x3 | ~x5) : (x3 | x5);
  assign n2180 = (~x0 | ~x3 | ~x4 | x5) & (x0 | x3 | x4 | ~x5);
  assign z098 = n2193 | ~n2196 | (x0 ? ~n2182 : ~n2187);
  assign n2182 = ~n2184 & (~n1295 | n2183) & (x5 | n2185);
  assign n2183 = (~x2 | ((~x3 | x4 | x6 | ~x7) & (x3 | ~x4 | ~x6 | x7))) & (x3 | x4 | ((~x6 | ~x7) & (x2 | x6 | x7)));
  assign n2184 = ~n271 & ((n606 & n921) | (~n542 & ~n1193));
  assign n2185 = (~x1 | n2186) & (x1 | x2 | x3 | n485);
  assign n2186 = (x2 | ~x3 | ~x4 | ~x6 | ~x7) & (~x2 | x3 | x4 | x6 | x7);
  assign n2187 = x4 ? (~n2192 & (x2 | n2191)) : n2188;
  assign n2188 = n2189 & ~n2190 & (n542 | n1116);
  assign n2189 = (x1 | x2 | x3 | ~n656) & (~x1 | ~x2 | ~x3 | ~n280);
  assign n2190 = ~n310 & ((n725 & n327) | (n438 & n328));
  assign n2191 = x6 ? ((~x1 | x3 | x5 | ~x7) & (x1 | (x3 ? (x5 | x7) : (~x5 | ~x7)))) : ((x3 | ~x5 | x7) & (~x1 | (x3 ? (~x5 | ~x7) : x7)));
  assign n2192 = n426 & ((n717 & n346) | (~n542 & ~n1417));
  assign n2193 = ~n565 & ((~x2 & ~n2194) | (n340 & ~n2195));
  assign n2194 = x4 ? ((~x0 | ~x1 | x3 | ~x5) & (x0 | ~x3 | (~x1 ^ x5))) : ((x0 | x1 | x3 | x5) & (~x0 | ~x3 | (x1 & x5)));
  assign n2195 = (x0 | ((~x4 | x5) & (~x1 | x4 | ~x5))) & (x1 | (x0 ? (x4 | x5) : ~x4));
  assign n2196 = n2199 & (x0 | (x4 & n2198) | (~x4 & n2197));
  assign n2197 = (~x3 | ~x6 | (x1 ^ (~x2 & ~x5))) & (~x1 | x3 | x6 | (x2 & x5));
  assign n2198 = (x1 | x2 | x3 | x5 | x6) & (~x1 | ~x5 | ((x3 | ~x6) & (~x2 | ~x3 | x6)));
  assign n2199 = (n614 | n2200) & (~x0 | (~n2201 & n2202));
  assign n2200 = (x0 | x1 | ~x2 | x3 | x6) & (~x0 | ~x1 | x2 | (~x3 ^ x6));
  assign n2201 = n346 & ((x2 & x4 & (x3 ^ x6)) | (~x2 & ~x3 & ~x4 & ~x6));
  assign n2202 = (~x1 | ~x2 | x3 | x4 | ~x6) & (x1 | x2 | ~x4 | (~x3 ^ x6));
  assign z099 = n2216 | ~n2218 | (x0 ? ~n2204 : ~n2210);
  assign n2204 = ~n2205 & (n1254 | n2208) & (~n923 | n2209);
  assign n2205 = ~x3 & ((~x7 & ~n2206) | (n789 & ~n2207));
  assign n2206 = (~x1 | x2 | x4 | ~x5 | ~x6) & (~x2 | ((~x5 | x6 | x1 | ~x4) & (~x1 | x5 | (~x4 ^ x6))));
  assign n2207 = (~x1 | ~x2 | x4 | x6) & (x1 | x2 | (x4 ^ ~x6));
  assign n2208 = (~x1 | x2 | ~x3 | x5 | ~x7) & (x1 | x3 | (x2 ? (~x5 | ~x7) : (x5 | x7)));
  assign n2209 = (x2 | x4 | x5 | x6 | x7) & (~x2 | ~x5 | (x4 ? (x6 | x7) : (~x6 ^ x7)));
  assign n2210 = ~n2211 & ~n2214 & ~n2215 & (n1263 | n2213);
  assign n2211 = n760 & ((n408 & n807) | (~n2212 & n1168));
  assign n2212 = x2 ? (~x3 | x5) : (x3 | ~x5);
  assign n2213 = (~x6 | x7) & (x3 | x6 | ~x7);
  assign n2214 = ~n542 & ((n725 & n547) | (n438 & n1265));
  assign n2215 = ~n1861 & (x1 ? (x2 & ~x6) : (~x2 & x6));
  assign n2216 = ~n688 & ~n2217;
  assign n2217 = x0 ? ((x1 | x5 | (~x2 & ~x3)) & (x2 | (x1 ? (x3 | x5) : ~x5))) : ((~x1 | ~x2 | ~x5) & (x3 | x5 | x1 | x2));
  assign n2218 = ~n2221 & ~n2223 & n2224 & (x2 | n2219);
  assign n2219 = (~n765 | ~n1187) & (~n2220 | n614 | n1556);
  assign n2220 = x3 & ~x7;
  assign n2221 = ~n2222 & (x0 ? (x2 & x5) : (~x2 ^ ~x5));
  assign n2222 = (x1 | ~x3 | ~x4 | ~x7) & (~x1 | x3 | x4 | x7);
  assign n2223 = ~n1024 & n387 & n501;
  assign n2224 = (~n364 | ~n1187) & (x0 | n350 | n1119);
  assign z100 = ~n2226 | n2230 | ~n2232 | (~n405 & ~n2231);
  assign n2226 = ~n2229 & (~x5 | n2227) & (~n709 | n2228);
  assign n2227 = ((~x3 ^ x6) | (x0 ? (~x1 | x2) : (x1 ^ x2))) & (~x3 | ~x6 | (x0 ? (x1 | ~x2) : (~x1 | x2)));
  assign n2228 = (x0 | ~x1 | x2 | ~x4 | ~x5) & (~x0 | ~x2 | (x1 ? (x4 | x5) : (~x4 | ~x5)));
  assign n2229 = n1241 & ((n656 & n606) | (x3 & n851));
  assign n2230 = ~x5 & ((~x1 & (x0 ? (x2 ^ x6) : (x2 & x6))) | (~x0 & x1 & ~x2 & ~x6));
  assign n2231 = (~x3 | ~x4 | ~x5 | x6 | ~x7) & (x3 | ~x6 | ((x5 | x7) & (x4 | ~x5 | ~x7)));
  assign n2232 = ~n2235 & (x6 | (~n2233 & (~n314 | n2234)));
  assign n2233 = ~n315 & ((n284 & n625) | (~x1 & ~n989));
  assign n2234 = (~x0 | ~x1 | ~x2 | x4) & (x0 | x1 | x2 | ~x4);
  assign n2235 = ~n315 & (x4 ? ~n2236 : ~n2237);
  assign n2236 = (~x1 | ~x3 | x5 | ~x6 | ~x7) & (x1 | x3 | ~x5 | x6 | x7);
  assign n2237 = (~x3 | (~x5 ^ x7) | (~x1 ^ ~x6)) & (~x1 | x3 | x6 | (x5 ^ x7));
  assign z101 = ~n2250 | ~n2248 | ~n2244 | n2239 | n2242;
  assign n2239 = ~n565 & (x0 ? ~n2241 : ~n2240);
  assign n2240 = x1 ? ((~x4 | ~x5 | x2 | ~x3) & (x4 | x5 | ~x2 | x3)) : (x2 ? (x3 ? (x4 | x5) : (~x4 | ~x5)) : (x3 | x4));
  assign n2241 = (~x1 | x2 | x3 | x4 | x5) & (x1 | ((~x2 | ~x3 | ~x4 | ~x5) & (x2 | (x3 ? (x4 | x5) : (~x4 | ~x5)))));
  assign n2242 = ~n542 & ((~n614 & ~n2243) | (n359 & n612));
  assign n2243 = x0 ? (x1 ? (x2 | ~x3) : (~x2 | x3)) : (x1 ? (x2 ^ x3) : (x2 | ~x3));
  assign n2244 = n2247 & (n602 | n2246) & (n598 | n2245);
  assign n2245 = x0 ? (x1 ^ ~x3) : (x1 | x3);
  assign n2246 = x0 ? (x1 ? (x2 | ~x3) : (~x2 | x3)) : (~x1 | (x2 ^ x3));
  assign n2247 = ~n408 | (x0 ? ~n1761 : ~n757);
  assign n2248 = (x0 | n2249) & (n585 | n2246);
  assign n2249 = (x1 | ~x2 | ~x3 | ~x4 | x6) & (~x1 | ((x2 | ~x3 | x4 | ~x6) & (~x2 | x3 | ~x4 | x6)));
  assign n2250 = x0 ? (~n2254 & ~n2255) : (~n2251 & ~n2252);
  assign n2251 = x1 & ((n656 & n892) | (n280 & n1453));
  assign n2252 = ~x1 & (x2 ? ~n2253 : (n443 & n313));
  assign n2253 = (x3 | ~x4 | x5 | ~x6 | x7) & (~x3 | x4 | ~x5 | x6 | ~x7);
  assign n2254 = ~x1 & (x2 ? (n280 & n588) : ~n2253);
  assign n2255 = n1986 & n1145;
  assign z102 = ~n2259 | (x7 & ~n2257);
  assign n2257 = (x0 | n2258) & (n614 | n2243) & (~x0 | n2241);
  assign n2258 = x1 ? ((~x4 | ~x5 | x2 | ~x3) & (x4 | x5 | ~x2 | x3)) : ((x4 | x5 | x2 | x3) & (~x2 | (x3 ? (x4 | x5) : (~x4 | ~x5))));
  assign n2259 = ~n2262 & ~n2264 & (x5 ? n2260 : n2268);
  assign n2260 = (n565 | n2261) & (~x3 | ~n408 | n1945);
  assign n2261 = (x0 | ~x2 | ~x3 | (~x1 ^ ~x4)) & (x3 | ((~x0 | (x1 ? (x2 | x4) : (~x2 | ~x4))) & (x0 | ~x1 | ~x2 | x4)));
  assign n2262 = ~n1274 & (x7 ? ~n2263 : (n725 & ~n602));
  assign n2263 = (x1 | ~x2 | ~x4 | x5 | ~x6) & (x2 | ((x1 | x4 | ~x5 | x6) & (~x1 | (x4 ? (~x5 | x6) : (x5 | ~x6)))));
  assign n2264 = ~x7 & (n2265 | ~n2266 | (~n736 & ~n2245));
  assign n2265 = ~x0 & ((x3 & x4 & ~x1 & x2) | (x1 & (x2 ? (~x3 & x4) : (x3 & ~x4))));
  assign n2266 = x1 | (x0 ? ~n974 : (x5 | n2267));
  assign n2267 = x2 ? (x3 | ~x4) : (~x3 | x4);
  assign n2268 = ~n2269 & ~n2270 & (~n443 | ~n717 | ~n359);
  assign n2269 = ~n607 & n700 & ~x7 & n324;
  assign n2270 = ~n736 & ~n542 & (n1177 | (x0 & n276));
  assign z103 = ~n2274 | (n441 & (x3 ? ~n2273 : ~n2272));
  assign n2272 = x2 ? ((x6 | x7 | x4 | ~x5) & (~x6 | ~x7 | ~x4 | x5)) : (~x5 | (x4 ? (x6 | x7) : (~x6 | ~x7)));
  assign n2273 = (~x2 | x4 | x5 | x6 | x7) & (x2 | ((~x6 | ~x7 | x4 | x5) & (~x4 | (x5 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n2274 = ~n2275 & n2276 & ~n2279 & (n677 | n2280);
  assign n2275 = n624 & (x0 ? (x1 & n465) : (~x1 & n2070));
  assign n2276 = (x0 | (n2277 & (~x1 | ~x6 | n2278))) & (~x6 | n2277) & (~x0 | x1 | n2278);
  assign n2277 = (~x1 | x2 | x3 | x4 | ~x5) & (x1 | ~x2 | ~x3 | ~x4 | x5);
  assign n2278 = (~x4 | x5 | x2 | ~x3) & (~x2 | x3 | x4 | ~x5);
  assign n2279 = ~n668 & (x0 ? (x1 ? ~x2 : n740) : (~x1 ^ x2));
  assign n2280 = x1 ? ((x2 | ~x3 | ~x6) & (x0 | ((~x3 | ~x6) & (x2 | (~x3 & ~x6))))) : ((~x0 | (x2 ^ x3)) & (~x2 | x3 | (x0 & ~x6)));
  assign z104 = n2282 | ~n2287 | ~n2293 | (~n534 & ~n2286);
  assign n2282 = ~n379 & (~n2283 | n2285 | (~x1 & ~n2284));
  assign n2283 = x0 ? ((x1 | ~x2 | x3 | ~x4) & (x2 | (x1 ? (x3 ^ x4) : (~x3 | x4)))) : (x2 ? ((x3 | x4) & (~x1 | ~x3 | ~x4)) : (x3 | ~x4));
  assign n2284 = (x0 | ~x2 | ~x3 | ~x4 | x7) & ((x0 ^ ~x7) | (x2 ? (~x3 | x4) : (x3 ^ x4)));
  assign n2285 = n1369 & ((~x0 & ~x2 & x3 & ~x4) | (~x3 & (x0 ? (x2 ^ x4) : (x2 & x4))));
  assign n2286 = (x1 | ((~x2 | (x0 ? ~x3 : (x3 | ~x7))) & (~x0 | x3 | (x2 & x7)))) & (~x1 | x2 | ~x3 | x7) & (x0 | ((x2 | ~x3) & (~x1 | x7 | (x2 & ~x3))));
  assign n2287 = ~n2291 & (~x1 | (~n2288 & ~n2290));
  assign n2288 = ~n315 & (n2289 | (n587 & n443));
  assign n2289 = ~x6 & x5 & ~x3 & x4;
  assign n2290 = n606 & ((n587 & n579) | (n324 & n1039));
  assign n2291 = n1369 & (x0 ? (n339 & n273) : ~n2292);
  assign n2292 = (~x2 | x3 | x4 | x5 | ~x6) & (x2 | ~x3 | ~x4 | ~x5 | x6);
  assign n2293 = x1 | (n2294 & ~n2298 & (~x3 | n2296));
  assign n2294 = x0 ? n2292 : n2295;
  assign n2295 = (x2 | x3 | x4 | x5 | ~x6) & (~x2 | ((~x4 | ~x5 | x6) & (~x3 | x4 | x5 | ~x6)));
  assign n2296 = (x7 | n2297) & (x0 | ~n366 | ~n313);
  assign n2297 = (x0 | ~x2 | x4 | ~x5 | ~x6) & (~x0 | ((x5 | ~x6 | x2 | x4) & (~x2 | ~x4 | ~x5 | x6)));
  assign n2298 = ~n2299 & n284 & ~x6 & n339;
  assign n2299 = x0 ^ ~x7;
  assign z105 = n2302 | n2307 | ~n2309 | (~n555 & ~n2301);
  assign n2301 = x1 ? ((x2 | ~x3 | x4) & (x0 | ((~x2 | x3 | ~x4) & (~x3 | x4) & (x2 | (~x3 & x4))))) : ((~x2 | (x3 ^ x4)) & (x3 | (x4 ? x2 : ~x0)));
  assign n2302 = ~n542 & (~n2303 | n2305 | (x4 & ~n2306));
  assign n2303 = n2304 & (n668 | (~n438 & (x0 | ~n725)));
  assign n2304 = (x1 | x2 | x3 | x4 | ~x5) & (~x1 | ((~x2 | x3 | x4 | ~x5) & (x2 | ~x3 | ~x4 | x5)));
  assign n2305 = ~n677 & (n514 | (~x2 & ~n607));
  assign n2306 = (~x0 | x1 | x2 | x3 | x5) & (x0 | ~x2 | ~x3 | (~x1 ^ x5));
  assign n2307 = ~n2308 & (n514 | (~x2 & ~n703));
  assign n2308 = (~x3 | ~x5 | ~x6 | x7) & (x3 | x5 | x6 | ~x7);
  assign n2309 = x3 ? n2312 : n2310;
  assign n2310 = (~n270 | ~n742) & (x7 | ~n327 | n2311);
  assign n2311 = (x0 & (x4 ? x1 : x2)) | (x1 & x2 & x4) | (~x1 & (~x4 | (~x0 & ~x2)));
  assign n2312 = (~n300 | ~n714) & (~x7 | ~n328 | n2313);
  assign n2313 = (x1 | (x2 ^ ~x4)) & (x0 | ((~x2 | ~x4) & (~x1 | x2 | x4)));
  assign z106 = ~n2324 | n2323 | n2315 | n2318;
  assign n2315 = ~x5 & ((n579 & n345) | n2316);
  assign n2316 = x0 & ((~x6 & ~n2317) | (n1658 & n622));
  assign n2317 = (x4 | ~x7 | x1 | ~x3) & (x3 | ((~x1 | ~x2 | ~x4 | x7) & (x2 | x4 | ~x7)));
  assign n2318 = ~n542 & (n2320 | ~n2321 | (x5 & ~n2319));
  assign n2319 = (x0 | ((~x3 | ~x4 | x1 | ~x2) & (x2 | x3 | x4))) & (x4 | ((~x0 | x1 | ~x2 | ~x3) & (~x1 | x2 | x3)));
  assign n2320 = ~n283 & (x0 ? ~x1 : x3);
  assign n2321 = (n677 | n2322) & (~n579 | ~n1265);
  assign n2322 = x3 ? (x2 | (~x0 & ~x1)) : (~x2 | (x0 & x1));
  assign n2323 = n1476 & (x0 ? (~x1 & x2) : (~x2 ^ x3));
  assign n2324 = (n1517 | n2326) & (n555 | n2325);
  assign n2325 = (x0 & ((x1 & x3) | (~x2 & ~x4))) | (~x0 & ~x3 & (x2 | (~x1 & x4))) | (x2 & x4) | (~x2 & x3 & ~x4);
  assign n2326 = (x0 & (x3 ? x2 : x1)) | (x1 & x2 & x3) | (~x2 & (~x3 | (~x0 & ~x1)));
  assign z107 = ~n2336 | (x4 ? ~n2332 : ~n2328);
  assign n2328 = n2331 & (x1 ? n2329 : (n566 | n1502));
  assign n2329 = (~n556 | ~n661) & (x6 | n2330);
  assign n2330 = (~x0 | ~x2 | x3 | x5 | ~x7) & (~x3 | ((~x5 | ~x7 | x0 | ~x2) & (x2 | (x0 ? (x5 ^ x7) : (x5 | ~x7)))));
  assign n2331 = (~n394 | ~n882) & (~n280 | ~n728);
  assign n2332 = ~n2334 & (~n394 | ~n2333);
  assign n2333 = x7 & ~x6 & ~x3 & ~x5;
  assign n2334 = ~x0 & ((x3 & n656) | (~x7 & ~n2335));
  assign n2335 = (~x1 | ((x3 | ~x5 | ~x6) & (~x2 | ~x3 | x5 | x6))) & (x3 | ~x6 | ((x1 | x2 | x5) & (~x2 | ~x5)));
  assign n2336 = ~n2338 & (n731 | n2337) & (n565 | n2344);
  assign n2337 = x0 ? ((x4 | x5 | x1 | ~x2) & (x2 | (x1 ? (x4 ^ x5) : (~x4 | x5)))) : (x1 ? (~x4 | x5) : (x4 | ~x5));
  assign n2338 = ~n542 & (n2342 | ~n2343 | n2339 | n2341);
  assign n2339 = ~n331 & (x0 ? ~n2340 : ~n668);
  assign n2340 = x3 ? (~x4 | x5) : (x4 ^ x5);
  assign n2341 = n443 & ((~x0 & (x1 ? (x2 & x5) : (~x2 & ~x5))) | (x0 & ~x1 & ~x2 & x5));
  assign n2342 = ~x0 & ((x4 & x5 & ~x1 & x3) | (~x4 & ~x5 & x1 & ~x3));
  assign n2343 = ~x1 | (x0 ? ~n1458 : (~x2 | ~n356));
  assign n2344 = n2347 & (x2 | n2346) & (x0 | n2345);
  assign n2345 = (~x4 | x5 | x1 | ~x3) & (~x1 | x3 | x4 | ~x5);
  assign n2346 = (x0 | x1 | x3 | ~x4 | ~x5) & (~x0 | x5 | (x1 ? (x3 | ~x4) : (~x3 | x4)));
  assign n2347 = (~n514 | ~n1270) & (~n363 | ~n612);
  assign z108 = ~n2352 | (x1 & ((n661 & n1755) | n2349));
  assign n2349 = x4 & (x3 ? (n647 & n2350) : ~n2351);
  assign n2350 = ~x5 & (~x6 ^ x7);
  assign n2351 = (x6 | x7 | ~x2 | x5) & (x0 | x2 | ~x5 | (x6 ^ x7));
  assign n2352 = n2356 & ~n2361 & ~n2364 & (x1 | n2353);
  assign n2353 = (n605 | n2354) & (x7 | n388 | ~n2355);
  assign n2354 = (x0 | ~x3 | x4 | ~x6 | x7) & (~x0 | ~x7 | (x3 ? (~x4 | x6) : (x4 | ~x6)));
  assign n2355 = ~x6 & ~x5 & ~x0 & ~x4;
  assign n2356 = (n555 | n2357) & (x0 | (~n2358 & ~n2359));
  assign n2357 = ((x2 & x3) | ((~x1 | x4) & (~x0 | x1 | ~x4))) & (x3 | ~x4 | x1 | x2) & (x0 | ~x2 | (~x1 ^ ~x4));
  assign n2358 = x1 & ((n624 & n875) | (n1207 & n876));
  assign n2359 = n913 & (x2 ? ~n2360 : (x5 & n717));
  assign n2360 = x5 ? (~x6 | ~x7) : (x6 | x7);
  assign n2361 = ~n1291 & ((~x3 & ~n820) | n2362 | (x3 & ~n2363));
  assign n2362 = ~n836 & ((x0 & (~x1 ^ ~x2)) | (~x1 & (x2 ? ~x3 : ~x0)));
  assign n2363 = (~x0 | x1 | x2 | x4) & (x0 | (x1 ? (x4 ^ x6) : (~x2 | ~x4)));
  assign n2364 = x0 & (x1 ? (n1207 & n875) : ~n2365);
  assign n2365 = (~x2 | ~x4 | ~x5 | ~x6 | ~x7) & (x4 | ((x5 | x6 | x7) & (~x6 | ~x7 | x2 | ~x5)));
  assign z109 = n2377 | ~n2382 | (x2 ? ~n2367 : ~n2372);
  assign n2367 = ~n2368 & (~n367 | n2371);
  assign n2368 = x6 & ((~x1 & ~n2369) | (n387 & ~n2370));
  assign n2369 = (x4 | (x0 ? (x3 ? (x5 | x7) : (~x5 | ~x7)) : (~x5 | x7))) & (x0 | x3 | ((~x4 | x5 | ~x7) & (~x5 | x7)));
  assign n2370 = (~x3 | ((~x5 | x7) & (~x4 | x5 | ~x7))) & (x7 | ((~x4 | ~x5) & (x3 | x4 | x5)));
  assign n2371 = (x1 | x3 | ((x5 | ~x7) & (x4 | ~x5 | x7))) & (~x3 | ((x4 | x5 | ~x7) & (~x1 | ((x5 | ~x7) & (~x4 | ~x5 | x7)))));
  assign n2372 = x5 ? (~n2374 & (~x6 | n2373)) : n2375;
  assign n2373 = (x0 | ~x1 | ~x3 | x4 | ~x7) & (x7 | ((x0 | x1 | ~x3 | ~x4) & (~x0 | (~x1 & (x3 | x4)))));
  assign n2374 = ~x6 & n625 & (x0 ? n1074 : n760);
  assign n2375 = x0 ? (~x7 | n2376) : (~n620 | ~n635);
  assign n2376 = (~x1 & x3) | (x6 & (~x3 | x4));
  assign n2377 = ~n542 & (n2379 | ~n2380 | (x2 & ~n2378));
  assign n2378 = (x0 | ~x1 | ~x3 | x4 | x5) & (x3 | (x0 ? (x1 ? (x4 | ~x5) : (~x4 | x5)) : (x1 | (x4 ^ x5))));
  assign n2379 = ~x2 & ((~x0 & ~x1 & x3 & ~x5) | (x5 & (x0 ? (x1 ^ ~x3) : (x1 & ~x3))));
  assign n2380 = n2381 & (~x4 | x5 | ~n579 | n954);
  assign n2381 = (~x0 | x1 | ~x2 | ~x3 | x5) & ((x0 ^ ~x2) | (x1 ? (x3 | x5) : (~x3 | ~x5)));
  assign n2382 = (n555 | n2385) & (n565 | (~n2383 & ~n2384));
  assign n2383 = n923 & (x0 ? (x2 ? x5 : (~x4 & ~x5)) : (x2 ? (x4 & ~x5) : (~x4 & x5)));
  assign n2384 = ~x4 & n625 & (x0 ? (x2 & ~x5) : (x2 ^ ~x5));
  assign n2385 = (x1 | (x0 ? (x2 ? x3 : (~x3 | ~x4)) : (x2 | x3))) & (x0 | x2 | (x3 ? ~x1 : ~x4));
  assign z110 = ~n2387 | n2399 | n2402 | (~x3 & ~n2394);
  assign n2387 = n2390 & (x2 | (x0 & n2388) | (~x0 & n2389));
  assign n2388 = (x1 | x3 | ~x4 | ~x5 | x6) & (~x1 | ~x3 | x4 | x5 | ~x6);
  assign n2389 = (x1 | ~x3 | ~x4 | x5 | x6) & (x3 | ((x1 | x4 | x5 | ~x6) & (~x1 | (x4 ? (~x5 | ~x6) : (x5 | x6)))));
  assign n2390 = ~n2393 & (~n782 | n2391) & (~x3 | n2392);
  assign n2391 = (x1 | ~x3 | ~x4 | ~x5 | x6) & (x3 | (x1 ^ ~x6) | (x4 ^ ~x5));
  assign n2392 = (x0 | ~x1 | ~x6 | (x2 ^ x4)) & (x1 | x6 | ((x2 | x4) & (~x0 | ~x2 | ~x4)));
  assign n2393 = n1064 & ((n438 & n1683) | (x1 & ~n902));
  assign n2394 = n2397 & (n542 | n2396) & (n1974 | n2395);
  assign n2395 = (x1 | ~x2 | ~x4 | ~x6 | x7) & (~x1 | ((~x4 | x6 | x7) & (x2 | ((x6 | x7) & (x4 | ~x6 | ~x7)))));
  assign n2396 = (~x0 | ~x1 | x2 | x4 | ~x5) & (x0 | x5 | (x1 ? (x2 | ~x4) : (~x2 | x4)));
  assign n2397 = (~n514 | ~n1022) & (x4 | ~n363 | ~n2398);
  assign n2398 = ~x5 & ~x7 & (~x2 ^ ~x6);
  assign n2399 = ~n565 & (x1 ? ~n2401 : ~n2400);
  assign n2400 = (x0 | (x2 ? (~x3 | x4) : (x3 | ~x5))) & (x2 | x3 | (~x4 ^ x5)) & (~x2 | ((~x3 | x4 | x5) & (~x4 | ~x5 | ~x0 | x3)));
  assign n2401 = (x0 | ~x2 | x3 | x4 | x5) & (x2 | ~x3 | (~x4 & (~x0 | ~x5)));
  assign n2402 = x3 & ((~n542 & ~n2403) | (~x1 & n2404));
  assign n2403 = (~x2 | x4 | x0 | ~x1) & (x1 | x2 | ~x4 | (~x0 & ~x5));
  assign n2404 = x7 & ~n998 & (x0 ? n424 : n425);
  assign z111 = ~n2413 | (x3 ? (n2406 | n2408) : ~n2409);
  assign n2406 = x5 & (x0 ? ~n2407 : (n282 & n633));
  assign n2407 = (x1 | ~x2 | x4 | (x6 ^ x7)) & (x2 | ((x1 | x4 | x6 | ~x7) & (~x1 | ~x6 | (x4 ^ x7))));
  assign n2408 = n425 & n441 & (x2 ? (~x6 & ~x7) : (~x6 ^ ~x7));
  assign n2409 = ~n2410 & (~n730 | n2412);
  assign n2410 = ~x5 & (x0 ? ~n2411 : (n282 & n633));
  assign n2411 = (x1 | ~x2 | x6 | (x4 ^ x7)) & (x2 | (x1 ? (~x4 | (x6 ^ x7)) : (x4 | (~x6 ^ x7))));
  assign n2412 = x1 ? (~x4 | (x2 ? (~x6 | x7) : (x6 ^ x7))) : ((~x2 | ~x4 | x6 | ~x7) & (~x6 | x7 | x2 | x4));
  assign n2413 = ~n2414 & ~n2416 & n2419 & (x0 | n2418);
  assign n2414 = ~x7 & (x2 ? (n363 & ~n766) : ~n2415);
  assign n2415 = (x0 | x1 | ~x3 | ~x4 | ~x5) & (x3 | (~x4 ^ x5) | (x0 ^ ~x1));
  assign n2416 = x7 & ~n2417;
  assign n2417 = (x0 | ~x2 | x3 | (~x4 ^ x5)) & (x2 | ((x4 | x5 | x0 | x3) & (~x0 | (x3 ? (x4 | x5) : (~x4 | ~x5)))));
  assign n2418 = (~x3 | x4 | (~x2 ^ x7)) & (x1 | ~x4 | (x2 ? (~x3 | ~x7) : (x3 | x7)));
  assign n2419 = ~n2420 & (x0 ? n2421 : (~n426 | ~n662));
  assign n2420 = ~n847 & ((n387 & n588) | (x0 & ~n357));
  assign n2421 = (~x1 | x2 | ~x3 | ~x4 | x7) & (x1 | ~x2 | x3 | x4 | ~x7);
  assign z112 = ~n2427 | ~n2437 | (x1 & (n2423 | n2425));
  assign n2423 = ~x6 & ((n659 & n1187) | (~x3 & ~n2424));
  assign n2424 = x0 ? ((~x5 | ~x7 | x2 | x4) & (~x2 | ~x4 | x5 | x7)) : (~x4 | (x2 ? (~x5 | x7) : (x5 | ~x7)));
  assign n2425 = ~n2426 & x6 & n601;
  assign n2426 = (x5 | ~x7 | x2 | ~x3) & (~x2 | x7 | (x3 ^ x5));
  assign n2427 = ~n2428 & ~n2433 & ~n2435 & (~n387 | n2436);
  assign n2428 = ~x1 & (~n2430 | (x6 & n857 & ~n2429));
  assign n2429 = (x2 | x4 | ~x5 | x7) & (~x2 | ~x4 | x5 | ~x7);
  assign n2430 = (~n344 | ~n595) & (n2432 | (~n807 & ~n2431));
  assign n2431 = x6 & ~x3 & x5;
  assign n2432 = (~x4 | x7 | x0 | ~x2) & (~x0 | x2 | x4 | ~x7);
  assign n2433 = ~n1254 & ((n1241 & n1876) | (n744 & ~n2434));
  assign n2434 = (~x1 | x2 | ~x3 | ~x5) & (x1 | ~x2 | x3 | x5);
  assign n2435 = ~n673 & (n1471 | (~n271 & n1064));
  assign n2436 = (~x3 | ~x4 | ~x5 | ~x6) & (~x2 | x3 | x4 | x5 | x6);
  assign n2437 = n2438 & ~n2442 & (n377 | n2441);
  assign n2438 = x4 ? n2440 : n2439;
  assign n2439 = x1 ? (x0 ? (x2 ? (x3 | ~x5) : (~x3 | x5)) : (x2 | (x3 ^ x5))) : (~x2 | (x0 ? (~x3 | x5) : (x3 ^ x5)));
  assign n2440 = (x0 | ~x1 | ~x2 | x3 | x5) & (x1 | ((x0 | x2 | x3 | ~x5) & (~x0 | ((~x3 | ~x5) & (x2 | x3 | x5)))));
  assign n2441 = (x0 | ~x2 | (x1 ? (~x3 | x4) : (x3 | ~x4))) & (x2 | ((x0 | ~x1 | x3 | ~x4) & (~x0 | ~x3 | (~x1 ^ ~x4))));
  assign n2442 = ~x1 & ((~x4 & ~n2443) | (n301 & n413));
  assign n2443 = (x0 | x2 | x3 | x5 | ~x6) & (~x0 | x6 | (x2 ? (~x3 | ~x5) : (x3 | x5)));
  assign z113 = ~n2459 | ~n2455 | n2452 | n2445 | n2448;
  assign n2445 = ~x0 & ((n296 & n628) | n2446);
  assign n2446 = ~x5 & ((n345 & n628) | (x6 & ~n2447));
  assign n2447 = (x1 | ~x2 | ~x3 | x4 | x7) & (~x1 | x3 | ~x4 | (~x2 ^ x7));
  assign n2448 = x3 & (n2450 | n2451 | (x6 & ~n2449));
  assign n2449 = (x0 | ~x1 | x2 | x4 | x7) & (x1 | ((~x0 | ~x4 | (~x2 ^ x7)) & (x4 | ~x7 | x0 | ~x2)));
  assign n2450 = ~n1254 & (x2 ? (x7 & n387) : (~x7 & n363));
  assign n2451 = ~n409 & n438 & n700;
  assign n2452 = ~x3 & (x0 ? ~n2453 : ~n2454);
  assign n2453 = (~x7 | ((x1 | x2 | ~x4 | ~x6) & (~x1 | (x2 ? (x4 | ~x6) : (~x4 | x6))))) & (x1 | ((x4 | x6 | (x2 & x7)) & (~x2 | ~x4 | ~x6 | x7)));
  assign n2454 = (x1 | ~x2 | ~x4 | x6 | x7) & (~x1 | x2 | x4 | ~x6 | ~x7) & ((x1 ? (~x2 | x4) : (x2 | ~x4)) | (~x6 ^ x7));
  assign n2455 = (n614 | n2457) & (n836 | n2456);
  assign n2456 = (x0 | x1 | ~x2 | x3 | ~x7) & (x2 | ((~x0 | ~x1 | ~x3 | ~x7) & (x0 | (x1 ? (x3 | x7) : (~x3 | ~x7)))));
  assign n2457 = (x2 | x7 | n2458) & (n1402 | (x2 ? (x3 ^ ~x7) : (~x3 | ~x7)));
  assign n2458 = x0 ? (x1 ? x6 : (x3 | ~x6)) : (x1 | x6);
  assign n2459 = ~n2462 & (n677 | (~n2461 & (~x6 | n2460)));
  assign n2460 = (x2 | (~x0 ^ ~x1) | (~x3 ^ x7)) & (x1 | ~x2 | (x0 ? ~x7 : (x3 | x7)));
  assign n2461 = n367 & ((~x1 & x2 & x3 & x7) | (x1 & (x2 ? ~x7 : (~x3 & x7))));
  assign n2462 = x0 & (x4 ? (n625 & n2465) : ~n2463);
  assign n2463 = (~n280 | ~n1127) & (~x5 | ~n923 | n2464);
  assign n2464 = x2 ? (x6 | ~x7) : (~x6 | x7);
  assign n2465 = ~x7 & (x2 ? (~x5 & ~x6) : (x5 & x6));
  assign z114 = ~n2478 | ~n2475 | ~n2472 | n2467 | n2470;
  assign n2467 = ~n1291 & (~n2469 | (x6 & ~n2468));
  assign n2468 = (x4 | ((x0 | x1 | ~x2 | ~x3) & (~x0 | (x1 ? (~x2 | x3) : (x2 | ~x3))))) & (x0 | ~x3 | ~x4 | (x1 ^ x2));
  assign n2469 = ((x0 ^ ~x2) | (x1 ? x6 : (x3 | ~x6))) & (x2 | (x0 ? (~x1 | ~x3) : (x1 | x6)));
  assign n2470 = ~n542 & (x3 ? ~n2471 : (n335 & n295));
  assign n2471 = (x0 | ~x1 | x2 | ~x5) & (x1 | ((~x4 | x5 | x0 | ~x2) & (~x0 | (x2 ? ~x5 : (~x4 | x5)))));
  assign n2472 = (n2473 | n2474) & (~n295 | ~n443 | ~n450);
  assign n2473 = x2 ? (~x6 | x7) : (x6 | ~x7);
  assign n2474 = (x0 | ~x1 | ~x5 | (x3 ^ ~x4)) & (~x0 | x1 | x3 | x5);
  assign n2475 = ~n2477 & (x3 | ((~n295 | ~n1422) & ~n2476));
  assign n2476 = n786 & (n394 | (n366 & n387));
  assign n2477 = n625 & ((x2 & ~n960) | (x0 & ~x2 & n327));
  assign n2478 = ~n2482 & (x3 ? n2479 : (~n2485 & ~n2487));
  assign n2479 = (~n425 | ~n521 | ~n295) & (x1 | n2480);
  assign n2480 = (x7 | n2481) & (~x0 | ~n624 | ~n656);
  assign n2481 = (x0 | x2 | x4 | ~x5 | ~x6) & (x5 | (x0 ^ ~x2) | (x4 ^ x6));
  assign n2482 = ~x1 & (x0 ? ~n2483 : ~n2484);
  assign n2483 = (x6 | x7 | x3 | x5) & (~x3 | ((~x6 | x7 | ~x2 | x5) & (x6 | ~x7 | x2 | ~x5)));
  assign n2484 = (x2 | x3 | x5 | ~x6 | x7) & (~x7 | ((x2 | x3 | ~x5 | ~x6) & (~x2 | x6 | (x3 ^ x5))));
  assign n2485 = x1 & (n2486 | (~x0 & n1207 & n875));
  assign n2486 = n335 & (x0 ? ~n2464 : n521);
  assign n2487 = n913 & ((n656 & n647) | (~x0 & n2465));
  assign z115 = ~n2500 | ~n2509 | (x5 ? ~n2496 : ~n2489);
  assign n2489 = x0 ? (~n2491 & (x1 | n2490)) : n2493;
  assign n2490 = (~x2 | x3 | x4 | x6 | x7) & (~x3 | ~x4 | ((~x6 | ~x7) & (x2 | x6 | x7)));
  assign n2491 = n725 & (n2492 | (~x3 & n626));
  assign n2492 = ~x7 & ~x6 & x3 & ~x4;
  assign n2493 = x1 ? (x3 ? (x4 | n2495) : n2494) : (~x3 | n2494);
  assign n2494 = (x2 | x4 | (x6 ^ x7)) & (~x2 | ~x4 | ~x6 | ~x7);
  assign n2495 = (x6 | x7) & (~x2 | ~x6 | ~x7);
  assign n2496 = n2498 & (x2 | n2497);
  assign n2497 = (x0 | x1 | x3 | ~n626) & (~x0 | ~x1 | n638);
  assign n2498 = (n607 | n2499) & (~n300 | ~n717 | ~n356);
  assign n2499 = (x0 | x2 | x4 | x6 | x7) & (~x4 | (x0 ^ ~x2) | (x6 ^ x7));
  assign n2500 = n2505 & (n565 | (n2501 & ~n2502 & ~n2503));
  assign n2501 = x0 ? (x4 | (x1 ? (~x2 | x3) : (x2 ^ x3))) : ((x1 | ~x2 | x3 | ~x4) & (~x1 | x2 | ~x3 | x4));
  assign n2502 = ~x0 & ((n725 & n429) | (n438 & n1458));
  assign n2503 = n559 & ((n725 & n464) | (n346 & ~n2504));
  assign n2504 = ~x2 ^ ~x3;
  assign n2505 = n2508 & (x0 | n2507) & (n506 | n2506);
  assign n2506 = (~x0 | x1 | ~x2 | ~x4 | ~x5) & (x0 | ((x4 | x5 | x1 | ~x2) & (~x4 | ~x5 | ~x1 | x2)));
  assign n2507 = (x1 | x2 | ~x3 | ~x4 | x6) & (~x1 | ~x2 | x3 | x4 | ~x6);
  assign n2508 = (~n428 | ~n825) & (~n782 | ~n464 | n1087);
  assign n2509 = (n614 | n2510) & (~n339 | n2511);
  assign n2510 = (x0 | x1 | x2 | x3 | ~x6) & (x6 | ((x0 | ~x1 | ~x2 | ~x3) & (~x0 | (x1 ? (x2 | ~x3) : (~x2 | x3)))));
  assign n2511 = (x0 | ~x1 | ~x4 | x5 | x6) & (~x6 | ((~x0 | (x1 ? (x4 | x5) : (~x4 | ~x5))) & (x0 | x1 | x4 | x5)));
  assign z116 = n2513 | ~n2518 | ~n2525 | (~x5 & ~n2516);
  assign n2513 = ~x1 & ((~x3 & ~n2515) | (n1183 & n2514));
  assign n2514 = x3 & ~x0 & ~x2;
  assign n2515 = (x0 | ~x2 | x5 | (x4 ^ x7)) & (x2 | ((x0 | x4 | ~x5 | x7) & (~x4 | (x0 ? (~x5 ^ x7) : (x5 ^ x7)))));
  assign n2516 = ~n2517 & (x0 | ((~n269 | ~n1498) & ~n632));
  assign n2517 = n394 & n308 & n588;
  assign n2518 = n2520 & n2521 & ~n2523 & (n2519 | n2524);
  assign n2519 = x4 ? (~x5 | x6) : (x5 | ~x6);
  assign n2520 = (~n394 | ~n890) & (n736 | n409 | n607);
  assign n2521 = (n436 | n1119 | n2299) & (n310 | n2522);
  assign n2522 = (x0 | ~x1 | ~x2 | ~x4) & (~x0 | x1 | x2 | x4);
  assign n2523 = ~n542 & ((n364 & n1458) | (n300 & n429));
  assign n2524 = (~x0 | ~x1 | x2 | ~x3 | x7) & (x0 | x1 | ~x2 | x3 | ~x7);
  assign n2525 = n2527 & (~x5 | ~n601 | n2526);
  assign n2526 = (~x3 | ((~x1 | ~x2 | ~x6 | x7) & (x1 | x2 | x6 | ~x7))) & (~x1 | x2 | x3 | (~x6 ^ x7));
  assign n2527 = (n602 | n2529) & (x4 | ~n620 | n2528);
  assign n2528 = (~x0 | x2 | ~x5 | x7) & (x0 | ~x7 | (x2 ^ ~x5));
  assign n2529 = (x0 | ~x1 | x2 | ~x3 | x7) & (~x0 | ~x7 | (x1 ? (x2 | ~x3) : (~x2 | x3)));
  assign z117 = ~n2537 | (x6 ? ~n2534 : ~n2531);
  assign n2531 = (~x1 | x7 | n2533) & (~x7 | ((~n330 | n2532) & (x1 | n2533)));
  assign n2532 = (x1 | ~x2 | ~x3 | ~x5) & (~x1 | x2 | x3 | x5);
  assign n2533 = (~x2 | x3 | ~x4 | x5) & (x0 | ~x3 | ~x5 | (~x2 ^ x4));
  assign n2534 = (~n790 | ~n443 | ~n359) & (~x2 | n2535);
  assign n2535 = (n2340 | n2536) & (x7 | n677 | ~n1706);
  assign n2536 = x0 ? (x1 | x7) : (~x1 | ~x7);
  assign n2537 = ~n2540 & n2541 & (~x0 | (~n2538 & ~n2539));
  assign n2538 = ~x2 & ((n301 & n923) | (x1 & ~n1670));
  assign n2539 = n438 & ((x3 & ~x4 & x5 & x6) | (~x3 & ~x5 & (x4 ^ ~x6)));
  assign n2540 = n282 & ((~x3 & n424) | (~x0 & x3 & ~n677));
  assign n2541 = ~n2543 & (x2 | n2542) & (~n441 | n2544);
  assign n2542 = x1 ? (x3 ? (~x4 | x5) : ((~x4 | ~x5) & (x0 | x4 | x5))) : ((x3 | ~x4 | x5) & (x4 | ~x5 | ~x0 | ~x3));
  assign n2543 = ~n467 & ((n725 & n1019) | (~x1 & ~n1249));
  assign n2544 = (~x2 | ~x3 | x4 | ~x5 | ~x6) & ((x4 ^ x6) | (x2 ? (x3 | x5) : (~x3 | ~x5)));
  assign z118 = n2550 | ~n2552 | (~x3 & ~n2546);
  assign n2546 = (~x0 | n2547) & (x0 | ~x5 | ~x6 | n2549);
  assign n2547 = (~x1 | x2 | ~x4 | ~n294) & (x4 | n2548);
  assign n2548 = (~x1 | ((~x2 | ~x5 | ~x6 | ~x7) & (x6 | x7 | x2 | x5))) & (x1 | ~x2 | x5 | ~x6 | x7);
  assign n2549 = (x1 | ~x2 | x4 | x7) & (x2 | ~x4 | ~x7);
  assign n2550 = ~n688 & (x6 ? ~n2551 : ~n469);
  assign n2551 = (x0 & (x1 | (x3 & x5))) | (~x2 & (x3 | x5)) | (x2 & ~x3 & ~x5) | (x3 & ((x1 & x5) | (~x0 & ~x1 & ~x5)));
  assign n2552 = n2558 & n2559 & (x5 ? n2556 : n2553);
  assign n2553 = (~x6 | n2554) & (~x3 | x6 | n2555);
  assign n2554 = x0 ? (~x1 | x3 | (~x2 ^ x4)) : (~x3 | ((x2 | ~x4) & (x1 | ~x2 | x4)));
  assign n2555 = x4 ? (~x2 | (x0 & x1)) : x2;
  assign n2556 = x3 ? (~x6 | n2557) : (x6 | (n2557 & (~n441 | n1011)));
  assign n2557 = (x4 & (~x2 | (x0 & x1))) | (~x0 & ~x1) | (x2 & ~x4);
  assign n2558 = (~n595 | ~n1284) & (~n789 | ~n356 | ~n428);
  assign n2559 = ~n2562 & (n2561 | (~n2431 & ~n2560));
  assign n2560 = x3 & (~x5 ^ ~x6);
  assign n2561 = (x0 | ~x1 | ~x2 | x4 | x7) & (~x0 | ((x2 | ~x4 | ~x7) & (x4 | x7 | x1 | ~x2)));
  assign n2562 = ~x0 & (n2564 | (x5 & n923 & ~n2563));
  assign n2563 = x2 ? (~x4 | ~x7) : (x4 | x7);
  assign n2564 = ~x3 & ~x5 & (x2 ? (~x4 & ~x7) : (x4 & x7));
  assign z119 = ~n2572 | (~x4 & (~n2567 | (~n542 & ~n2566)));
  assign n2566 = (x0 | x1 | x3 | ~x5) & (x5 | (x0 ? (x1 ? (~x2 | x3) : (x2 | ~x3)) : (~x1 | ~x3)));
  assign n2567 = (~x6 | x7 | ~n359 | ~n464) & (x6 | n2568);
  assign n2568 = n2570 & (~x7 | n467 | (n470 & ~n2569));
  assign n2569 = ~x2 & x0 & x1;
  assign n2570 = x0 | (x1 ? ~n2571 : (~x2 | ~n2220));
  assign n2571 = ~x7 & x3 & x5;
  assign n2572 = ~n2573 & ~n2577 & ~n2581 & (n565 | n2579);
  assign n2573 = ~n498 & (n2574 | n2576 | (n626 & ~n2575));
  assign n2574 = ~n271 & ((x4 & (~x6 ^ x7)) | (~x7 & (x0 ? ~x6 : (~x4 & x6))));
  assign n2575 = (x1 | x2) & (x0 | ~x1 | ~x2);
  assign n2576 = n1683 & ((x2 & ~x7 & ~x0 & x1) | (x0 & (x1 ? (~x2 & x7) : ~x7)));
  assign n2577 = ~n566 & ((n1114 & n622) | (~x2 & ~n2578));
  assign n2578 = (x3 | ~x4 | ~x6 | x7) & (~x3 | x6 | ((~x4 | ~x7) & (x1 | x4 | x7)));
  assign n2579 = (x3 | n2580) & (~x3 | ~x4 | x5 | n2052);
  assign n2580 = (~x0 | ~x1 | ~x2 | x4 | ~x5) & (x0 | ((~x4 | ~x5) & (x4 | x5 | x1 | x2)));
  assign n2581 = ~n2582 & ((x2 & x4 & ~x6) | (~x4 & x6));
  assign n2582 = x0 ? ((~x5 | ~x7 | x1 | ~x3) & (x5 | x7 | ~x1 | x3)) : (~x3 | ~x7 | (~x1 ^ ~x5));
  assign z120 = ~n2592 | (x1 ? ~n2584 : (n2588 | n2590));
  assign n2584 = ~n2585 & (~n329 | ~n876) & (x4 | n2587);
  assign n2585 = ~x3 & ((n280 & n898) | (n330 & ~n2586));
  assign n2586 = (x2 | x5 | ~x6 | ~x7) & (~x2 | (x5 ? (~x6 | ~x7) : (x6 | x7)));
  assign n2587 = (~x5 | ~x7 | x0 | ~x2) & (x2 | ((x6 | x7 | ~x0 | x5) & (~x5 | ~x6 | ~x7)));
  assign n2588 = x4 & ((~x7 & ~n2589) | (~x0 & n875));
  assign n2589 = (~x0 | ~x2 | ~x3 | ~x5 | ~x6) & (x6 | ((x2 | x3 | x5) & (x0 | (x5 & (x2 | ~x3)))));
  assign n2590 = ~x4 & ((n324 & n876) | (x7 & ~n2591));
  assign n2591 = x0 ? (~x6 | ((~x2 | ~x3) & ~x5)) : (x5 | x6 | (x2 ^ ~x3));
  assign n2592 = (n555 | n2593) & (n1291 | (~n2594 & n2595));
  assign n2593 = (x0 | ~x1 | ~x2 | ~x3 | ~x4) & ((x1 & x2) | (~x0 ^ ~x4));
  assign n2594 = ~x1 & ((n324 & n590) | (n367 & ~n986));
  assign n2595 = ~n2597 & n2598 & (~x0 | x4 | ~n2596);
  assign n2596 = ~x6 & (~x1 ^ ~x2);
  assign n2597 = ~x4 & n480 & (x2 ? ~x3 : (x3 & x6));
  assign n2598 = (x0 | ((~x4 | ~x6) & (~x1 | x4 | x6))) & (x1 | x2 | ((~x4 | ~x6) & (~x0 | x4 | x6)));
  assign z121 = n2610 | n2613 | (x4 ? ~n2604 : ~n2600);
  assign n2600 = x0 ? n2601 : (n2603 & (x1 | n2602));
  assign n2601 = (x2 | x3 | n555) & (x1 | (n555 & (~x2 | x3 | n2360)));
  assign n2602 = (x2 | x3 | x5 | ~x6 | ~x7) & (~x2 | ~x3 | (x5 ? (x6 | x7) : (~x6 | ~x7)));
  assign n2603 = (x1 | ~x2 | n563) & (x2 | ((~x3 | n563) & (~x1 | (n563 & (x3 | ~n313)))));
  assign n2604 = n2607 & (x0 | (n2606 & (~x2 | n2605)));
  assign n2605 = (~x1 | ~x3 | ~x5 | x6 | ~x7) & (x1 | ((x6 | x7 | x3 | ~x5) & (~x6 | ~x7 | ~x3 | x5)));
  assign n2606 = (~n294 & ~n556) | (n271 & (~n272 | ~n294));
  assign n2607 = (n998 | n2608) & (~n363 | n2609);
  assign n2608 = (x0 | x1 | ~x3 | ~x5 | x7) & (~x0 | ((~x5 | ~x7 | x1 | ~x3) & (x3 | x5 | x7)));
  assign n2609 = x2 ? ((x5 | ~x6 | x7) & (x3 | ~x5 | ~x7)) : ((~x5 | x6 | ~x7) & (~x3 | x5 | x7));
  assign n2610 = ~n565 & (n2611 | ~n2612);
  assign n2611 = ~x0 & ((x1 & x2 & ~x5) | (~x3 & x5 & ~x1 & ~x2));
  assign n2612 = ~x5 | ~n480 | (x2 ^ (~x3 & ~x4));
  assign n2613 = ~n542 & (n2614 | ~n2616 | (n330 & ~n2615));
  assign n2614 = ~x1 & (x0 ? (x2 ? (x3 & ~x5) : (~x3 & x5)) : (~x5 & (~x2 ^ ~x3)));
  assign n2615 = (~x1 | ~x2 | x3 | x5) & (x1 | x2 | ~x3 | ~x5);
  assign n2616 = (~x0 | ~x1 | x2 | x5) & (x0 | (x1 ? ~x5 : (x2 | ~n1265)));
  assign z122 = ~n2620 | ~n2628 | (x4 ? ~n2619 : ~n2618);
  assign n2618 = (~x0 | ((x3 | x6 | x1 | ~x2) & (~x3 | ~x6 | ~x1 | x2))) & (~x1 | ~x2 | x3 | ~x6) & (x0 | (x1 ? (x2 ? ~x6 : (x3 | x6)) : (x2 ? (~x3 | x6) : (x3 | ~x6))));
  assign n2619 = (~x0 | x2 | ~x3 | (~x1 ^ ~x6)) & (~x2 | ((x3 | x6 | ~x0 | x1) & (x0 | (x1 ? (x3 | ~x6) : (~x3 | x6)))));
  assign n2620 = ~n2621 & ~n2626 & (~n329 | n2627);
  assign n2621 = ~x4 & (n2623 | n2625 | (~n542 & ~n2622));
  assign n2622 = (x2 | ~x3 | x0 | ~x1) & (~x0 | ((~x3 | ~x5 | x1 | ~x2) & (~x1 | x2 | x3)));
  assign n2623 = ~n2624 & ~x3 & n387;
  assign n2624 = (x2 | ~x5 | ~x6 | ~x7) & (~x2 | x5 | x6 | x7);
  assign n2625 = n400 & n717 & n394;
  assign n2626 = x0 & ((n1658 & n458) | (n301 & n1986));
  assign n2627 = (~x1 | ~x2 | ~x3 | x5 | ~x6) & (x1 | x3 | (x2 ? (~x5 | x6) : (x5 | ~x6)));
  assign n2628 = ~n2629 & (~x4 | (~n2632 & (n542 | n2631)));
  assign n2629 = ~n565 & ((n514 & n612) | n2630);
  assign n2630 = ~x1 & ((~x0 & (x2 ? (~x3 & ~x4) : x3)) | (~x2 & (x3 ? ~x4 : x0)));
  assign n2631 = (~x0 | x1 | ~x2 | ~x3) & (~x1 | x2 | (x0 & (x3 | x5)));
  assign n2632 = ~x3 & ((n364 & n921) | n2633);
  assign n2633 = n441 & (x2 ? (~x5 & n308) : (x5 & n521));
  assign z123 = ~n2639 | (~x5 & ~n2635) | (x5 & n339 & ~n2638);
  assign n2635 = ~n2637 & (~x2 | (~n2636 & (~x0 | n1692)));
  assign n2636 = n285 & (x1 ? (~x4 & n521) : (x4 & ~n565));
  assign n2637 = n359 & n996;
  assign n2638 = (x0 | x1 | ~x4 | ~x6 | ~x7) & (~x1 | (x0 ? (~x4 | (~x6 ^ x7)) : (x4 | (x6 ^ x7))));
  assign n2639 = n2641 & ~n2644 & ~n2645 & (~x4 | n2640);
  assign n2640 = (x2 | (x0 ? (~x3 | x7) : (x1 ? (~x3 | ~x7) : (x3 | x7)))) & (~x0 | x1 | ~x2 | (x3 ^ x7));
  assign n2641 = ~n2642 & (x4 | n2524) & (~n339 | n2643);
  assign n2642 = ~n1597 & (x0 ? (~x1 & n1151) : (x1 & ~n478));
  assign n2643 = (~x0 | ~x1 | ~x4 | x5 | ~x7) & (x0 | x4 | x7 | (~x1 ^ x5));
  assign n2644 = ~n478 & (x0 ? (~x3 & ~x4) : (~x1 & x3));
  assign n2645 = x2 & (n2646 | (x5 & n285 & n1065));
  assign n2646 = ~n1034 & x3 & ~n570;
  assign z124 = ~n2657 | ~n2651 | n2648 | n2650;
  assign n2648 = ~x3 & (x4 ? ~n2649 : (n387 & n1121));
  assign n2649 = x0 ? (x2 | (x1 ? (~x5 | ~x6) : (x5 | x6))) : (~x2 | (x1 ? (~x5 | x6) : (x5 | ~x6)));
  assign n2650 = ~x2 & (x0 ? (x1 ? (x3 & ~x4) : (~x3 ^ x4)) : (x1 ? (~x3 & x4) : (x3 & ~x4)));
  assign n2651 = ~n2654 & n2655 & (n2652 | ~n2653);
  assign n2652 = (~x1 | ~x2 | x3 | ~x6 | x7) & (x1 | x2 | (x3 ? (x6 | x7) : (~x6 | ~x7)));
  assign n2653 = x5 & ~x0 & x4;
  assign n2654 = n624 & (x0 ? (~x1 & ~n498) : (x1 & n314));
  assign n2655 = (~n295 | ~n757) & (n826 | ~n2656);
  assign n2656 = x3 & ~x1 & x2;
  assign n2657 = x4 ? n2658 : ((~n394 | ~n882) & ~n2659);
  assign n2658 = (~x0 | ~x1 | x2 | ~x3 | x5) & (x0 | ((~x3 | x5 | x1 | x2) & (~x2 | (x1 ? (x3 ^ x5) : (x3 | ~x5)))));
  assign n2659 = ~x5 & ((n387 & ~n2661) | (x0 & ~n2660));
  assign n2660 = (x1 | ~x2 | ~x3 | ~x6 | ~x7) & (~x1 | x2 | x3 | x6 | x7);
  assign n2661 = (~x6 | x7 | x2 | ~x3) & (~x2 | x3 | x6 | ~x7);
  assign z125 = ~n2663 | n2676 | (~x2 & ~n2674);
  assign n2663 = ~n2664 & ~n2666 & n2669 & (n444 | n2668);
  assign n2664 = ~x0 & ((~x1 & ~n2665) | (n628 & n764));
  assign n2665 = (x2 | ~x3 | x4 | ~x5 | x6) & (~x2 | ~x4 | (x3 ? (~x5 | x6) : (x5 | ~x6)));
  assign n2666 = x0 & ((n1658 & n764) | (n709 & ~n2667));
  assign n2667 = (x2 | (x1 ? (x4 ^ x5) : (~x4 | x5))) & (x4 | ~x5 | x1 | ~x2);
  assign n2668 = (x1 | x2 | ~x3 | ~x4 | ~x5) & (x3 | x4 | (x1 ? (~x2 ^ x5) : (x2 | x5)));
  assign n2669 = ~n2671 & ~n2672 & n2673 & (x1 | n2670);
  assign n2670 = (x0 | ~x2 | ~x3 | ~x4 | x5) & (x2 | (~x3 ^ x5) | (~x0 ^ ~x4));
  assign n2671 = ~n1503 & ((n363 & n1270) | (n387 & n609));
  assign n2672 = ~n677 & ((n423 & n480) | (n782 & ~n954));
  assign n2673 = (n405 | n668) & (~n514 | ~n1458);
  assign n2674 = (~n335 | n2675) & (~x5 | n967 | n1163);
  assign n2675 = (x0 | ~x1 | ~x3 | ~x6 | ~x7) & (x3 | ((x0 | x1 | x6 | ~x7) & (~x0 | (x1 ? (x6 | ~x7) : (~x6 | x7)))));
  assign n2676 = x2 & ((~x4 & ~n2677) | (n1063 & n1476));
  assign n2677 = (x3 | n2678) & (~n382 | n1255 | x0 | ~x3);
  assign n2678 = (~x0 | ((x1 | ~x5 | x6 | ~x7) & (~x1 | x5 | ~x6 | x7))) & (x0 | ~x1 | x5 | x6 | ~x7);
  assign z126 = n2680 | ~n2682 | n2691 | (n387 & ~n2695);
  assign n2680 = ~x1 & (x0 ? ~n1237 : ~n2681);
  assign n2681 = (~x4 | (x2 ? (x6 | (~x3 ^ x5)) : (x3 ? (~x5 | ~x6) : x5))) & (x5 | ~x6 | (x2 ? (~x3 | x4) : x3));
  assign n2682 = n2686 & (n379 | n2683) & (~x1 | n2684);
  assign n2683 = (x4 | (x0 ? (x1 ? (x2 | ~x3) : (~x2 | x3)) : (x1 ? (x2 ^ x3) : (x2 | ~x3)))) & (~x0 | x2 | ~x4 | (~x1 ^ x3));
  assign n2684 = ~n2685 & (n315 | n1670) & (~n312 | ~n512);
  assign n2685 = n329 & (x2 ? ~n966 : (x5 & ~n1163));
  assign n2686 = ~n2687 & ~n2689 & (n978 | n2688);
  assign n2687 = ~n534 & ((~x1 & (x0 ? (~x2 ^ x3) : (x2 & ~x3))) | (~x2 & x3 & ~x0 & x1));
  assign n2688 = (~x0 | ~x5 | (x1 ? (x2 | ~x3) : (~x2 | x3))) & (x5 | (~x1 ^ x3) | (x0 ^ ~x2));
  assign n2689 = ~n2690 & ((n717 & n718) | (n382 & n913));
  assign n2690 = (x0 | x2 | ~x3 | x5) & (~x0 | x3 | (~x2 ^ x5));
  assign n2691 = ~x1 & ((n270 & n344) | n2692 | n2694);
  assign n2692 = x5 & ((~x7 & ~n2693) | (n2131 & n2514));
  assign n2693 = (x0 | ~x2 | x3 | x4 | ~x6) & (~x0 | ((x4 | ~x6 | x2 | x3) & (~x2 | ~x3 | ~x4 | x6)));
  assign n2694 = ~n2504 & ((n313 & n330) | (~x0 & n1611));
  assign n2695 = (~x4 | x5 | x6 | ~n2696) & (~x5 | n2697);
  assign n2696 = ~x7 & (x2 ^ ~x3);
  assign n2697 = (x2 | ~x3 | x4 | ~x6 | x7) & (~x7 | ((~x2 | (x3 ? (x4 | x6) : (~x4 | ~x6))) & (x2 | x3 | ~x4 | x6)));
  assign z127 = ~n2703 | ~n2714 | (~x2 & (n2699 | n2701));
  assign n2699 = ~x4 & (n2700 | (~x5 & n387 & ~n1262));
  assign n2700 = ~n409 & ((n328 & n923) | (n327 & n625));
  assign n2701 = ~n2702 & x5 & n588;
  assign n2702 = (x0 | x1 | x6 | ~x7) & (~x0 | (x1 ? (~x6 | ~x7) : (x6 | x7)));
  assign n2703 = n2705 & n2708 & (n736 | n2704);
  assign n2704 = (x5 | ((~x0 | x1 | x3 | ~x6) & (x0 | (x1 ? (~x3 | ~x6) : (x3 | x6))))) & (~x0 | ~x5 | ~x6 | (x1 ^ ~x3));
  assign n2705 = ~n2707 & (n731 | n2706) & (~n300 | ~n1687);
  assign n2706 = (x0 | ~x1 | x2 | ~x4 | ~x5) & (~x0 | x5 | (x1 ? (x2 | x4) : (~x2 | ~x4)));
  assign n2707 = ~n2267 & ((x0 & ~x1 & x5 & ~x6) | (~x0 & (x1 ? (~x5 & ~x6) : x6)));
  assign n2708 = ~n2709 & (n542 | (~n2711 & n2712));
  assign n2709 = x1 & ((~x6 & ~n2710) | (n273 & n344));
  assign n2710 = x0 ? (x2 | (x3 ? ~x4 : (x4 | ~x5))) : (~x2 | ~x5 | (x3 ^ x4));
  assign n2711 = ~n736 & ((~x0 & ~x1 & ~x3 & x5) | (x0 & ~x5 & (~x1 ^ ~x3)));
  assign n2712 = (x1 | n2713) & (~x5 | n2267 | x0 | ~x1);
  assign n2713 = (~x0 | x2 | x3 | x4) & (x0 | ~x2 | ~x3 | ~x4 | ~x5);
  assign n2714 = (~x2 | n2718) & (n565 | (n2716 & (x2 | n2715)));
  assign n2715 = (x0 | ~x1 | x3 | ~x4 | x5) & (~x5 | ((x0 | x1 | x3 | x4) & (~x0 | (x1 ? (~x3 | x4) : (x3 | ~x4)))));
  assign n2716 = x3 ? (x4 ? n2717 : (~n782 | n1255)) : (x4 | n2717);
  assign n2717 = (~x0 | x1 | ~x2 | ~x5) & (x0 | x5 | (x1 ^ x2));
  assign n2718 = ~n2719 & (~n593 | ~n728);
  assign n2719 = ~x1 & (x5 ? ~n2720 : (n329 & ~n1262));
  assign n2720 = (~x0 | ((~x6 | ~x7 | x3 | ~x4) & (x6 | x7 | ~x3 | x4))) & (x0 | ~x3 | x4 | x6 | ~x7);
  assign z128 = ~n2726 | ~n2732 | (x7 & ~n2722);
  assign n2722 = (~x4 | n2724) & (x2 | x4 | n467 | n2723);
  assign n2723 = ~x1 ^ ~x6;
  assign n2724 = (~x5 | n2723 | x2 | ~x3) & (~x2 | n2725);
  assign n2725 = (x0 | ~x1 | x3 | (~x5 ^ x6)) & (x1 | ((x3 | x5 | x6) & (~x0 | ~x6 | (x3 ^ ~x5))));
  assign n2726 = ~n2730 & (n1527 | n2729) & (x7 | n2727);
  assign n2727 = (~n327 | ~n443 | ~n394) & (~n339 | n2728);
  assign n2728 = x1 ? (~x6 | ((x4 | x5) & (x0 | ~x4 | ~x5))) : (x6 | ((~x4 | ~x5) & (~x0 | x4 | x5)));
  assign n2729 = (x1 | x4 | x5 | ~x7) & (~x4 | (x1 ? (~x5 | x7) : (x5 ^ x7)));
  assign n2730 = ~n1977 & ((n413 & n629) | (~x7 & ~n2731));
  assign n2731 = x2 ? ((x3 | ~x4 | x5) & (x4 | ~x5 | x0 | ~x3)) : (~x3 | (x4 ^ x5));
  assign n2732 = x5 ? n2735 : (x1 ? n2733 : n2734);
  assign n2733 = x2 ? (x4 | ((x3 | ~x7) & (x0 | ~x3 | x7))) : (~x4 | (~x3 ^ x7));
  assign n2734 = (~x4 | ~x7 | x2 | ~x3) & (x4 | x7 | ~x2 | x3) & ((~x4 ^ x7) | (x0 ? (~x2 | ~x3) : (x2 | x3)));
  assign n2735 = ~n2737 & (~n742 | ~n842) & (x1 | n2736);
  assign n2736 = (x4 | x7 | x2 | ~x3) & (x3 | ((~x2 | x4 | ~x7) & (x0 | ~x4 | (~x2 ^ x7))));
  assign n2737 = ~n487 & (x0 ? ~n468 : n718);
  assign z129 = ~n2741 | (~x3 & (n2739 | (n284 & ~n2740)));
  assign n2739 = ~n478 & ((n1039 & n329) | (~x4 & ~n379));
  assign n2740 = (~x0 | x1 | x2 | x6 | ~x7) & (~x6 | ((~x0 | ((x2 | x7) & (x1 | ~x2 | ~x7))) & (~x1 | ((x2 | x7) & (x0 | ~x2 | ~x7)))));
  assign n2741 = n2744 & ((x0 & x1 & n2743) | (n2742 & (~x0 | ~x1)));
  assign n2742 = x2 ? (x3 ? (x4 ? (~x5 | x6) : (x5 ^ x6)) : (x4 ? (x5 | ~x6) : (~x5 | x6))) : (x4 ? ((x5 | x6) & (~x3 | ~x5 | ~x6)) : (x5 | ~x6));
  assign n2743 = (x6 | ((~x2 | x3 | x4 | ~x5) & (x2 | ~x4 | (x3 & x5)))) & (x2 | ~x6 | ((~x3 | ~x4 | ~x5) & (x4 | x5)));
  assign n2744 = (~n2745 | n2746) & (~n327 | ~n356 | ~n359);
  assign n2745 = x3 & (x4 ? (~x5 & x6) : (x5 & ~x6));
  assign n2746 = x7 ? (~x2 | (x0 & x1)) : x2;
  assign z130 = n2748 | ~n2754 | ~n2756 | (~n542 & ~n2752);
  assign n2748 = ~n271 & ((n921 & n2749) | ~n2750 | n2751);
  assign n2749 = x4 & ~x0 & x3;
  assign n2750 = (x3 | ~x4 | ~x5 | x6 | ~x7) & (~x3 | ((~x4 | x5 | x6 | ~x7) & (x4 | ~x6 | x7)));
  assign n2751 = ~n542 & ((x0 & n314) | n400 | n669);
  assign n2752 = (~x5 | n2753) & (n2575 | (x3 ? x5 : ~n424));
  assign n2753 = (~x0 | ~x1 | ~x2 | x3 | x4) & (x0 | x1 | x2 | ~x3 | ~x4);
  assign n2754 = (~n592 | ~n296) & (n498 | n978 | n2755);
  assign n2755 = x2 & x0 & x1;
  assign n2756 = ~n2757 & (n2575 | n2750);
  assign n2757 = n403 & ((n387 & n301) | (x0 & ~n2758));
  assign n2758 = (~x1 | ~x2 | x4 | x5 | x6) & (x1 | x2 | ~x4 | ~x5 | ~x6);
  assign z131 = ~n2767 | n2766 | n2760 | n2764;
  assign n2760 = ~x7 & ((n519 & n2761) | (~x3 & ~n2762));
  assign n2761 = (~x4 | x5) & (x4 | ~x5) & (~x0 | ~x1 | ~x2);
  assign n2762 = (~n764 | ~n742) & (~x6 | (~n2761 & ~n2763));
  assign n2763 = ~x5 & ~x4 & x2 & x0 & x1;
  assign n2764 = ~n614 & ((n428 & n1768) | (~x0 & ~n2765));
  assign n2765 = (x6 | x7) & (x1 | ~x6 | (x2 & x3) | ~x7);
  assign n2766 = ~n271 & ((~x4 & n308) | (x0 & n626));
  assign n2767 = n2770 & (~x7 | n2768) & (~n399 | n2769);
  assign n2768 = (x0 | ~x1 | ((~x4 | ~x6) & (~x2 | x4 | x6))) & (x1 | x2 | ((x4 | x6) & (~x0 | ~x4 | ~x6)));
  assign n2769 = (x1 | x2 | ~x3 | ~x4 | x7) & (~x1 | ~x2 | x3 | x4 | ~x7);
  assign n2770 = ~n717 | ((~n300 | ~n588) & (~n424 | ~n1284));
  assign z132 = ~n2774 | (~x1 & ((n595 & n713) | n2772));
  assign n2772 = n2773 & (n319 | (n339 & n512));
  assign n2773 = ~x0 & x7;
  assign n2774 = ~n2775 & n2779 & (~n981 | (~n2596 & ~n2778));
  assign n2775 = ~n570 & ((~n687 & n507) | ~n2776 | n2777);
  assign n2776 = x0 ? ((~x6 & (x2 | x3)) | (x1 & (x2 | ~x6))) : (~x1 & (x6 | (~x2 & ~x3)));
  assign n2777 = n330 & (x3 ? (~x6 & n408) : (x6 & n282));
  assign n2778 = ~x6 & ((x1 & x2 & ~x3 & ~x4) | (~x1 & ~x2 & x3 & x4));
  assign n2779 = ~n2780 & ((x3 & x4) | ~n587 | ~n300);
  assign n2780 = x6 & ~x5 & ~x2 & ~x0 & ~x1;
  assign z133 = n2782 | ~n2784 | ~n2785 | (~n271 & ~n389);
  assign n2782 = x0 & ((n282 & n2783) | (n272 & n634));
  assign n2783 = ~x3 & ~x4 & (~x6 ^ x7);
  assign n2784 = ~x0 | x1 | x2 | (~n717 & ~n1766);
  assign n2785 = ~n2787 & ~n2788 & (~n1052 | ~n2786);
  assign n2786 = x3 & ~x2 & x0 & ~x1;
  assign n2787 = ~x0 & ((~x1 & ~x6 & x7) | (x6 & (x1 ^ (~x2 & ~x7))));
  assign n2788 = n278 & ((n1063 & n875) | (n457 & n876));
  assign z134 = ~n2791 | (~x1 & ((n413 & n1422) | n2790));
  assign n2790 = n366 & (x0 ? (x3 & ~n1291) : (~x3 & n790));
  assign n2791 = ~n2792 & ~n2796 & n2797 & (~n441 | n2794);
  assign n2792 = ~x7 & (n2793 | (~x0 & ~x1 & ~n986));
  assign n2793 = x0 & ((x3 & x4 & ~x1 & ~x2) | (x1 & x2 & ~x3 & ~x4));
  assign n2794 = (x2 | x3 | x4 | ~n280) & (~x2 | ~x3 | ~x4 | ~n2795);
  assign n2795 = x5 & (~x6 ^ x7);
  assign n2796 = ~x1 & ((~x3 & x7 & x0 & ~x2) | (~x0 & ~x7 & (~x2 ^ ~x3)));
  assign n2797 = (~x0 | x7 | (x1 ^ ~x2)) & ~n1420 & (x0 | ~x1 | ~x7);
  assign z135 = ~n2802 | (~x1 & (~n2799 | ~n2800)) | ~n2804;
  assign n2799 = (x0 | x2 | x3 | x4 | ~x5) & (~x3 | ((x0 | x2 | x4 | x5) & (~x0 | (x2 ? (~x4 | x5) : (x4 | ~x5)))));
  assign n2800 = x0 ? (~n340 | ~n320) : (~x6 | n2801);
  assign n2801 = (~x2 | ~x3 | ~x4 | ~x5) & (x2 | x3 | x4 | x5);
  assign n2802 = n2803 & (n736 | n1468) & (~n990 | ~n1476);
  assign n2803 = (x2 | ~x3 | x0 | ~x1) & (~x0 | x1 | ~x2 | x3);
  assign n2804 = ~n2805 & (~n285 | ~n328 | n2806);
  assign n2805 = ~x0 & ~x2 & ~x3 & (x1 ^ x4);
  assign n2806 = (~x1 | ~x2 | ~x4 | x7) & (x1 | x2 | x4 | ~x7);
  assign z136 = n2808 | n2812 | (~x1 & ~n2810);
  assign n2808 = n782 & (x1 ? ~n2809 : (n588 & n556));
  assign n2809 = (x3 & x4 & x5 & x6 & x7) | (~x3 & (~x4 | (~x5 & ~x6 & ~x7)));
  assign n2810 = (x2 & (x4 ? n2811 : x3)) | (~x2 & ~x3) | (x3 & ~x4 & ~n424);
  assign n2811 = (~x3 | ~x5 | ~x6 | ~x7) & (x3 | x5 | x6 | x7);
  assign n2812 = x1 & ~x2 & (~x3 | (~x4 & ~x5));
  assign z137 = ~n2819 | (~x2 & ~n2814) | (x4 & ~n2815);
  assign n2814 = (~x0 | ~x1 | ~x3 | ~x4 | x5) & (x4 | ((~x1 | x3 | x5) & (~x0 | (x5 ? ~x1 : x3))));
  assign n2815 = n2817 & (n2816 | (x0 ? (x2 | x7) : (~x2 | ~x7)));
  assign n2816 = (x3 | x5 | x6) & (~x1 | ~x3 | ~x5 | ~x6);
  assign n2817 = (~x2 | ~x7 | ~n363 | n966) & (x2 | x7 | n2818);
  assign n2818 = (~x0 | x1 | ~x3 | ~x5 | ~x6) & (x5 | x6 | x0 | x3);
  assign n2819 = n2075 & ~n2820 & (~x4 | (~n2823 & ~n2824));
  assign n2820 = ~n470 & (n2821 | (~x2 & (n1458 | n2822)));
  assign n2821 = x2 & (x3 ? (~x4 & ~x5) : (x4 & x5));
  assign n2822 = x3 & (~x4 ^ ~x5);
  assign n2823 = ~n470 & ((n587 & n426) | (n423 & n1039));
  assign n2824 = n464 & ~n678;
  assign z138 = ~n2828 | (x4 & (n2826 | (~x1 & ~n2827)));
  assign n2826 = ~n1331 & (n2333 | (x3 & ~n2360));
  assign n2827 = (~x0 | x3 | ~x5 | ~x6 | x7) & (x0 | x5 | x6 | (~x3 ^ x7));
  assign n2828 = ~n2829 & n2831 & ~n2834 & (~x4 | n2833);
  assign n2829 = ~x7 & (n2830 | (~x0 & ~n1113));
  assign n2830 = n2569 & ((x5 & ~n1597) | (x4 & ~x5 & ~n1163));
  assign n2831 = (~n270 | ~n765) & (x4 | n2832);
  assign n2832 = x5 ? (~x3 | (x0 & x1)) : (x3 | (~x0 & ~x1 & ~x6));
  assign n2833 = (x0 | x1 | ~x3 | ~x5 | ~x6) & (x3 | (x0 & x1) | (~x5 ^ x6));
  assign n2834 = n480 & n1151 & (~n668 | n754);
  assign z139 = n2836 | n2841 | n2842 | (~n350 & ~n2838);
  assign n2836 = ~x3 & ((n359 & n2837) | (n1747 & n1944));
  assign n2837 = x7 & ~x6 & x4 & ~x5;
  assign n2838 = n2839 & ~n2840 & (x2 | ~n480 | n379);
  assign n2839 = (x5 | x6 | x0 | ~x1) & (x1 | ((~x2 | x5 | x6) & (~x0 | (x5 ^ x6))));
  assign n2840 = n659 & ((n282 & n327) | (n408 & n328));
  assign n2841 = ~n534 & ~n2755;
  assign n2842 = x5 & (n2843 | (~x3 & n1019 & n742));
  assign n2843 = x6 & n329 & (~n331 | n1127);
  assign z140 = n2848 | n2849 | n2850 | (n725 & ~n2845);
  assign n2845 = ~n2846 & (~n659 | ~n556) & (n2051 | ~n2847);
  assign n2846 = x0 & ((~x5 & x6 & ~x7) | (x3 & (x5 ? (~x6 ^ x7) : (~x6 & x7))));
  assign n2847 = x4 & x0 & ~x3;
  assign n2848 = ~n1896 & (~n2051 | (n282 & n280));
  assign n2849 = ~n2051 & ((~x0 & (~x3 | ~x4)) | (~x1 & (x4 ? x0 : x3)));
  assign n2850 = n521 & ((n387 & n314) | (~x1 & ~n1974));
  assign z141 = ~n2853 | (~x6 & ((n359 & n649) | n2852));
  assign n2852 = n282 & ((n659 & n1074) | (x0 & n606));
  assign n2853 = n2854 & n2855 & ~n2856 & (~n601 | n2189);
  assign n2854 = ~n1420 & (x0 | ~n308 | (~x1 & ~x2));
  assign n2855 = (x6 & (x0 | x7)) | (x1 & x2) | (~x0 & ~x6);
  assign n2856 = ~x0 & ((n282 & n1766) | (n408 & n2857));
  assign n2857 = x7 & x3 & ~x6;
  assign z142 = ~n2861 | (~x0 & (~n2859 | (~x4 & ~n2860)));
  assign n2859 = (~x1 & (x7 | (~x2 & ~x3 & ~x4))) | (x7 & (~x2 | ~x3 | ~x4)) | (x1 & x2 & x3 & ~x7);
  assign n2860 = (x1 | x2 | x3 | ~n962) & (~x1 | ~x2 | ~x3 | ~n2795);
  assign n2861 = (~x0 | ~x7 | n2863) & (x0 | x4 | x7 | n2862);
  assign n2862 = (~x1 | ~x2 | ~x3 | x5) & (x1 | x2 | x3 | ~x5);
  assign n2863 = x1 & x2 & (x3 | x4);
  assign z143 = n2093 | ~n2865 | (n782 & n2867);
  assign n2865 = n2866 & (~n514 | ~n1259) & (~x2 | n1468);
  assign n2866 = ~x1 | (x2 & (~x0 | x3 | x4));
  assign n2867 = x3 & (x1 ? (~x4 & ~x5) : (x4 & x5));
  assign z144 = ~n2871 | (n1151 & (x0 ? ~n2869 : ~n2870));
  assign n2869 = (~x1 | x3 | ~x4 | ~x5 | x6) & (x1 | ~x3 | x4 | x5 | ~x6);
  assign n2870 = (~x1 | ~x3 | ~x4 | x5 | x6) & (x1 | ((~x3 | ~x4 | ~x5 | ~x6) & (x5 | x6 | x3 | x4)));
  assign n2871 = n1931 & ~n2873 & n2875 & (~x3 | n2872);
  assign n2872 = (~x0 | x1 | x2 | x4 | ~x5) & (x0 | ((~x1 | (x2 ? (x4 | x5) : (~x4 | ~x5))) & (x1 | ~x2 | ~x4 | x5)));
  assign n2873 = x1 & ((n301 & n661) | (n659 & ~n2874));
  assign n2874 = (x5 | ~x6 | x2 | ~x4) & (~x2 | x4 | ~x5 | x6);
  assign n2875 = (~x0 | ~x1 | x2 | ~x3) & (~x2 | x3 | (x0 & x1 & ~n411));
  assign z145 = ~n2882 | (~x5 & ~n2877) | (x1 & ~n2881);
  assign n2877 = ~n2879 & (x6 | ((~n359 | ~n2006) & ~n2878));
  assign n2878 = (n312 | n2514) & (x1 | n760) & (~x1 | n1074);
  assign n2879 = n740 & ~n2880;
  assign n2880 = (x0 | ~x1 | x3 | ~x4 | ~x7) & (~x0 | ~x3 | (x1 ? (~x4 | ~x7) : (x4 | x7)));
  assign n2881 = (x0 | ~x2 | x3 | ~x4 | x5) & (x2 | ((x4 | ~x5 | x0 | ~x3) & (~x0 | ~x4 | (x3 ^ x5))));
  assign n2882 = n2890 & ~n2888 & ~n2887 & ~n2883 & ~n2886;
  assign n2883 = ~x1 & ((~n761 & ~n2884) | (n519 & ~n2885));
  assign n2884 = x0 ? (x4 | x5) : (~x4 | ~x5);
  assign n2885 = (~x0 | ~x2 | ~x4 | ~x5) & (x0 | x2 | x4 | x5);
  assign n2886 = ~x3 & x5 & (x0 ? (x1 ^ x4) : (x1 & x4));
  assign n2887 = (~x0 ^ ~x3) & (x1 ? (~x4 & ~x5) : (x4 ^ x5));
  assign n2888 = ~n2889 & n1207 & n790;
  assign n2889 = (~x0 | ~x1 | x3 | x6) & (x0 | x1 | ~x3 | ~x6);
  assign n2890 = (~n514 | ~n1259) & (~n300 | ~n1270);
  assign z146 = ~n2905 | ~n2898 | n2892 | n2896;
  assign n2892 = ~x2 & (n2893 | (n480 & ~n2895));
  assign n2893 = ~x0 & (x1 ? (n606 & n313) : ~n2894);
  assign n2894 = (x3 | x4 | x5 | x6 | ~x7) & (~x3 | ~x4 | ~x5 | ~x6 | x7);
  assign n2895 = (x3 | ~x5 | x6 | (~x4 ^ x7)) & (~x3 | ~x4 | x5 | ~x6 | x7);
  assign n2896 = n426 & (n2897 | (~x0 & n473 & n875));
  assign n2897 = ~x6 & n1921 & (x1 ? (x4 & ~x7) : (x4 ^ ~x7));
  assign n2898 = ~n2899 & ~n2902 & (n703 | n2901);
  assign n2899 = ~n2900 & x4 & n363;
  assign n2900 = (x2 | x3 | ~x5 | x6) & (~x3 | (x6 ? x5 : ~x2));
  assign n2901 = (x0 | ~x2 | ~x3 | ~x5 | ~x6) & (~x0 | x2 | x5 | (x3 & x6));
  assign n2902 = ~x0 & ((n725 & ~n2903) | (~n1163 & ~n2904));
  assign n2903 = (~x3 | x4 | ~x5 | ~x6) & (x3 | ~x4 | x5 | x6);
  assign n2904 = (x1 | x2 | ~x4 | x5) & (~x1 | ~x2 | x4 | ~x5);
  assign n2905 = (n2158 | n2907) & (n1016 | n2906);
  assign n2906 = (x5 & ((x2 & x3) | (~x0 & x6 & (x2 | x3)))) | (~x2 & ((~x5 & ~x6) | (~x3 & (~x5 | (x0 & ~x6))))) | (x0 & ~x5 & (x3 | ~x6));
  assign n2907 = (~x0 | x1 | ~x3 | x4 | ~x6) & (x0 | ((x4 | x6 | x1 | ~x3) & (~x1 | ~x4 | (~x3 ^ x6))));
  assign z147 = n2914 | n2919 | (x0 ? ~n2924 : ~n2909);
  assign n2909 = x2 ? n2912 : (x4 ? n2910 : n2911);
  assign n2910 = (~x1 | x5 | x7 | (~x3 ^ x6)) & (~x5 | ((x1 | (x3 ? (~x6 | x7) : (x6 | ~x7))) & (~x1 | ~x3 | x6 | ~x7)));
  assign n2911 = (x1 | x3 | x5 | x6 | ~x7) & ((x5 ^ x7) | (x1 ? (x3 | ~x6) : (~x3 | x6)));
  assign n2912 = (n1291 | n2913) & (x6 | ~n588 | n1188);
  assign n2913 = (~x1 | x3 | ~x4 | ~x6) & (x1 | x4 | (~x3 ^ x6));
  assign n2914 = x3 & (~n2916 | (~x0 & ~n2915));
  assign n2915 = (x1 | x2 | ~x4 | ~x5 | x6) & (x4 | ((~x1 | x6 | (~x2 ^ ~x5)) & (x1 | x2 | ~x5 | ~x6)));
  assign n2916 = ~n2917 & ~n2918 & (~n273 | ~n364);
  assign n2917 = x6 & ((x0 & ~x1 & ~x2 & x5) | (~x0 & ((x2 & ~x5) | (x1 & ~x2 & x5))));
  assign n2918 = x0 & ~x6 & ((~x2 & ~x5) | (~x1 & x2 & x5));
  assign n2919 = ~x3 & (n2922 | n2923 | (n2920 & ~n2921));
  assign n2920 = ~x0 & x6;
  assign n2921 = (~x4 | x5 | x1 | ~x2) & (~x5 | (x1 ? (x2 ^ ~x4) : (x2 | x4)));
  assign n2922 = ~n605 & ((x0 & (~x1 | ~x4) & x6) | (~x6 & (x1 ? ~x0 : x4)));
  assign n2923 = ~n902 & (x0 ? n1494 : n1295);
  assign n2924 = n2926 & (n731 | n2925);
  assign n2925 = (~x1 | x2 | ~x4 | x5) & (x1 | x4 | (~x2 ^ ~x5));
  assign n2926 = (n791 | n1262) & (~n356 | n2927);
  assign n2927 = (~x1 | ~x2 | x5 | x6 | x7) & (x1 | x2 | ~x5 | ~x6 | ~x7);
  assign z148 = n2929 | ~n2935 | ~n2945 | (~n283 & ~n2934);
  assign n2929 = ~x3 & (n2932 | (~x6 & (n2930 | n2931)));
  assign n2930 = n2773 & ((n335 & n408) | (n282 & n284));
  assign n2931 = ~x7 & n559 & ((x2 & ~x5) | (x1 & ~x2 & x5));
  assign n2932 = ~n2933 & n521 & n387;
  assign n2933 = x2 ? (~x4 | ~x5) : (x4 | x5);
  assign n2934 = (x0 | ~x1 | x3 | (~x6 ^ x7)) & (~x3 | ((~x0 | x1 | x6 | ~x7) & (x0 | (x1 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n2935 = ~n2936 & n2937 & n2942 & (n868 | n2941);
  assign n2936 = ~n565 & ((n480 & n1453) | (n441 & n892));
  assign n2937 = ~n2938 & ~n2940 & (~n521 | ~n443 | ~n394);
  assign n2938 = ~n2939 & (x1 ? n1683 : n700);
  assign n2939 = (x3 | ~x5 | x0 | ~x2) & (~x0 | x2 | ~x3 | x5);
  assign n2940 = ~n645 & n913 & ~x5 & x6;
  assign n2941 = (~x2 | ~x3 | x4 | x6 | ~x7) & (x2 | x3 | ~x4 | (~x6 ^ x7));
  assign n2942 = (x6 | n2943) & (~x5 | ~n1064 | n2944);
  assign n2943 = x0 ? ((~x4 | ~x5 | x1 | ~x3) & (x4 | x5 | ~x1 | x3)) : ((~x1 | ~x3 | x4 | ~x5) & (~x4 | x5 | x1 | x3));
  assign n2944 = x1 ? (x2 ? (x4 | x6) : (~x4 | ~x6)) : (~x6 | (x2 ^ x4));
  assign n2945 = n2948 & (~x3 | ((~n364 | ~n714) & ~n2946));
  assign n2946 = ~x1 & (n2947 | (x0 & n366 & n294));
  assign n2947 = n521 & ((~x0 & ~x2 & x4 & x5) | (x0 & ~x5 & (~x2 ^ x4)));
  assign n2948 = ~n2949 & (n542 | (x2 & n2953) | (~x2 & n2952));
  assign n2949 = ~x0 & (x2 ? ~n2951 : ~n2950);
  assign n2950 = (x1 | ~x3 | x4 | ~x5 | ~x6) & (x6 | ((x1 | x3 | x4 | ~x5) & (~x1 | (x3 ? (x4 | x5) : (~x4 | ~x5)))));
  assign n2951 = (x1 | ~x3 | ~x4 | ~x5 | ~x6) & (~x1 | x5 | (x3 ? (~x4 | x6) : (x4 | ~x6)));
  assign n2952 = x0 ? (x3 | (x1 ? (~x4 ^ x5) : (x4 | x5))) : (x1 ? (~x3 | ~x4) : (x3 ? (x4 | x5) : (~x4 | ~x5)));
  assign n2953 = (~x0 | x1 | x3 | x4) & (x0 | ~x3 | (x1 ? (~x4 | ~x5) : x4));
  assign z149 = n2955 | n2961 | ~n2965 | (~x2 & ~n2964);
  assign n2955 = ~x1 & (~n2958 | (~x0 & ~n2956));
  assign n2956 = (x4 | n2957) & (~x3 | ~x4 | ~x7 | n903);
  assign n2957 = (x2 | ~x3 | ~x5 | x6 | x7) & (~x6 | ((x2 | x3 | x5 | ~x7) & (~x2 | (x3 ? (x5 | x7) : (~x5 | ~x7)))));
  assign n2958 = (n2107 | n2959) & (~n857 | n2960);
  assign n2959 = (~x4 | x7 | x0 | ~x3) & (~x0 | (x3 ? (x4 | ~x7) : (~x4 | x7)));
  assign n2960 = (~x2 | x5 | ~x6 | (~x4 ^ ~x7)) & (x2 | x4 | ~x5 | x6 | x7);
  assign n2961 = x1 & ((~n350 & ~n2962) | (n1837 & ~n2963));
  assign n2962 = (~x0 | x2 | x3 | ~x5 | ~x6) & (x0 | ~x3 | (x2 ? (x5 | x6) : (~x5 | ~x6)));
  assign n2963 = (~x5 | ~x7 | ~x3 | x4) & (x3 | ((x0 | x4 | x5 | ~x7) & (~x5 | x7 | ~x0 | ~x4)));
  assign n2964 = (x1 | x3 | x4 | ~x5 | ~x7) & (x5 | (x1 ? (x3 ? (x4 | ~x7) : (~x4 | x7)) : (x3 ? (x4 | x7) : (~x4 | ~x7))));
  assign n2965 = n2967 & ~n2969 & ~n2971 & (~x4 | n2966);
  assign n2966 = x1 ? (x7 | ((x2 | ~x3) & (x0 | ~x2 | x3))) : (~x7 | ((~x2 | x3) & (~x0 | x2 | ~x3)));
  assign n2967 = (~n624 | n2968) & (~x5 | n350 | ~n2656);
  assign n2968 = x1 ? (~x7 | (x0 & x3)) : (x3 | x7);
  assign n2969 = ~x7 & ((n359 & n609) | (~n2970 & ~n1548));
  assign n2970 = x2 ? (~x3 | ~x4) : (x3 | x4);
  assign n2971 = n1151 & ((n625 & ~n2884) | (n441 & n2822));
  assign z150 = ~n2982 | (x2 ? ~n2977 : (n2973 | n2975));
  assign n2973 = ~x5 & ((n387 & n842) | (~x1 & ~n2974));
  assign n2974 = (x0 | ~x3 | x4 | x6 | x7) & (~x4 | ((x0 | ~x3 | x6 | ~x7) & (~x0 | (x3 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n2975 = x5 & ((n633 & n765) | (x1 & ~n2976));
  assign n2976 = (~x0 | x3 | x6 | (x4 ^ x7)) & (~x3 | ((~x6 | x7 | ~x0 | x4) & (x0 | (x4 ? (~x6 | x7) : (x6 | ~x7)))));
  assign n2977 = x6 ? (~n2978 & ~n2980) : (x1 | n2981);
  assign n2978 = ~x0 & ((n923 & n1555) | (x1 & ~n2979));
  assign n2979 = (~x3 | ~x4 | x5 | x7) & (x3 | x4 | ~x5 | ~x7);
  assign n2980 = n363 & (x3 ? ~n1663 : n284);
  assign n2981 = (~x0 | ~x3 | x5) & (~x5 | ((x0 | ~x3 | x4 | ~x7) & (x3 | (x0 ? (x4 ^ x7) : (~x4 | x7)))));
  assign n2982 = ~n2983 & n2987 & (x0 ? n2985 : n2986);
  assign n2983 = x2 & ((~x6 & ~n2984) | (n875 & n2749));
  assign n2984 = (x0 | ~x3 | x4 | x5 | x7) & (x3 | ((~x5 | ~x7 | x0 | ~x4) & (~x0 | (x4 ? (x5 | x7) : (~x5 | ~x7)))));
  assign n2985 = (~x2 | x3 | x4 | ~x5 | ~x6) & (x2 | ((~x3 | ~x5 | (~x4 & x6)) & (x5 | ((x4 | ~x6) & (x3 | (x4 & ~x6))))));
  assign n2986 = x2 ? (x3 ? (x4 ? (x5 | x6) : (~x5 | ~x6)) : (~x5 | (x4 ^ x6))) : (x3 ? ((x5 | ~x6) & (~x4 | ~x5 | x6)) : (~x4 | x5));
  assign n2987 = (~n270 | ~n344) & (n1291 | n2988);
  assign n2988 = (~x0 | x2 | x3 | ~x4 | x6) & (x0 | x4 | (x2 ? (x3 | ~x6) : (~x3 | x6)));
  assign z151 = n2990 | ~n2995 | ~n3002 | (~x2 & ~n2993);
  assign n2990 = ~x1 & (n2991 | (~n1578 & ~n2179));
  assign n2991 = ~x3 & (x0 ? ~n2992 : (n366 & n294));
  assign n2992 = (x2 | x5 | ~x7 | (~x4 ^ ~x6)) & (~x2 | x4 | ~x5 | ~x6 | x7);
  assign n2993 = (~n1064 | n1417 | x4 | ~x6) & (~x4 | n2994);
  assign n2994 = (x0 | x1 | x3 | x5 | ~x6) & (~x1 | ~x5 | (x0 ? (x3 ^ x6) : (~x3 | x6)));
  assign n2995 = ~n2996 & ~n2997 & n3000 & (n1254 | n2999);
  assign n2996 = ~n1163 & ((x0 & ~x1 & ~x4 & ~x5) | (~x0 & (x1 ? (~x4 ^ ~x5) : (x4 & x5))));
  assign n2997 = ~n565 & (~n2998 | (x5 & n620 & ~n510));
  assign n2998 = (~x0 | x1 | ~x3 | ~x4 | x5) & (x0 | x3 | x4 | (~x1 ^ x5));
  assign n2999 = (x0 | x1 | ~x2 | x3 | x5) & (~x0 | ~x3 | (x1 ? (x2 | x5) : ~x5));
  assign n3000 = (n485 | n3001) & (~n300 | ~n1687);
  assign n3001 = (x0 | x1 | x2 | ~x3 | x5) & (~x0 | ~x2 | x3 | (~x1 ^ x5));
  assign n3002 = ~n3003 & (~x1 | ((~n713 | ~n2837) & ~n3006));
  assign n3003 = ~n542 & ((~x4 & ~n3004) | (n356 & ~n3005));
  assign n3004 = (~x1 | ((x0 | x2 | ~x3 | x5) & (~x0 | x3 | ~x5))) & (x0 | x1 | ~x3 | (~x2 & ~x5));
  assign n3005 = (~x0 | x1 | (x2 ^ ~x5)) & (~x1 | (x0 ? (x2 | x5) : (~x2 | ~x5)));
  assign n3006 = ~x0 & ((~n1254 & ~n3007) | (n556 & n1453));
  assign n3007 = (~x2 | ~x3 | x5 | x7) & (x2 | x3 | ~x5 | ~x7);
  assign z152 = ~n3010 | ~n3015 | ~n3020 | (~n566 & ~n3009);
  assign n3009 = (x2 | (x1 ? (x4 ^ x7) : (x3 | (~x4 ^ x7)))) & (x4 | x7 | ~x1 | x3) & (x1 | ~x2 | ~x3 | ~x4 | ~x7);
  assign n3010 = n3012 & (n1254 | (~n3011 & (~x0 | n2208)));
  assign n3011 = n579 & ((n789 & n923) | (x1 & n790));
  assign n3012 = (n688 | n3014) & (~n364 | ~n3013);
  assign n3013 = ~x7 & ~x5 & x3 & x4;
  assign n3014 = (~x1 | ((x3 | x5 | ~x0 | x2) & (x0 | ~x2 | ~x5))) & (~x0 | x1 | (x2 ? x5 : ~x3));
  assign n3015 = x2 ? (~n3016 & ~n3018) : (x1 | n3019);
  assign n3016 = ~x6 & (n3017 | (x0 & n276 & n1555));
  assign n3017 = x7 & ~n1278 & (~x0 ^ ~x4);
  assign n3018 = n1177 & n425 & n521;
  assign n3019 = (x0 | x3 | ~x4 | ~n313) & (~x0 | (x3 ? n1851 : (x4 | ~n313)));
  assign n3020 = ~n3023 & (x0 | (~n3022 & (x4 | n3021)));
  assign n3021 = (x1 | ~x5 | x7) & (~x3 | ((~x2 | x5 | x7) & (~x5 | ~x7 | ~x1 | x2)));
  assign n3022 = x7 & n913 & (x2 ? ~x3 : x5);
  assign n3023 = ~n836 & ((n579 & ~n3025) | (x2 & ~n3024));
  assign n3024 = (x0 | ~x1 | ~x3 | x5 | ~x7) & (x7 | ((~x0 | (x1 ? (x3 | x5) : (~x3 | ~x5))) & (x0 | x1 | x3 | x5)));
  assign n3025 = (~x1 | x3 | ~x5 | ~x7) & (x1 | ~x3 | x5 | x7);
  assign z153 = ~n3034 | ~n3039 | (x0 ? ~n3031 : ~n3027);
  assign n3027 = (x7 | n3028) & (~x6 | ~x7 | n3030);
  assign n3028 = (~x1 | x2 | x5 | n580) & (~x2 | n3029);
  assign n3029 = (x1 | ~x3 | ~x4 | x5 | ~x6) & (~x5 | ((x1 | x3 | x4 | x6) & (~x1 | ~x6 | (x3 ^ ~x4))));
  assign n3030 = (x1 | x2 | x3 | ~x4 | x5) & (~x2 | ((~x4 | ~x5 | x1 | ~x3) & (~x1 | x5 | (x3 ^ ~x4))));
  assign n3031 = (x2 | n3032) & (x1 | ~x2 | n570 | n580);
  assign n3032 = (n3033 | n966) & (x1 | ~n294 | ~n443);
  assign n3033 = x1 ? (x4 | x7) : (~x4 | ~x7);
  assign n3034 = ~n3035 & (n377 | n3037) & (x2 | n3038);
  assign n3035 = ~x6 & n340 & (n3036 | (~x0 & ~n1731));
  assign n3036 = ~x5 & ~x4 & x0 & ~x1;
  assign n3037 = (~x0 | ~x1 | ~x2 | x3 | x4) & (x0 | ~x3 | (x1 ? (~x2 | ~x4) : x2));
  assign n3038 = x0 ? ((x5 | ~x6 | x1 | x3) & (~x1 | ~x3 | ~x5 | x6)) : (x3 | ~x5 | (~x1 ^ ~x6));
  assign n3039 = n3041 & (x2 | (~n3040 & (~x0 | n2236)));
  assign n3040 = n730 & ((n276 & n521) | (n308 & n620));
  assign n3041 = n3042 & ~n3043 & ~n3044 & (n405 | n966);
  assign n3042 = (~n364 | ~n1458) & (~n300 | (~n1314 & ~n2333));
  assign n3043 = ~n435 & ((n335 & n423) | (n284 & n426));
  assign n3044 = ~n3045 & (x1 ? n314 : n400);
  assign n3045 = x0 ? (x2 | ~x4) : (~x2 | x4);
  assign z154 = ~n3059 | n3056 | n3047 | ~n3050;
  assign n3047 = ~x1 & ((n579 & ~n3049) | (x0 & ~n3048));
  assign n3048 = (~x7 | n602 | x2 | ~x3) & (~x2 | x7 | n2903);
  assign n3049 = x3 ? (x7 | (x4 ? (~x5 | ~x6) : (x5 | x6))) : (x4 | ~x7 | (x5 ^ x6));
  assign n3050 = x6 ? (x7 ? (~n3051 & n3052) : n3053) : (x7 ? n3053 : (~n3051 & n3052));
  assign n3051 = x1 & ((n647 & n429) | (n285 & ~n2933));
  assign n3052 = (x4 | ((x0 | ~x1 | ~x2 | ~x3) & (~x0 | (x1 ? (x2 | ~x3) : (~x2 | x3))))) & (x0 | x1 | ~x4 | (x2 ^ x3));
  assign n3053 = ~n3055 & (x0 ? n3054 : (~n438 | ~n613));
  assign n3054 = (~x1 | x2 | x3 | x4 | x5) & (x1 | ~x4 | (x2 ? ~x3 : (x3 | ~x5)));
  assign n3055 = ~n614 & (n594 | (~x0 & (n628 | n1114)));
  assign n3056 = x1 & ((n296 & n713) | n3057);
  assign n3057 = ~x0 & (x2 ? (n313 & n356) : ~n3058);
  assign n3058 = (~x3 | ((~x4 | ~x5 | x6 | ~x7) & (~x6 | x7 | x4 | x5))) & (x3 | x4 | ~x5 | x6 | x7);
  assign n3059 = ~n3062 & ~n3064 & (x1 ? n3060 : n3061);
  assign n3060 = (x0 | ~x2 | ~x3 | ~x4 | ~x6) & (x3 | (x0 ? (x2 ? (x4 | ~x6) : (~x4 | x6)) : (x2 ? (x4 | x6) : (~x4 | ~x6))));
  assign n3061 = x0 ? (~x4 | (x2 ? (x3 | ~x6) : (~x3 | x6))) : (~x3 | x4 | (~x2 ^ x6));
  assign n3062 = ~x3 & (n3063 | (n700 & n782 & ~n1417));
  assign n3063 = n366 & (x0 ? ~n1029 : (x5 & ~n2723));
  assign n3064 = x3 & ((n273 & n394) | (~x2 & ~n3065));
  assign n3065 = (x0 | x1 | ~x4 | x5 | ~x6) & (~x0 | ~x5 | (x1 ? (~x4 | ~x6) : (x4 | x6)));
  assign z155 = n3067 | ~n3072 | ~n3074 | (x3 & ~n3071);
  assign n3067 = ~x4 & (n3068 | (n575 & ~n3070));
  assign n3068 = ~x1 & (x6 ? ~n3069 : (n579 & ~n453));
  assign n3069 = (~x0 | ~x2 | ~x3 | ~x5 | ~x7) & (x2 | ((~x3 | x5 | x7) & (x0 | ((x5 | x7) & (x3 | ~x5 | ~x7)))));
  assign n3070 = (~x6 | x7 | x3 | ~x5) & (~x3 | x5 | (x6 ^ x7));
  assign n3071 = x2 ? ((x1 | (x4 ^ x7)) & (x0 | ~x1 | (~x4 ^ x7))) : ((x0 | x1 | ~x4 | x7) & (~x0 | ~x1 | x4 | ~x7));
  assign n3072 = (~x2 | x3 | x4 | n1318) & (x2 | (x3 ? n3073 : (~x4 | n1318)));
  assign n3073 = x1 ? (~x7 | ((~x4 | x5) & (x0 | x4 | ~x5))) : (x7 | ((x4 | ~x5) & (~x0 | ~x4 | x5)));
  assign n3074 = ~n3075 & (~x4 | (n3079 & (n565 | n3078)));
  assign n3075 = ~x3 & (n3076 | ~n3077 | (~n570 & ~n2522));
  assign n3076 = ~n1291 & ((n278 & n441) | (n366 & n480));
  assign n3077 = (~n394 | ~n1555) & (~n295 | ~n1183);
  assign n3078 = (~x0 | x1 | ~x2 | x3 | x5) & (x0 | ~x1 | x2 | ~x3 | ~x5);
  assign n3079 = ~n3080 & (n2615 | (x0 ? (x6 | x7) : (~x6 | ~x7)));
  assign n3080 = ~n1318 & n647 & x3 & n327;
  assign z156 = n3083 | n3086 | ~n3091 | (~n3082 & ~n3090);
  assign n3082 = ~x0 & ~x1;
  assign n3083 = ~x1 & ((~x3 & ~n3084) | (n659 & ~n3085));
  assign n3084 = x0 ? ((~x5 | x6 | x2 | x4) & (~x2 | x5 | ~x6)) : (x5 | (x2 ^ ~x4));
  assign n3085 = x2 ? (x6 | (x4 ^ x5)) : (x4 | ~x5);
  assign n3086 = x6 & ((n394 & n451) | n3087 | n3089);
  assign n3087 = ~x7 & ((n300 & n612) | (~x2 & ~n3088));
  assign n3088 = (x0 | ~x1 | x3 | ~x4 | x5) & (~x0 | ((~x1 | ~x3 | x4 | ~x5) & (~x4 | x5 | x1 | x3)));
  assign n3089 = ~n2615 & (x0 ? n342 : n341);
  assign n3090 = (~x2 | x3 | x4 | x5 | x6) & (x2 | (x3 ? (x4 ? (~x5 | ~x6) : (~x5 ^ x6)) : (x4 ? (x5 | x6) : (~x5 | ~x6))));
  assign n3091 = ~n3092 & (n467 | n3096) & (~n387 | n3097);
  assign n3092 = ~x6 & ((~x4 & ~n3093) | (n588 & ~n3095));
  assign n3093 = x2 ? (x7 | (n504 & (x0 | n3094))) : (~x7 | n504);
  assign n3094 = x1 ? (~x3 | x5) : (x3 | ~x5);
  assign n3095 = (x0 | x1 | x2 | x5 | x7) & (~x0 | ~x5 | (x1 ? (x2 | ~x7) : (~x2 | x7)));
  assign n3096 = (x0 | ((~x2 | ~x4) & (x4 | ~x6 | x1 | x2))) & (x1 | ~x2 | ~x4) & (~x0 | ~x1 | x2 | x4 | x6);
  assign n3097 = (x2 | ~x3 | x4 | ~x5 | ~x6) & (~x2 | ((x5 | ~x6 | x3 | x4) & (~x3 | ~x4 | ~x5 | x6)));
  assign z157 = ~n3106 | (x1 ? (n3102 | n3104) : ~n3099);
  assign n3099 = ~n3100 & (~n413 | ~n595);
  assign n3100 = ~x3 & (x0 ? (n1207 & n313) : ~n3101);
  assign n3101 = (x2 | x4 | x5 | ~x6 | x7) & (x6 | ((x2 | x4 | x5 | ~x7) & (~x2 | (x4 ? (x5 | x7) : (~x5 | ~x7)))));
  assign n3102 = ~n3103 & (x2 ? n403 : n2220);
  assign n3103 = (~x0 | x4 | x5 | ~x6) & (x0 | (x4 ? (x5 | ~x6) : (~x5 | x6)));
  assign n3104 = ~x0 & (n3105 | (x2 & n280 & n588));
  assign n3105 = n339 & (n1145 | (x4 & n851));
  assign n3106 = n3109 & (n487 | (x0 & n3107) | (~x0 & n3108));
  assign n3107 = (x5 | x6 | x1 | x4) & (~x5 | ((x1 | ((x4 | ~x6) & (~x2 | ~x4 | x6))) & (x2 | ((x4 | ~x6) & (~x1 | ~x4 | x6)))));
  assign n3108 = (~x1 | ~x2 | x4 | x5 | x6) & (x1 | ~x4 | ((~x5 | ~x6) & (x2 | x5 | x6)));
  assign n3109 = n3110 & ~n3113 & ((~x1 & x2) | n3112 | (x1 & ~x2));
  assign n3110 = (~n428 | ~n2289) & (n271 | n3111);
  assign n3111 = x3 ? ((x0 | x4 | x5 | ~x6) & (~x4 | ((x5 | x6) & (~x0 | ~x5 | ~x6)))) : (x0 ? (x4 ? (x5 | ~x6) : (~x5 | x6)) : (x4 ? (~x5 | x6) : (x5 ^ x6)));
  assign n3112 = (~x0 | x3 | x4 | ~x5 | x6) & (x0 | ((~x3 | x4 | x5 | ~x6) & (x3 | ~x5 | (~x4 ^ x6))));
  assign n3113 = x3 & (x4 ? ~n3114 : ~n3115);
  assign n3114 = (x0 | ~x1 | ((~x5 | ~x6) & (~x2 | x5 | x6))) & (x1 | (x0 ? (x2 | (x5 ^ x6)) : (x5 | ~x6)));
  assign n3115 = (x0 | x1 | x2 | ~x5 | x6) & (~x0 | x5 | (x1 ? (x2 | x6) : ~x6));
  assign z158 = n3117 | n3124 | ~n3127 | (~n542 & ~n3126);
  assign n3117 = ~x4 & (n3118 | ~n3122 | (n1747 & n3121));
  assign n3118 = x1 & ((x5 & ~n3119) | (n1921 & ~n3120));
  assign n3119 = (~x0 | ~x2 | x3 | ~x6 | ~x7) & (x0 | x7 | (x2 ? (~x3 | x6) : (x3 | ~x6)));
  assign n3120 = (x2 | ~x3 | ~x6 | ~x7) & (~x2 | x3 | x6 | x7);
  assign n3121 = ~x3 & (~x5 ^ ~x7);
  assign n3122 = (~n359 | ~n3123) & (~n382 | ~n300 | ~n465);
  assign n3123 = ~x7 & x3 & ~x5;
  assign n3124 = ~x1 & (~n3125 | (~x0 & (n1226 | n2837)));
  assign n3125 = ~x0 | (~n270 & ~n1476 & (~n278 | ~n313));
  assign n3126 = (~x5 | (x1 & x2) | (x0 ^ ~x4)) & (~x4 | x5 | (x0 ? (x1 | x2) : ~x1));
  assign n3127 = ~n3128 & ~n3131 & (n555 | n3130);
  assign n3128 = n1074 & (~n3129 | (~n881 & ~n1548));
  assign n3129 = (~n300 | ~n807) & (~n2431 | ~n364);
  assign n3130 = (~x1 | (x0 ? (x2 | ~x4) : x4)) & (x0 | ~x2 | x4) & (x1 | ((x0 | x2 | x3 | ~x4) & (~x0 | (x2 ^ x4))));
  assign n3131 = x1 & (~n3132 | (n308 & ~n736 & n924));
  assign n3132 = (x0 | ~x2 | ~x4 | ~x5 | ~x6) & (~x0 | x2 | x4 | x5 | x6);
  assign z159 = n3134 | n3139 | ~n3147 | (~n542 & ~n3143);
  assign n3134 = ~x6 & (n3135 | ~n3138 | (~x5 & ~n3137));
  assign n3135 = x0 & ((~x5 & ~n3136) | (n1114 & n2007));
  assign n3136 = (x1 | x2 | ~x3 | x4 | ~x7) & (x7 | ((x1 | ~x2 | ~x3 | ~x4) & (~x1 | x3 | (~x2 ^ ~x4))));
  assign n3137 = (x3 | ~x7 | x1 | x2) & (x0 | ~x2 | (x1 ? ~x7 : (~x3 | x7)));
  assign n3138 = (~n2571 | ~n514) & (~n588 | ~n359 | ~n786);
  assign n3139 = x6 & (n3140 | (n789 & n588 & n514));
  assign n3140 = x5 & ((n387 & n3141) | (~x1 & ~n3142));
  assign n3141 = x2 & ~x7;
  assign n3142 = (~x0 | ((~x2 | ~x3 | ~x4 | ~x7) & (x2 | x3 | x7))) & (x4 | ((~x3 | ~x7 | x0 | ~x2) & (x2 | x3 | x7)));
  assign n3143 = ~n3144 & n3145 & (n868 | (~n306 & n1757));
  assign n3144 = ~x2 & ((x0 & x1 & x3 & ~x5) | (~x0 & ~x1 & x5));
  assign n3145 = ~n3146 & (n736 | ~n480 | ~n465);
  assign n3146 = x5 & ~x3 & x2 & ~x0 & ~x1;
  assign n3147 = ~n3148 & (n555 | n3149);
  assign n3148 = ~n565 & ~n1255 & (n2514 | (x0 & ~n1235));
  assign n3149 = x2 ? (x1 | (x0 & ~x3 & ~x4)) : (~x1 | (x3 & (~x0 | x4)));
  assign z160 = n3151 | n3154 | ~n3160 | (~x4 & ~n3156);
  assign n3151 = ~n878 & (n3153 | (~x1 & ~n3152));
  assign n3152 = (~x4 | ((x3 | x5 | x7) & (~x5 | ~x7 | x0 | ~x3))) & (~x5 | x7 | x3 | x4) & (~x0 | ((x4 | x5 | x7) & (x3 | (x7 & (x4 | x5)))));
  assign n3153 = x1 & ~x3 & (x0 ? ~x4 : ~x7);
  assign n3154 = x3 & ((~x0 & ~n2104) | (n744 & ~n3155));
  assign n3155 = (~x4 | x6 | x1 | ~x2) & (x2 | ((~x4 | ~x6) & (~x1 | x4 | x6)));
  assign n3156 = (~x2 | n3157) & (~x0 | x2 | ~n327 | n3159);
  assign n3157 = x0 ? (~n276 | ~n656) : (x7 | n3158);
  assign n3158 = (~x1 | ~x3 | ~x5 | x6) & (x1 | x3 | x5 | ~x6);
  assign n3159 = x1 ? (x3 | ~x7) : (~x3 | x7);
  assign n3160 = ~n3161 & ~n3163 & n3164 & (~n2847 | n3162);
  assign n3161 = ~n998 & ((~x1 & x3 & (x0 ^ ~x7)) | (~x0 & x7 & (x1 | ~x3)));
  assign n3162 = (x6 | ~x7 | x1 | ~x2) & (~x1 | x2 | (x6 ^ x7));
  assign n3163 = n740 & ((x3 & ~x7 & ~x0 & x1) | (x0 & x7 & (~x1 ^ x3)));
  assign n3164 = (~n300 | ~n2857) & (~x6 | n453 | ~n3165);
  assign n3165 = x4 & ~x2 & ~x0 & ~x1;
  assign z161 = ~n3170 | (~x4 & (n3169 | (x0 & ~n3167)));
  assign n3167 = (~x3 | ~x5 | ~n438 | n565) & (x3 | n3168);
  assign n3168 = (~x1 | x2 | ~x5 | ~x6 | ~x7) & (x1 | ((~x6 | ~x7 | x2 | x5) & (~x2 | ~x5 | x6 | x7)));
  assign n3169 = n387 & n501 & (x3 ? (~x6 ^ ~x7) : (~x6 & ~x7));
  assign n3170 = ~n3171 & n3176 & (x0 | (~n3174 & ~n3175));
  assign n3171 = x4 & (n3173 | (x5 & n441 & ~n3172));
  assign n3172 = (~x2 | x3 | (x6 ^ ~x7)) & (~x3 | (x2 ? (~x6 | ~x7) : (x6 | x7)));
  assign n3173 = n742 & n382 & n465;
  assign n3174 = x2 & ((n620 & n886) | (n276 & n629));
  assign n3175 = x4 & n408 & (x3 ? (~x5 ^ x7) : (~x5 ^ ~x7));
  assign n3176 = ~n3178 & n3179 & (~x2 | n3177);
  assign n3177 = (~x0 | ~x1 | x3 | x4 | x7) & (x0 | ((~x1 | x3 | x4 | ~x7) & (x1 | ~x3 | ~x4 | x7)));
  assign n3178 = ~n310 & ((x4 & (x1 ? (~x0 | n725) : x0)) | (~x0 & ~x4 & (~x1 | n725)));
  assign n3179 = x4 | ((n487 | ~n2569) & (~n363 | n3180));
  assign n3180 = x3 ? ((x5 | ~x7) & (x2 | ~x5 | x7)) : (x5 ^ x7);
  assign z162 = (x4 | ~n3182) & (n3190 | ~n3191 | ~x4 | n3188);
  assign n3182 = x3 ? (~n3186 & n3187) : n3183;
  assign n3183 = x1 ? n3184 : n3185;
  assign n3184 = (x2 | (x0 & (~x5 | ~x6 | ~x7))) & (~x0 | ~x2 | x5 | x6 | x7) & (x0 | (~x5 & ~x6 & ~x7));
  assign n3185 = (~x0 & x5 & (~x2 | x6)) | (~x6 & ~x7 & ~x2 & ~x5) | (x0 & ((x2 & (~x5 | (~x6 & ~x7))) | (~x5 & (~x6 | ~x7))));
  assign n3186 = x2 & ((x5 & x6 & x0 & ~x1) | (~x0 & (x1 ? (~x5 & x6) : (x5 & ~x6))));
  assign n3187 = (x1 & (x0 | (x2 & ~x5))) | (~x0 & ~x1 & x5 & ~n900) | (x0 & (x2 | ~x5));
  assign n3188 = ~n3189 & x3 & ~n878;
  assign n3189 = (~x0 | x1 | ~x5 | x7) & (x0 | (x1 ? (x5 | x7) : (~x5 | ~x7)));
  assign n3190 = x0 & (x1 ? ~x2 : (~x5 | (x2 & ~x6)));
  assign n3191 = (x0 | n3192) & (~x5 | n878 | ~n1706);
  assign n3192 = (~x1 | ~x2 | x5 | x6) & (x1 | x2 | ~x5 | ~x6);
  assign z163 = n3197 | ~n3204 | (x6 ? ~n3200 : ~n3194);
  assign n3194 = ~n3195 & (~n790 | ~n588 | ~n364);
  assign n3195 = ~x1 & ((n312 & n2007) | (n423 & ~n3196));
  assign n3196 = (x0 | ~x5 | ~x7) & (~x4 | ((~x5 | ~x7) & (~x0 | x5 | x7)));
  assign n3197 = ~x0 & (x3 ? ~n3199 : (n282 & n3198));
  assign n3198 = x4 & (~x5 ^ ~x6);
  assign n3199 = (~x1 | ~x2 | ~x5 | x6) & (x4 | ((x1 | x2 | ~x5 | ~x6) & (x5 | (~x1 ^ (x2 & ~x6)))));
  assign n3200 = x0 ? ((~n269 | ~n1183) & ~n3201) : n3202;
  assign n3201 = ~n570 & ((n725 & n606) | (n438 & n588));
  assign n3202 = (~n1658 | ~n1187) & (x4 | n3203);
  assign n3203 = (x1 | ~x2 | ~x3 | ~x5 | ~x7) & (~x1 | x7 | (x2 ? (~x3 | ~x5) : (x3 | x5)));
  assign n3204 = ~n3210 & ~n3209 & ~n3208 & ~n3205 & ~n3207;
  assign n3205 = ~n3206 & (x1 ? (~x5 ^ ~x7) : (~x5 & ~x7));
  assign n3206 = (x0 | ~x3 | ~x4 | (~x2 ^ ~x6)) & (x4 | x6 | ~x2 | x3);
  assign n3207 = ~n1417 & ((~x2 & (x3 ? (x4 & x6) : (~x4 & ~x6))) | (x2 & ~x3 & ~x4 & x6));
  assign n3208 = ~x1 & ((n340 & n764) | (n339 & n494));
  assign n3209 = ~n1230 & ((n438 & ~n379) | (~x2 & ~n1417));
  assign n3210 = n364 & n1687;
  assign z164 = n3212 | ~n3216 | n3225 | (~x6 & ~n3224);
  assign n3212 = ~x2 & (n3215 | (~x5 & (n3213 | n3214)));
  assign n3213 = x0 & ((n620 & n634) | (n276 & n633));
  assign n3214 = n601 & ((x1 & ~x3 & x6 & x7) | (x3 & ~x6 & (~x1 | x7)));
  assign n3215 = n285 & n2038 & (~x1 | x7);
  assign n3216 = n3219 & (n565 | (~n3217 & n3218));
  assign n3217 = n601 & ((n725 & n464) | (~x1 & ~n469));
  assign n3218 = x2 ? (x3 | x4 | (~x0 & ~x1)) : (~x3 | ~x4);
  assign n3219 = ~n3221 & n3223 & (~n663 | n3220);
  assign n3220 = (~x3 | x5 | ~x6 | x7) & (~x5 | ((x3 | ~x6 | ~x7) & (x1 | (x3 ? (x6 | x7) : ~x6))));
  assign n3221 = (n356 | n889) & (~x0 | n1837) & (x0 | n3222);
  assign n3222 = x2 & x6;
  assign n3223 = (~n295 | ~n635) & (~n1370 | (~n413 & ~n394));
  assign n3224 = (x4 | x7 | ~x0 | x2) & (x0 | ~x4 | (x2 ? (~x3 | x7) : x3));
  assign n3225 = x0 & ((n1658 & n634) | (x6 & ~n3226));
  assign n3226 = (~x1 | x2 | x3 | x4 | ~x7) & (x1 | ~x2 | (x3 ? x4 : (~x4 | x7)));
  assign z165 = n3228 | ~n3231 | (~n271 & ~n3230);
  assign n3228 = ~x2 & ((~x0 & x3 & n1863) | (~x3 & ~n3229));
  assign n3229 = x0 ? ((x5 | ~x7 | x1 | x4) & (~x1 | ~x4 | ~x5 | x7)) : (x4 | (x1 ? (x5 | ~x7) : (~x5 | x7)));
  assign n3230 = (~x0 | x4 | (~x3 ^ x7)) & (~x4 | ((x0 | x3 | x7) & (~x3 | ~x7)));
  assign n3231 = n3233 & ~n3235 & ~n3236 & (~x0 | n3232);
  assign n3232 = (~x1 | ~x2 | x3 | x4 | ~x7) & (x1 | ((x3 | ~x4 | x7) & (x2 | ~x3 | (x4 ^ x7))));
  assign n3233 = ~n3234 & ((~n408 & ~n282) | ~n329 | n487);
  assign n3234 = ~n566 & ~n506 & n408 & n760;
  assign n3235 = n663 & ((~x5 & ~n310) | (~x1 & x5 & ~n487));
  assign n3236 = x1 & (n3237 | (n424 & n782 & n1390));
  assign n3237 = ~n3238 & ~x7 & ~n1163;
  assign n3238 = (~x0 | x2 | ~x4 | x5) & (x0 | x4 | ~x5);
  assign z166 = ~n3242 | (~x2 & (x0 ? ~n3240 : ~n3241));
  assign n3240 = (x1 & ((x4 & x7) | (~x6 & ~x7 & ~x4 & ~x5))) | (~x1 & ((x6 & x7 & ~x4 & x5) | (x4 & ~x7))) | (x4 & (x7 ? (~x5 | ~x6) : (x5 | x6)));
  assign n3241 = x4 ? ((~x5 & (~x6 | ~x7)) | (x1 & (~x5 | (~x6 & ~x7)))) : ((x5 & (x6 | x7)) | (~x1 & (~x6 ^ x7)));
  assign n3242 = ~n1420 & (x4 | n3243) & (~x2 | n3246);
  assign n3243 = (~x2 | x3 | ~x5 | ~n480) & (x5 | n3244);
  assign n3244 = (~x2 | x3 | ~x6 | ~n480) & (x6 | n3245);
  assign n3245 = (x0 | x1 | x2 | ~x3 | x7) & (~x0 | ~x1 | x3 | (x2 ^ x7));
  assign n3246 = (x1 | (x0 ? x4 : (~x4 | ~x5))) & (x0 | (x4 ? (~x5 | ~x6) : (x5 & (~x1 | x6))));
  assign z167 = ~n3251 | (~x3 & (n3250 | (~x5 & ~n3248)));
  assign n3248 = (x6 | n3249) & (n847 | ~n363 | x4 | ~x6);
  assign n3249 = (~x0 | ~x1 | x2 | ~x4 | x7) & (x0 | ((~x1 | ~x2 | x4 | ~x7) & (~x4 | x7 | x1 | x2)));
  assign n3250 = n424 & n480 & (x2 ^ (~x6 & ~x7));
  assign n3251 = n3254 & (x2 ? (x3 ? n3252 : n3253) : (x3 ? n3253 : n3252));
  assign n3252 = (x0 | ((~x1 | (x5 ? (x6 | x7) : ~x6)) & (x5 | ~x6 | x7))) & (x1 | ((x0 | x5 | x6 | ~x7) & (~x0 | ~x5 | (x6 & x7))));
  assign n3253 = x0 ? ((x6 | x7 | ~x1 | x5) & (x1 | ~x5 | (x6 & x7))) : ((~x1 | (x5 ? (x6 | x7) : ~x6)) & (x5 | (x6 ? x7 : x1)));
  assign n3254 = n3257 & (~x7 | n3255) & (~n441 | n3256);
  assign n3255 = ((x2 ^ x5) | (x0 ? (x1 | ~x6) : (~x1 | x6))) & (~x0 | ~x1 | x2 | ~x5) & (x0 | x1 | ~x2 | x5 | ~x6);
  assign n3256 = (~x2 | ~x3 | x5 | x6 | x7) & (x2 | x3 | ~x5 | ~x6 | ~x7);
  assign n3257 = (~n364 | ~n556) & (~n424 | ~n717 | ~n1471);
  assign z168 = n3259 | n3262 | ~n3264 | (x2 & ~n3261);
  assign n3259 = x5 & ((n514 & n1586) | (n1752 & ~n3260));
  assign n3260 = (x0 | x2 | ~x3 | ~x4 | ~x7) & (~x0 | x3 | x4 | (~x2 ^ ~x7));
  assign n3261 = (x0 & (~x6 | (~x3 & ~x4))) | (x1 & x6) | (~x6 & (~x1 | (~x3 & ~x4)));
  assign n3262 = ~n3263 & (x1 ? (~x6 ^ x7) : (~x6 ^ ~x7));
  assign n3263 = (x0 & ~x2 & ~x3 & ~x4) | (x2 & (~x0 | x3 | x4));
  assign n3264 = n3265 & (n561 | ~n1064 | x7 | ~n328);
  assign n3265 = x3 | x4 | (x6 ? ~n364 : n3266);
  assign n3266 = (~x2 | x7 | x0 | ~x1) & (~x0 | x1 | x2 | ~x7);
  assign z169 = ~n3269 | ~n3275 | (n606 & ~n3268);
  assign n3268 = (x0 | ~x1 | ~x2 | ~x5 | ~x7) & (x1 | ((x2 | ~x5 | x7) & (~x0 | x5 | (~x2 ^ x7))));
  assign n3269 = ~n3270 & n3272 & (x7 | ~n465 | n3271);
  assign n3270 = n426 & ((n387 & n341) | (x0 & ~n3033));
  assign n3271 = (x0 | x1 | x2 | x4 | ~x6) & (~x0 | ~x1 | ~x2 | ~x4 | x6);
  assign n3272 = ~n3273 & ~n3274 & (~n359 | ~n3013);
  assign n3273 = x3 & ((x2 & x7 & ~x0 & x1) | (x0 & ~x1 & ~x2 & ~x7));
  assign n3274 = (~x0 | x3) & (x1 ? (~x2 & ~x7) : (x2 & x7));
  assign n3275 = ~n3277 & (x2 | n3276);
  assign n3276 = (x0 | x1 | ~x3 | x4 | x7) & (x3 | ((x1 | ~x4 | x7) & (~x0 | ((~x4 | x7) & (~x1 | x4 | ~x7)))));
  assign n3277 = ~n542 & ((n394 & n1458) | (~x0 & ~n670));
  assign z170 = ~n3281 | (x0 & (~n3280 | (~x1 & n3279)));
  assign n3279 = x2 & ~x4 & x5 & (x3 ^ x6);
  assign n3280 = x3 ? (x4 | (x1 ? x2 : x5)) : ((x2 | ~x4) & (x1 | (~x4 & (x2 | ~x5))));
  assign n3281 = n3283 & (x0 | (x3 & n2758) | (~x3 & n3282));
  assign n3282 = (x1 & x2 & ~x4 & ~x5 & ~x6) | (~x1 & ((x4 & x5 & x6) | (~x2 & (x4 ? x5 : (~x5 & ~x6)))));
  assign n3283 = ~n3284 & (x7 | (~n3210 & (n878 | n3285)));
  assign n3284 = n270 & n2076;
  assign n3285 = (~x0 | x1 | ~x3 | x4 | ~x5) & (x0 | ((~x4 | ~x5 | x1 | x3) & (~x1 | ~x3 | x4 | x5)));
  assign z171 = ~n3288 | ~n3294 | (~n409 & ~n3287);
  assign n3287 = (x1 | x4 | ~x5 | (~x2 ^ ~x6)) & (~x1 | x2 | ~x4 | x5 | x6);
  assign n3288 = n3289 & n3290 & n3291 & (n868 | n1249);
  assign n3289 = (x0 | ~x1 | x4 | ~x5) & (~x0 | ~x4 | (x1 ? (x2 | ~x5) : x5));
  assign n3290 = x0 | x1 | ~x2 | (~n335 & ~n512);
  assign n3291 = (~x1 | ~x2 | ~x6 | ~n3293) & (x2 | (x6 ? n3292 : ~n3293));
  assign n3292 = (~x0 | ~x1 | ~x4 | x5) & (x0 | x1 | (x4 ^ x5));
  assign n3293 = x7 & ~x5 & ~x0 & ~x4;
  assign n3294 = ~n3296 & (n878 | (~n3295 & (~n662 | ~n728)));
  assign n3295 = n1295 & ((~n436 & n744) | (n2773 & ~n1597));
  assign n3296 = n450 & ((n359 & n3297) | (x1 & ~n3298));
  assign n3297 = ~x6 & x3 & ~x4;
  assign n3298 = (x0 | ~x2 | ~x3 | ~x4 | ~x6) & (~x0 | x3 | x6 | (~x2 ^ x4));
  assign z172 = ~n3303 | (x1 & (~n3301 | (~n1291 & ~n3300)));
  assign n3300 = (x0 | ~x2 | ~x3 | x4 | ~x6) & (x6 | (x0 ? (x2 ? (x3 | x4) : (~x3 | ~x4)) : (x2 | (x3 ^ ~x4))));
  assign n3301 = (~n661 | ~n1514) & (~n329 | n3302);
  assign n3302 = (x2 | ~x3 | x5 | x6 | ~x7) & (~x2 | ~x6 | (x3 ? (x5 | ~x7) : (~x5 | x7)));
  assign n3303 = ~n3304 & ~n3307 & n3310 & (~x2 | n3309);
  assign n3304 = ~x1 & ((~x4 & ~n3306) | (~n570 & ~n3305));
  assign n3305 = x0 ? (~x3 | (x2 ? (~x4 | ~x6) : x6)) : (x3 | ~x4 | (~x2 ^ ~x6));
  assign n3306 = x0 ? (~x2 | n2811) : (n1424 | (x2 ^ x6));
  assign n3307 = x4 & (x5 ? (n380 & ~n878) : ~n3308);
  assign n3308 = x0 ? (x3 | (x1 ? (x2 | ~x6) : (~x2 | x6))) : (x1 | ~x3 | (x2 ^ x6));
  assign n3309 = (x0 | (x1 ? ((~x5 | x6) & (x3 | x5 | ~x6)) : (x5 | x6))) & (x1 | ((~x3 | x5 | x6) & (~x5 | ~x6 | ~x0 | x3)));
  assign n3310 = (x2 | n3311) & (x5 | ~n718 | n3312);
  assign n3311 = (~x5 & (~x1 | (x0 & ~x3 & x6))) | (x1 & x5) | (~x6 & (~x0 | x3));
  assign n3312 = (~x0 | (x2 ? (x3 | ~x6) : (~x3 | x6))) & (x0 | x2 | x3 | x6);
  assign z173 = n3314 | ~n3320 | (x6 & (n3318 | n3319));
  assign n3314 = ~x0 & (n3316 | (~n703 & ~n3315));
  assign n3315 = (~x6 | ~x7 | ~x3 | x5) & (~x2 | ((~x6 | ~x7 | x3 | ~x5) & (~x3 | x6 | x7)));
  assign n3316 = x2 & ((n1933 & n921) | (~n542 & ~n3317));
  assign n3317 = x1 ? (~x3 | x4) : (x3 | ~x4);
  assign n3318 = n473 & ((~x0 & ~x2 & x3 & x5) | (x2 & (x0 ? (~x3 ^ ~x5) : (~x3 & ~x5))));
  assign n3319 = ~n469 & x4 & n387;
  assign n3320 = n3323 & (n565 | (n3322 & (x5 | n3321)));
  assign n3321 = (x0 | x2 | ~x3 | (~x1 ^ ~x4)) & (~x0 | x1 | ~x2 | x3 | x4);
  assign n3322 = (~x1 | x4 | (x0 ? (~x2 | x3) : (x2 | ~x3))) & (x2 | (x1 & ~x4) | (~x0 ^ ~x3));
  assign n3323 = n3326 & (~x0 | (~n3325 & (n542 | n3324)));
  assign n3324 = (~x1 | x2 | x3 | x4 | x5) & (x1 | ~x2 | ~x3 | (~x4 & ~x5));
  assign n3325 = n606 & ((n725 & n921) | (n438 & n313));
  assign n3326 = x0 ? n3328 : n3327;
  assign n3327 = x1 ? (x3 | x4 | (~x2 ^ ~x6)) : (~x3 | ~x4 | (~x2 ^ x6));
  assign n3328 = (~x1 | x2 | ~x3 | x4 | x6) & (x3 | ((x2 | ~x4 | x6) & (x1 | (x2 ? (~x4 | ~x6) : x6))));
  assign z174 = ~n3334 | ~n3331 | (n441 & n1019 & ~n3330);
  assign n3330 = (x5 | ~x7 | x2 | ~x3) & (~x2 | ~x5 | (~x3 ^ ~x7));
  assign n3331 = x0 | (n3332 & (n703 | n3333));
  assign n3332 = (~x4 | ~x7 | x2 | x3) & (x1 | ((x2 | x3 | ~x7) & (~x2 | ~x3 | ~x4 | x7)));
  assign n3333 = (~x3 | (x2 ? (x5 | ~x7) : (~x5 | x7))) & (~x2 | x3 | (x5 ^ x7));
  assign n3334 = n3337 & (n565 | n3335) & (~n330 | n3336);
  assign n3335 = x4 ? (n605 | ~n380) : (~n1064 | n791);
  assign n3336 = (~x1 | x2 | x3 | x5 | ~x7) & (x1 | ~x2 | (x3 ? (x5 ^ x7) : (~x5 | x7)));
  assign n3337 = x3 ? ((~x7 | n3339) & (x2 | x7 | n3338)) : ((x7 | n3339) & (~x2 | ~x7 | n3338));
  assign n3338 = x0 ? (~x1 | x4) : (x1 | ~x4);
  assign n3339 = x0 ? ((x2 | ~x4) & (x1 | (x2 & ~x4))) : (~x1 | x4);
  assign z175 = ~n3343 | ~n3350 | (x0 & ~n3341);
  assign n3341 = (~x1 | x3 | x4 | n903) & (~x4 | ~n3342 | x1 | ~x3);
  assign n3342 = x6 & (x2 ^ ~x5);
  assign n3343 = ~n3344 & n3345 & n3346 & (~n363 | ~n2821);
  assign n3344 = ~x2 & (x1 ? (~x4 & (~x3 ^ x5)) : (x4 & x5));
  assign n3345 = (n605 | ~n2920 | n3317) & (~n282 | ~n1458);
  assign n3346 = (x2 | n3348) & (~n3347 | n3349);
  assign n3347 = x3 & (x2 ^ ~x5);
  assign n3348 = (x0 | ~x1 | x3 | x4 | ~x5) & (~x0 | x5 | (x1 ? (~x3 | x4) : (x3 | ~x4)));
  assign n3349 = (~x0 | x1 | ~x4 | x6 | ~x7) & (x0 | x4 | (x1 ? (x6 | ~x7) : (~x6 | x7)));
  assign n3350 = ~n3353 & (n703 | (~n3352 & (x3 | n3351)));
  assign n3351 = (~x0 | x2 | ~x5 | ~x6 | ~x7) & (~x2 | x5 | (x0 & (x6 | x7)));
  assign n3352 = ~x0 & x3 & ((x2 & (~x5 | ~x6)) | (~x5 & ~x6));
  assign n3353 = n426 & ((n313 & n1483) | (~x4 & ~n3354));
  assign n3354 = (x0 | ((x6 | x7 | x1 | ~x5) & (~x6 | ~x7 | ~x1 | x5))) & (x6 | ~x7 | ~x0 | x5);
  assign z176 = ~n3359 | (~n506 & ~n3358) | (~x4 & ~n3356);
  assign n3356 = (~n308 | ~n400 | ~n514) & (~n343 | n3357);
  assign n3357 = (~x1 | ((~x2 | x3 | ~x5) & (x2 | ~x3 | x5 | ~x7))) & (x3 | ((~x2 | ~x5 | x7) & (x1 | x2 | x5 | ~x7)));
  assign n3358 = (~x0 | ((x2 | ~x5) & (x1 | ~x2 | x5))) & (~x5 | ~x7 | ~x1 | x2) & (~x2 | ((x1 | x5 | ~x7) & (x0 | (x1 ? x5 : (~x5 | x7)))));
  assign n3359 = ~n3360 & n3363 & n3367 & (x1 | n3362);
  assign n3360 = ~n605 & ((n1063 & n1370) | (~x6 & ~n3361));
  assign n3361 = x0 ? ((~x1 | x3 | x4 | ~x7) & (x1 | ~x3 | ~x4 | x7)) : (~x4 | ~x7 | (x1 ^ x3));
  assign n3362 = (~x0 | ~x2 | ~x3 | x5 | x6) & (x0 | x2 | (x3 ? (x5 | x6) : (~x5 | ~x6)));
  assign n3363 = n3364 & ~n3365 & (~n425 | ~n285 | n3366);
  assign n3364 = (~n295 | ~n2431) & (n420 | n753);
  assign n3365 = ~n761 & ((n363 & n786) | (n387 & n450));
  assign n3366 = (~x1 | ~x2 | ~x6 | ~x7) & (x1 | x2 | x6 | x7);
  assign n3367 = ~n3369 & (x7 | (~n3368 & (~n1064 | n3192)));
  assign n3368 = n659 & ((n587 & n408) | (n282 & n1039));
  assign n3369 = ~n3370 & ((n601 & ~n506) | (n1964 & n1064));
  assign n3370 = (~x1 | x2 | ~x5 | x7) & (x1 | (x2 ? (x5 | x7) : (~x5 | ~x7)));
  assign z177 = ~n3376 | (~x3 & (x1 ? ~n3374 : ~n3372));
  assign n3372 = (x2 | n3373) & (~x0 | ~x2 | ~x4 | n565);
  assign n3373 = (~x0 | ~x4 | x5 | x6 | ~x7) & (x4 | (x0 ? ((~x5 | x6 | ~x7) & (~x6 | x7)) : (x5 ? (x6 | x7) : (~x6 | ~x7))));
  assign n3374 = x4 ? n3375 : (~n782 | ~n962);
  assign n3375 = x0 ? (x7 | (x2 ? (x5 | x6) : (~x5 | ~x6))) : (~x6 | ~x7 | (x2 ^ x5));
  assign n3376 = n3381 & (~x3 | (~n3377 & (~n725 | n3380)));
  assign n3377 = ~x1 & ((x4 & ~n3378) | (n601 & ~n3379));
  assign n3378 = x0 ? ((x6 | x7 | x2 | ~x5) & (~x6 | ~x7 | ~x2 | x5)) : (~x2 | ((x6 | ~x7) & (x5 | ~x6 | x7)));
  assign n3379 = (~x5 | ~x6 | x7) & (x2 | (x6 ^ ~x7));
  assign n3380 = (x4 | ((~x0 | ((x6 | ~x7) & (x5 | ~x6 | x7))) & (x6 | x7 | x0 | x5))) & (x0 | ~x4 | ~x5 | (~x6 ^ x7));
  assign n3381 = ~n3382 & n3386 & n3388 & (x0 | n3385);
  assign n3382 = ~n542 & (x1 ? ~n3383 : ~n3384);
  assign n3383 = (~x3 | x4 | x0 | ~x2) & (x3 | ((x0 | x2 | ~x4 | ~x5) & (~x0 | x4 | (~x2 & x5))));
  assign n3384 = (~x0 | ~x2 | ~x3 | ~x4 | ~x5) & ((~x4 ^ x5) | (x0 ? (x2 | ~x3) : (~x2 | x3)));
  assign n3385 = x1 ? (n614 | n761) : (~n273 | ~n426);
  assign n3386 = (n506 | n3387) & (~n428 | ~n590);
  assign n3387 = (x0 | x1 | x2 | ~x4) & (~x0 | (x1 ? (x2 | ~x4) : (~x2 | x4)));
  assign n3388 = (n506 | n3390) & (x0 | n3389);
  assign n3389 = (x1 | ~x2 | ~x3 | x4 | x6) & (~x1 | ((x4 | ~x6 | x2 | x3) & (~x2 | ~x3 | ~x4 | x6)));
  assign n3390 = (x0 | x1 | ~x2 | ~x4 | ~x5) & (~x0 | x2 | x4 | (~x1 ^ ~x5));
  assign z178 = ~n3399 | ~n3404 | (x0 ? ~n3396 : ~n3392);
  assign n3392 = ~n3393 & (~x5 | ~n278 | n3395);
  assign n3393 = ~x4 & (x7 ? (n1295 & ~n800) : ~n3394);
  assign n3394 = (x1 | ~x6 | (x2 ? (~x3 | ~x5) : (x3 | x5))) & (x6 | ((x1 | x2 | x3 | ~x5) & (~x1 | (x2 ? (x3 | ~x5) : (~x3 | x5)))));
  assign n3395 = (x1 | ~x3 | ~x6 | ~x7) & (~x1 | x3 | (x6 ^ ~x7));
  assign n3396 = ~n3398 & (x1 | ((~n1453 | ~n875) & ~n3397));
  assign n3397 = ~x5 & ((n340 & n622) | (~n350 & ~n800));
  assign n3398 = n411 & n1127;
  assign n3399 = ~n3400 & ~n3402 & (~x3 | n3403);
  assign n3400 = ~n566 & ((n345 & n1114) | (~x2 & ~n3401));
  assign n3401 = (x1 | ~x3 | ~x4 | x6 | x7) & (~x1 | ~x6 | (x3 ? (x4 | ~x7) : (~x4 | x7)));
  assign n3402 = ~n1016 & (n1734 | (~x0 & ~n384));
  assign n3403 = (~x7 | (x0 ? (x1 ? (x2 | ~x4) : (~x2 | x4)) : (~x4 | (x1 ^ x2)))) & (x2 | x4 | x7 | (~x0 ^ ~x1));
  assign n3404 = x1 ? n3407 : (~n3405 & (~x0 | n3406));
  assign n3405 = ~n315 & ((x3 & ~x4 & ~x5 & x7) | (~x3 & (x4 ? (~x5 ^ x7) : (x5 & ~x7))));
  assign n3406 = x2 ? ((x5 | ~x7 | x3 | x4) & (~x3 | ~x4 | ~x5 | x7)) : (~x3 | x7 | (x4 ^ ~x5));
  assign n3407 = x3 ? (~n579 | n3408) : n3409;
  assign n3408 = x4 ? (x5 ^ ~x7) : (~x5 | ~x7);
  assign n3409 = (x0 | x2 | ~x4 | ~x5 | x7) & ((x0 ^ ~x2) | (x4 ? (x5 | ~x7) : (x5 ^ x7)));
  assign z179 = ~n3420 | (x0 ? (n3411 | n3413) : ~n3415);
  assign n3411 = ~x2 & ((~n2723 & n3013) | (x7 & ~n3412));
  assign n3412 = x1 ? (~x5 | (x3 ? (x4 | ~x6) : (~x4 | x6))) : (x3 | x5 | (x4 ^ x6));
  assign n3413 = x2 & (x1 ? (n606 & n921) : ~n3414);
  assign n3414 = (~x3 | ~x4 | ~x5 | ~x6 | x7) & (x4 | (x3 ? (x6 | (~x5 ^ x7)) : (~x6 | (x5 ^ x7))));
  assign n3415 = x5 ? n3417 : (x1 ? n893 : n3416);
  assign n3416 = (x2 | ~x4 | (x3 ? (x6 | ~x7) : (~x6 | x7))) & (x4 | ((x2 | x3 | x6 | ~x7) & (~x2 | (x3 ? (x6 | x7) : (~x6 | ~x7)))));
  assign n3417 = x2 ? n3418 : (x7 | n3419);
  assign n3418 = x1 ? (x6 | (x3 ? (~x4 | x7) : (x4 | ~x7))) : (~x6 | (x3 ? (~x4 | ~x7) : (x4 | x7)));
  assign n3419 = (x1 | ~x3 | x4 | x6) & (~x1 | (x3 ? (x4 | ~x6) : (~x4 | x6)));
  assign n3420 = n3422 & n3426 & (~x1 | n3421);
  assign n3421 = (x0 | ~x2 | x3 | ~x5 | ~x6) & (x2 | ((x0 | x3 | x5 | ~x6) & (~x0 | (x3 ? (x5 | x6) : (~x5 | ~x6)))));
  assign n3422 = ~n3424 & ~n3425 & (~x5 | ~n659 | n3423);
  assign n3423 = (~x1 | x2 | ~x4 | ~x6) & (x1 | (x2 ? (x4 | ~x6) : (~x4 | x6)));
  assign n3424 = ~n1091 & ((x3 & ~x6 & ~x0 & x1) | (x0 & ~x1 & (~x3 ^ x6)));
  assign n3425 = n441 & ((n423 & n587) | (n1039 & n426));
  assign n3426 = (n1011 | n3427) & (x3 | (~n2763 & ~n3428));
  assign n3427 = (x0 | ~x1 | x5 | (x3 ^ x6)) & (x1 | (x0 ? (x3 ? (~x5 | x6) : (x5 | ~x6)) : (x3 ? (x5 | x6) : (~x5 | ~x6))));
  assign n3428 = ~x2 & ((n441 & n764) | (n981 & ~n770));
  assign z180 = n3434 | ~n3437 | ~n3444 | (x1 & ~n3430);
  assign n3430 = ~n3433 & (x2 | (x3 & n3432) | (~x3 & n3431));
  assign n3431 = (x0 | ~x4 | ~x5 | ~x6 | ~x7) & (x5 | x6 | x7 | (~x0 & x4));
  assign n3432 = (~x6 | ~x7 | x4 | ~x5) & (x0 | ~x4 | x5 | x6 | x7);
  assign n3433 = n720 & n1755;
  assign n3434 = ~n542 & ((n276 & ~n3436) | (x3 & ~n3435));
  assign n3435 = (~x4 | ~x5 | x1 | ~x2) & (~x1 | x5 | (x0 ? (x2 | ~x4) : (~x2 | x4)));
  assign n3436 = (~x2 | x4 | ~x5) & (x0 | x2 | ~x4 | x5);
  assign n3437 = n3441 & (~x2 | (~n3439 & (x3 | n3438)));
  assign n3438 = (~x4 | ~x6 | x0 | ~x1) & (~x0 | x6 | (x1 ? (x4 | x5) : (~x4 | ~x5)));
  assign n3439 = n659 & ((n327 & n473) | (n3440 & ~n614));
  assign n3440 = x1 & ~x6;
  assign n3441 = ~n3443 & (~n359 | ~n2077) & (x1 | n3442);
  assign n3442 = (x2 | x4 | (x3 ? (x5 | x6) : (~x5 | ~x6))) & (~x4 | ((~x2 | x5 | (~x3 ^ ~x6)) & (~x5 | ~x6 | x2 | ~x3)));
  assign n3443 = n725 & (n1161 | (x3 & ~n2519));
  assign n3444 = (n565 | n3446) & (x1 | (n3448 & (n565 | n3445)));
  assign n3445 = (x0 | ~x2 | (x3 ? (x4 | x5) : (~x4 | ~x5))) & (x2 | ~x3 | ((x4 | ~x5) & (~x0 | ~x4 | x5)));
  assign n3446 = n3447 & (n1896 | (x1 ? (~x2 | ~x5) : (x2 | x5)));
  assign n3447 = (~x0 | x1 | ~x2 | ~x3 | x4) & (~x1 | x3 | ((x2 | ~x4) & (x0 | ~x2 | x4)));
  assign n3448 = x0 ? n3449 : ((~n313 | ~n1453) & ~n3451);
  assign n3449 = x4 ? (~n339 | n1308) : n3450;
  assign n3450 = (~x6 | ~x7 | x3 | x5) & (~x3 | ~x5 | (x2 ? (~x6 | ~x7) : (x6 | x7)));
  assign n3451 = ~x3 & ((n1207 & n921) | (x2 & ~n585));
  assign z181 = ~n3455 | (x2 & ((n728 & n1755) | n3453));
  assign n3453 = ~x1 & ((~x4 & ~n3454) | (n921 & n1589));
  assign n3454 = (x6 | x7 | x3 | x5) & (~x3 | ~x5 | (x0 ? (x6 | ~x7) : (~x6 | x7)));
  assign n3455 = ~n3460 & n3465 & (x2 ? n3463 : n3456);
  assign n3456 = x7 ? n3459 : (~n3458 & (~x1 | n3457));
  assign n3457 = (x3 | ((x5 | x6 | ~x0 | ~x4) & (x0 | ~x6 | (x4 ^ x5)))) & (~x0 | ~x3 | ~x5 | (x4 ^ x6));
  assign n3458 = x6 & n276 & ((~x4 & ~x5) | (~x0 & x4 & x5));
  assign n3459 = x0 ? (~x3 | ~n494) : (x1 ? (~x3 | ~n764) : (x3 | ~n494));
  assign n3460 = ~n878 & (x0 ? ~n3462 : ~n3461);
  assign n3461 = (~x1 | x4 | (x3 ? (~x5 | x7) : (x5 | ~x7))) & (~x4 | ~x7 | ((x3 | ~x5) & (x1 | ~x3 | x5)));
  assign n3462 = (x5 | ~x7 | x3 | x4) & (x1 | ((~x3 | x4 | ~x5 | x7) & (x3 | ~x4 | (x5 ^ x7))));
  assign n3463 = (~n1183 | ~n1008) & (x3 | n3464);
  assign n3464 = (x0 | ~x1 | ~x4 | ~x5 | x7) & (x1 | ((~x0 | ~x5 | (~x4 ^ x7)) & (x0 | x4 | x5 | ~x7)));
  assign n3465 = n3468 & (n570 | n3467) & (x0 | n3466);
  assign n3466 = x3 ? ((~x5 | x7 | x2 | ~x4) & (x5 | ~x7 | ~x2 | x4)) : (x2 ? (x4 ? (x5 | x7) : (~x5 | ~x7)) : (x4 ? (x5 | ~x7) : (~x5 | x7)));
  assign n3467 = (~x0 | ~x1 | ~x2 | x3 | x4) & (~x3 | ((x1 | ~x2 | ~x4) & (x0 | (x2 ^ x4))));
  assign n3468 = ~n647 | (n3469 & (~n284 | n3159));
  assign n3469 = x4 ? (x5 | ~x7) : (x7 | (x3 ^ ~x5));
  assign z182 = ~n3482 | (x1 ? ~n3471 : ~n3476);
  assign n3471 = x5 ? n3474 : (~n3473 & (x2 | n3472));
  assign n3472 = (~x0 | x4 | ~x6 | (~x3 ^ ~x7)) & (~x4 | (x0 ? (x6 | (~x3 ^ ~x7)) : (~x6 | (~x3 ^ x7))));
  assign n3473 = ~n836 & n324 & ~x3 & ~x7;
  assign n3474 = (~n634 | ~n713) & (x0 | n3475);
  assign n3475 = x3 ? (x4 ? (~x6 | ~x7) : (x6 | x7)) : ((x4 | x6 | ~x7) & (~x6 | x7 | ~x2 | ~x4));
  assign n3476 = x3 ? n3477 : (x0 ? n3481 : n3480);
  assign n3477 = x5 ? n3478 : n3479;
  assign n3478 = (~x0 | x2 | ~x4 | ~x6 | ~x7) & (x0 | ~x2 | x4 | x6 | x7);
  assign n3479 = (~x6 | x7 | x0 | ~x4) & (~x7 | (x0 ? ((~x4 | x6) & (~x2 | x4 | ~x6)) : (x4 | x6)));
  assign n3480 = (~x6 | ~x7 | ~x4 | x5) & (x4 | ((~x6 | x7 | x2 | ~x5) & (~x2 | x6 | (x5 ^ x7))));
  assign n3481 = (~x4 | x7 | (x5 ^ x6)) & (x2 | x4 | ~x5 | x6 | ~x7);
  assign n3482 = n3485 & (n331 | n3484) & (~n367 | n3483);
  assign n3483 = (x1 | x2 | x3 | x4 | ~x5) & (~x1 | ~x4 | ((~x3 | x5) & (~x2 | x3 | ~x5)));
  assign n3484 = (x3 | ~x4 | ~x5 | x6) & (~x3 | ((x0 | x4 | x5 | ~x6) & (~x0 | (x4 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n3485 = ~n3486 & (~x6 | (~n3487 & (~x0 | ~n1465)));
  assign n3486 = ~n379 & ((n441 & n588) | (n606 & ~n3082));
  assign n3487 = n782 & ((n424 & n276) | (x1 & n400));
  assign z183 = ~n3500 | (x1 ? (n3495 | ~n3497) : ~n3489);
  assign n3489 = x3 ? (x5 ? n3490 : n3491) : n3492;
  assign n3490 = (~x0 | x4 | (x6 ^ x7)) & (~x2 | ((~x6 | x7 | ~x0 | ~x4) & (x0 | (x4 ? (x6 | ~x7) : (~x6 | x7)))));
  assign n3491 = (~x6 | x7 | x0 | ~x4) & (x2 | ((x6 | x7 | x0 | x4) & (~x0 | ~x4 | (x6 ^ x7))));
  assign n3492 = ~n3493 & ~n3494 & (~x0 | ~n278 | ~n556);
  assign n3493 = n484 & ((x6 & ~x7 & ~x0 & x4) | (x7 & (x0 ? (~x4 ^ x6) : (~x4 & x6))));
  assign n3494 = ~n614 & ((n382 & n647) | (x2 & ~n389));
  assign n3495 = ~n3496 & x6 & n285;
  assign n3496 = (~x2 | ~x4 | x5 | ~x7) & (x2 | x7 | (x4 ^ ~x5));
  assign n3497 = (n1254 | n3499) & (n677 | n3498);
  assign n3498 = (~x0 | x2 | ~x3 | ~x6 | x7) & (x0 | x6 | (x2 & x3) | ~x7);
  assign n3499 = (x0 | ~x2 | ~x3 | x5 | ~x7) & (~x0 | x2 | x3 | ~x5 | x7);
  assign n3500 = n3503 & (n836 | (~n3502 & (~x5 | n3501)));
  assign n3501 = (~x0 | x1 | x2 | x3 | ~x7) & (x0 | ((~x1 | ~x2 | ~x3 | ~x7) & (x1 | x2 | x7)));
  assign n3502 = ~x7 & n1921 & (n1658 | n625);
  assign n3503 = n3506 & (x1 ? n3505 : n3504);
  assign n3504 = x0 ? ((~x2 | x4 | x6 | ~x7) & (x2 | ~x4 | ~x6 | x7)) : ((x2 | ~x4 | x6 | ~x7) & (~x2 | x4 | (x6 ^ x7)));
  assign n3505 = (x2 | ~x7 | (x0 ? (x4 ^ x6) : (x4 | ~x6))) & (x0 | x7 | ((~x2 | ~x4 | ~x6) & (x4 | x6)));
  assign n3506 = (n444 | n3507) & (~n438 | ~n341 | n1581);
  assign n3507 = (x1 | x2 | ~x3 | x4 | ~x7) & (~x1 | ((~x2 | x3 | x4 | ~x7) & (x2 | ~x3 | ~x4 | x7)));
  assign z184 = n3511 | ~n3516 | (~n1291 & ~n3509);
  assign n3509 = x2 ? (n3510 & (~n387 | n506)) : n435;
  assign n3510 = (~x0 | x1 | x3 | x4 | ~x6) & (x0 | ((~x1 | (x3 ? (x4 | x6) : (~x4 | ~x6))) & (x1 | ~x3 | ~x4 | x6)));
  assign n3511 = ~n570 & (~n3513 | (x0 & ~n3512));
  assign n3512 = (x1 | ~x2 | ~x3 | ~x4 | ~x6) & (~x1 | x4 | (x2 ? (x3 | ~x6) : (~x3 | x6)));
  assign n3513 = ~n3514 & (~n438 | n444) & (~n1706 | n3515);
  assign n3514 = ~x2 & (x1 ? ((~x3 & x6) | (x0 & (~x3 | x6))) : (x3 & (~x0 | ~x6)));
  assign n3515 = x2 ? (x4 | x6) : ~x4;
  assign n3516 = ~n3519 & ~n3523 & (x0 ? n3517 : n3521);
  assign n3517 = (x6 | n3518) & (~n438 | n1597 | x5 | ~x6);
  assign n3518 = (x1 | x2 | x3 | x5) & (~x1 | ~x5 | (x2 ? (x3 | x4) : (~x3 | ~x4)));
  assign n3519 = x3 & ((n514 & n2837) | (x0 & ~n3520));
  assign n3520 = (x1 | ~x2 | ~x4 | ~n313) & (~x1 | x2 | x4 | ~n921);
  assign n3521 = (~n269 | ~n273) & (~x5 | n3522);
  assign n3522 = (~x1 | x2 | ~x3 | ~x6) & (x1 | ~x2 | x6 | (x3 ^ ~x4));
  assign n3523 = n285 & ((n424 & ~n3524) | (n932 & n313));
  assign n3524 = (~x1 | ~x2 | ~x6 | x7) & (x1 | x6 | (~x2 ^ x7));
  assign z185 = n3526 | ~n3529 | n3534 | (~n542 & ~n3532);
  assign n3526 = x6 & ((n285 & ~n3528) | (x3 & ~n3527));
  assign n3527 = (x0 | ~x1 | ~x2 | ~x4 | x5) & (~x0 | ((~x4 | ~x5 | x1 | ~x2) & (x4 | x5 | ~x1 | x2)));
  assign n3528 = (~x1 | ~x2 | x4 | ~x5) & (x1 | (x2 ? (x4 | x5) : (~x4 | ~x5)));
  assign n3529 = (~x0 | n3531) & (~n410 | ~n411) & (x0 | n3530);
  assign n3530 = (~x3 | ((x1 | (x2 ? (~x4 | x6) : ~x6)) & (~x1 | ~x2 | x4 | ~x6))) & (~x1 | x3 | (x2 ? (~x4 | ~x6) : x6));
  assign n3531 = (~x1 | x2 | x3 | ~x6) & (x1 | x6 | (x2 ? (x3 | x4) : ~x3));
  assign n3532 = ~n1965 & (~x0 | ~n567) & (~x5 | n3533);
  assign n3533 = (x0 | ~x2 | (x1 ? (~x3 | ~x4) : (x3 | x4))) & (~x0 | ~x1 | x2 | ~x3 | x4);
  assign n3534 = ~n565 & (~n3536 | (~x5 & ~n3535));
  assign n3535 = (~x0 | x1 | ~x2 | ~x3 | ~x4) & (x0 | x3 | (x1 ? (~x2 | x4) : (x2 | ~x4)));
  assign n3536 = (x2 | ~x3 | x0 | ~x1) & (x1 | ((~x0 | ~x2 | (~x3 ^ x4)) & (x3 | x4 | x0 | x2)));
  assign z186 = n3538 | ~n3543 | ~n3544 | (x2 & ~n3542);
  assign n3538 = ~x6 & (n3540 | (~n1486 & ~n3539));
  assign n3539 = (x0 | ~x4 | (x2 ? (~x3 | x5) : (x3 | ~x5))) & (~x0 | x2 | ~x3 | x4 | x5);
  assign n3540 = x2 & ((~x3 & ~n3541) | (n1555 & n1008));
  assign n3541 = x0 ? ((~x5 | ~x7 | x1 | x4) & (~x1 | ~x4 | x5 | x7)) : (x4 | (x1 ? (~x5 | x7) : (x5 | ~x7)));
  assign n3542 = (~x0 | ~x1 | x3 | x4 | x7) & (x0 | x1 | ~x3 | ~x4 | ~x7) & ((x3 ^ ~x4) | ((x1 | x7) & (x0 | ~x1 | ~x7)));
  assign n3543 = (~n2076 | ~n1514) & (~x4 | ~n387 | n1699);
  assign n3544 = ~n3545 & (n570 | n3535) & (x2 | n3548);
  assign n3545 = ~x4 & (n3547 | (x0 & ~n3546));
  assign n3546 = (~x1 | x2 | ~x3 | ~x5 | x7) & (x1 | ~x2 | x3 | x5 | ~x7);
  assign n3547 = ~x7 & x5 & ~x3 & ~x0 & ~x1;
  assign n3548 = x3 ? (x1 ? (x7 | (x0 & ~x4)) : ~x7) : ((~x0 | (~x1 ^ ~x7)) & (~x1 | x4 | ~x7));
  assign z187 = ~n3554 | (x7 & (x1 ? ~n3552 : ~n3550));
  assign n3550 = (~n1837 | n3551) & (~x2 | n580 | n566);
  assign n3551 = (~x0 | ~x3 | x4 | x5) & (x0 | x3 | (x4 ^ x5));
  assign n3552 = (~n273 | ~n713) & (x0 | n3553);
  assign n3553 = (x2 | x3 | ~x4 | ~x5 | ~x6) & (~x2 | ((~x3 | ~x4 | x5 | ~x6) & (~x5 | x6 | x3 | x4)));
  assign n3554 = ~n3555 & ~n3558 & n3559 & (n566 | n3557);
  assign n3555 = ~x3 & (x0 ? (~x1 & n278) : ~n3556);
  assign n3556 = x1 ? ((~x2 | ~x4 | ~x5 | ~x6) & (x5 | x6 | x2 | x4)) : (~x5 | (x2 ? (x4 | x6) : (~x4 | ~x6)));
  assign n3557 = (x1 | ~x2 | ~x3 | ~x4 | ~x6) & (~x1 | x2 | (x3 ? (~x4 | x6) : (x4 | ~x6)));
  assign n3558 = n314 & (x0 ? (~x2 & n1019) : (x2 & ~n836));
  assign n3559 = n3560 & (~n443 | n998 | x5 | ~n363);
  assign n3560 = (x0 | ~x2 | ~x4 | (x3 ^ x5)) & (x2 | ((~x3 | x4 | (x0 & ~x5)) & (~x0 | x5 | (x3 ^ x4))));
  assign z188 = ~n3563 | ~n3569 | ~n3573 | (~x2 & ~n3562);
  assign n3562 = (x0 | ~x1 | ~x3 | ~x4 | ~x5) & (x1 | ((x0 | x3 | x4 | ~x5) & (~x4 | (x0 ? (x3 ^ x5) : (~x3 | x5)))));
  assign n3563 = n3564 & (n2723 | n3567) & (~n1122 | n3568);
  assign n3564 = (n485 | n3566) & (n677 | n3565);
  assign n3565 = x0 ? ((~x3 | ~x6 | x1 | ~x2) & (x3 | x6 | ~x1 | x2)) : (x1 | x2 | (~x3 ^ x6));
  assign n3566 = (~x0 | ((x1 | ~x2 | x3 | ~x5) & (~x1 | x2 | ~x3 | x5))) & (x0 | x1 | ~x2 | x3 | x5);
  assign n3567 = (~n661 | ~n662) & (~x7 | ~n329 | n2212);
  assign n3568 = (x2 | x4 | (x5 ? (~x6 | x7) : (x6 | ~x7))) & (~x2 | ~x4 | ~x5 | x6 | ~x7);
  assign n3569 = x1 ? (x2 ? n3572 : n3571) : (n3570 & (~x2 | n3571));
  assign n3570 = (~n312 | ~n458) & (n510 | (~n2431 & ~n2560));
  assign n3571 = x0 ? (x3 ? (x4 | ~x5) : (~x4 | x5)) : (x4 | (~x3 ^ x5));
  assign n3572 = (~x0 | x3 | x4 | x5) & (x0 | ~x3 | (x4 ^ x5));
  assign n3573 = ~n3574 & (x0 | ((~n1127 | ~n1145) & ~n3576));
  assign n3574 = x1 & (x0 ? (n423 & n301) : ~n3575);
  assign n3575 = (~x4 | x5 | ((x3 | x6) & (x2 | ~x3 | ~x6))) & (~x2 | x4 | ~x5 | (~x3 ^ x6));
  assign n3576 = ~x7 & (n3577 | (x6 & n923 & ~n2933));
  assign n3577 = x1 & ((n426 & n971) | (n423 & n512));
  assign z189 = ~n3595 | ~n3589 | n3579 | n3583;
  assign n3579 = ~x2 & (n3580 | (n1921 & ~n3582));
  assign n3580 = x5 & (x0 ? (n923 & n622) : ~n3581);
  assign n3581 = x1 ? (~x6 | (x3 ? (x4 | x7) : (~x4 | ~x7))) : (x6 | ((x4 | x7) & (x3 | ~x4 | ~x7)));
  assign n3582 = (x1 | x3 | x4 | x6 | ~x7) & (~x1 | ~x3 | (x4 ? (x6 | ~x7) : (x6 ^ x7)));
  assign n3583 = ~x2 & (n3585 | ~n3586 | (x0 & ~n3584));
  assign n3584 = (x1 | x3 | x4 | x5 | ~x6) & (~x4 | ((x1 | ~x3 | ~x5 | x6) & (~x1 | (x3 ? (~x5 | ~x6) : (x5 | x6)))));
  assign n3585 = ~n467 & ((x0 & ~x1 & (~x4 ^ ~x6)) | (x1 & (x0 ? (x4 & x6) : (~x4 & ~x6))));
  assign n3586 = ~n3587 & ~n3588 & (~n273 | ~n765);
  assign n3587 = ~x0 & ~x1 & x4 & (~x5 ^ x6);
  assign n3588 = x1 & ((x5 & ~x6 & x0 & ~x4) | (~x5 & x6 & ~x0 & x4));
  assign n3589 = ~n3591 & (n379 | (x0 & n3594) | (~x0 & n3590));
  assign n3590 = (x1 | ~x2 | ~x3 | ~x4 | ~x7) & (~x1 | x2 | x3 | x4 | x7);
  assign n3591 = x2 & (~n3592 | ~n3593 | (~n379 & ~n755));
  assign n3592 = (~n273 | ~n363) & (~n457 | ~n512);
  assign n3593 = x6 ? (n467 | ~n507) : (~n730 | n703);
  assign n3594 = (~x1 | ~x2 | x3 | x4 | x7) & (x1 | x2 | (x3 ? (x4 | ~x7) : (~x4 | x7)));
  assign n3595 = ~n3597 & (~x2 | (n3600 & (~n3596 | n3599)));
  assign n3596 = ~x1 & ~x6;
  assign n3597 = ~n688 & ((n300 & n1314) | (~x2 & ~n3598));
  assign n3598 = (x0 | ~x3 | (x1 ? (~x5 | x6) : (x5 | ~x6))) & (~x0 | ~x1 | x3 | x5 | ~x6);
  assign n3599 = (~x5 | ~x7 | ~x0 | ~x4) & (x0 | x5 | (x3 ? (x4 | x7) : (~x4 | ~x7)));
  assign n3600 = ~n3602 & (~n1514 | ~n1177) & (n542 | n3601);
  assign n3601 = (~x0 | x1 | x3 | x4 | ~x5) & (x0 | ~x1 | ~x3 | ~x4 | x5);
  assign n3602 = ~n534 & ((n363 & n2220) | (n387 & n403));
  assign z190 = n2377 | ~n2382 | (x2 ? ~n3604 : ~n2372);
  assign n3604 = ~n2368 & (~n367 | n3605);
  assign n3605 = (x1 | x3 | x5 | ~x7) & (~x3 | ((x4 | x5 | ~x7) & (~x1 | ((x5 | ~x7) & (~x4 | ~x5 | x7)))));
  assign z191 = ~n2387 | ~n3610 | (n3607 & (n3608 | n3609));
  assign n3607 = ~x3 & ~x7;
  assign n3608 = n1921 & (x1 ? (x4 & ~x6) : (x2 ? (~x4 ^ x6) : (~x4 & x6)));
  assign n3609 = n730 & ((x1 & ~x2 & x4 & ~x6) | (~x1 & (x2 ? (~x4 ^ x6) : (~x4 & x6))));
  assign n3610 = ~n3611 & ~n3614 & (~n923 | ~n2404);
  assign n3611 = ~n542 & (~n3613 | (~x0 & ~n3612));
  assign n3612 = x1 ? (x3 | (x2 ? (~x4 | ~x5) : (~x4 ^ x5))) : ((~x4 | ~x5 | x2 | ~x3) & (x4 | x5 | ~x2 | x3));
  assign n3613 = (x0 | ~x1 | ~x2 | ~x3 | x4) & (~x0 | x2 | (x1 ? (x3 | x4) : (~x3 | ~x4)));
  assign n3614 = ~n565 & (x1 ? ~n2401 : ~n3615);
  assign n3615 = (x3 | ((x2 | ~x4 | (x0 & x5)) & (~x0 | ~x5 | (~x2 ^ ~x4)))) & (~x2 | ~x3 | x4 | (x0 & x5));
  assign z192 = n3620 | ~n3622 | (x3 ? ~n3617 : ~n3619);
  assign n3617 = (~x0 | ~x5 | n2407) & (x0 | ~x4 | x5 | n3618);
  assign n3618 = (~x1 | x2 | ~x6 | x7) & (x1 | (x2 ? (x6 ^ x7) : (x6 | ~x7)));
  assign n3619 = (n1974 | n2411) & (~n387 | ~n3222 | n1435);
  assign n3620 = ~x7 & (x3 ? (n335 & n394) : ~n3621);
  assign n3621 = (~x0 | x1 | ~x2 | ~x4 | ~x5) & (x2 | (~x4 ^ x5) | (x0 ^ ~x1));
  assign n3622 = ~n2416 & n3625 & (x0 ? n3624 : n3623);
  assign n3623 = (x1 | x2 | x3 | ~x4 | x7) & (~x3 | (x2 ? ((x4 | x7) & (~x1 | ~x4 | ~x7)) : (x4 | ~x7)));
  assign n3624 = x2 ? (~x7 | ((x3 | x4) & (x1 | ~x3 | ~x4))) : (x7 | ((~x3 | ~x4) & (~x1 | x3 | x4)));
  assign n3625 = (~n3626 | n987) & (~n300 | ~n588 | ~n786);
  assign n3626 = ~x0 & ~x7;
  assign z193 = ~n3629 | n3637 | (x1 & (~n3628 | ~n3640));
  assign n3628 = (x0 | ~x2 | x3 | ~x4 | x5) & (x4 | (x0 ? (x2 ? (x3 | ~x5) : (~x3 | x5)) : ((~x3 | ~x5) & (x2 | x3 | x5))));
  assign n3629 = n3633 & (n1254 | n3631) & (x1 | n3630);
  assign n3630 = (x0 | ~x2 | x3 | x4 | x5) & (~x4 | ((x0 | x2 | x3 | ~x5) & (~x0 | ((~x3 | ~x5) & (x2 | x3 | x5)))));
  assign n3631 = (x2 | n3632) & (x1 | ~x2 | n487 | n1974);
  assign n3632 = (x0 | x1 | x3 | x5 | ~x7) & (~x0 | ~x1 | ~x3 | ~x5 | x7);
  assign n3633 = ~n3634 & (~n408 | ((~n280 | ~n2749) & ~n3636));
  assign n3634 = x0 & ((~x3 & ~n3635) | (~n1354 & n2560));
  assign n3635 = (x1 | x2 | x4 | x5 | x6) & ((x1 ^ ~x2) | (x4 ? (x5 | x6) : (~x5 | ~x6)));
  assign n3636 = n424 & ((~x6 & x7 & ~x0 & x3) | (x0 & x6 & (x3 ^ x7)));
  assign n3637 = ~x0 & (x2 ? ~n3638 : ~n3639);
  assign n3638 = x1 ? ((~x3 | ~x4 | ~x5 | ~x6) & (x5 | x6 | x3 | x4)) : (x3 ? (x4 ? (x5 | x6) : (~x5 | ~x6)) : (~x4 | (~x5 ^ x6)));
  assign n3639 = (x1 | ~x3 | ~x4 | x5 | x6) & ((~x1 ^ ~x4) | (x3 ? (~x5 | ~x6) : (~x5 ^ x6)));
  assign n3640 = (~x6 | ~n335 | ~n782 | n487) & (x6 | n3641);
  assign n3641 = (x3 | n2424) & (~x4 | n2158 | x0 | ~x3);
  assign z194 = ~n3655 | (x5 ? ~n3650 : ~n3643);
  assign n3643 = x1 ? n3646 : (x0 ? n3644 : n3645);
  assign n3644 = (x2 | x7 | ((~x4 | ~x6) & (x3 | x4 | x6))) & (~x3 | ~x4 | x6 | ~x7) & (~x2 | ((~x4 | x6 | ~x7) & (~x3 | (x4 ? x6 : (~x6 | ~x7)))));
  assign n3645 = ((x2 ^ ~x7) | ((x4 | ~x6) & (x3 | ~x4 | x6))) & (~x6 | ~x7 | x3 | x4) & (x2 | ~x3 | ~x4 | x6 | x7);
  assign n3646 = ~n3649 & ((x3 & (x2 | n3648)) | (n3647 & (n3648 | (~x2 & ~x3))));
  assign n3647 = (x0 | ~x2 | x4 | x6 | x7) & (x2 | (x0 ? (x4 ? (x6 | x7) : (~x6 | ~x7)) : (x4 | (~x6 ^ x7))));
  assign n3648 = x0 ? (x7 | (x4 ^ ~x6)) : (~x7 | (x4 ^ x6));
  assign n3649 = ~n1254 & n782 & x3 & ~x7;
  assign n3650 = n3653 & (n1254 | n3652) & (x2 | n3651);
  assign n3651 = (~x0 | x1 | x4 | ~x6 | x7) & (x0 | x6 | (x1 ? (~x4 | ~x7) : (x4 | x7)));
  assign n3652 = x0 ? (x1 ? (x2 | x7) : (~x2 | ~x7)) : (x1 | (x2 ? x7 : (x3 | ~x7)));
  assign n3653 = (~x2 | ~n387 | n485) & (n599 | ~n3654);
  assign n3654 = x7 & x6 & ~x2 & x4;
  assign n3655 = ~n3659 & (x0 ? n3656 : (~n3661 & n3663));
  assign n3656 = ~n3657 & (x4 ? (~n308 | ~n725) : n3658);
  assign n3657 = ~x1 & ((x2 & ~x7 & (~x4 ^ x6)) | (~x6 & x7 & ~x2 & ~x4));
  assign n3658 = (~x1 | ~x2 | x3 | ~x6 | ~x7) & (x1 | x2 | ~x3 | x6 | x7);
  assign n3659 = ~n3660 & (x1 ? (x3 & ~x4) : x4);
  assign n3660 = (~x0 | x2 | ~x6 | ~x7) & (x0 | (x2 ? (x6 | ~x7) : (~x6 | x7)));
  assign n3661 = x3 & ((n282 & n3662) | (n408 & n2131));
  assign n3662 = x6 & (x4 ^ ~x7);
  assign n3663 = (x1 | ~x2 | ~x3 | n485) & (~x1 | (x2 ? (x3 | ~n1498) : n485));
  assign z195 = ~n3679 | n3676 | n3673 | n3665 | n3669;
  assign n3665 = ~x7 & ((n514 & n2289) | n3666);
  assign n3666 = ~x5 & (x3 ? ~n3668 : ~n3667);
  assign n3667 = x0 ? ((~x1 | x2 | x4 | ~x6) & (~x2 | ((~x4 | x6) & (x1 | (~x4 & x6))))) : ((~x1 | (x2 ^ x6)) & (x2 | (x6 ? x1 : ~x4)));
  assign n3668 = (x1 | (x0 ? (~x2 | (x4 & ~x6)) : (x2 | ~x6))) & (x0 | ((x2 | ~x4 | ~x6) & (~x1 | (x2 ? (x4 | ~x6) : x6))));
  assign n3669 = ~n1291 & (n3671 | ~n3672 | (x6 & ~n3670));
  assign n3670 = (x0 | x1 | ~x2 | x3 | ~x4) & (~x1 | ((x3 | x4 | x0 | x2) & (~x0 | (x2 ? (x3 | x4) : (~x3 | ~x4)))));
  assign n3671 = n3596 & (n1416 | (~x0 & x3 & ~n736));
  assign n3672 = (x0 | x1 | ~x2 | x3 | x6) & ((~x1 ^ x6) | (x0 ? x2 : (~x2 | ~x3)));
  assign n3673 = ~x0 & (x2 ? ~n3674 : ~n3675);
  assign n3674 = (x1 | ~x3 | ~x4 | x5 | x6) & (x4 | ~x5 | (x1 ? (~x3 ^ ~x6) : (x3 | ~x6)));
  assign n3675 = (~x1 | x5 | ~x6 | (x3 ^ ~x4)) & (x1 | x3 | ~x4 | ~x5 | x6);
  assign n3676 = n786 & (n3677 | ~n3678);
  assign n3677 = ~x2 & ((~x0 & (x1 ? (x3 & ~x6) : x6)) | (x0 & ~x1 & x3 & ~x6));
  assign n3678 = x3 ? (~x6 | n405) : ((x6 | n405) & (~x2 | ~x6 | n755));
  assign n3679 = ~n3682 & (~x0 | (~n3681 & (x3 | n3680)));
  assign n3680 = (~x1 | ((~x5 | ~x6 | x2 | ~x4) & (x5 | x6 | ~x2 | x4))) & (x1 | ~x2 | x4 | x5 | ~x6);
  assign n3681 = ~x6 & n923 & (x2 ? x5 : (~x4 & ~x5));
  assign n3682 = ~n310 & ((n301 & n514) | (~x2 & ~n3683));
  assign n3683 = (x0 | x1 | x4 | ~x5 | x6) & (~x0 | ((x5 | x6 | x1 | ~x4) & (~x5 | ~x6 | ~x1 | x4)));
  assign z196 = ~n3698 | ~n3694 | ~n3690 | n3685 | n3687;
  assign n3685 = x2 & ((n728 & n1476) | (x3 & ~n3686));
  assign n3686 = (x5 | ~n3662 | x0 | ~x1) & (~x0 | x1 | n1851);
  assign n3687 = ~n565 & (~n3688 | (~x4 & ~n605 & n923));
  assign n3688 = ~n3689 & (n2504 | ~n913) & (~n514 | ~n1265);
  assign n3689 = ~x4 & ~x3 & x1 & x2;
  assign n3690 = n3692 & (~x4 | n1792 | ~n3691);
  assign n3691 = x2 & ~x0 & x1;
  assign n3692 = (~n595 | ~n2076) & (~n423 | n3693);
  assign n3693 = x1 ? (x6 | (~x4 & x7)) : (~x4 | ~x6);
  assign n3694 = (x4 | n3695) & (~n725 | n3697);
  assign n3695 = x3 ? (~n782 | n3696) : (~n382 | ~n428);
  assign n3696 = x1 ? (~x6 | ~x7) : (x6 | x7);
  assign n3697 = (x3 | ~x4 | ~x5 | x6 | x7) & (~x3 | x4 | ~x7 | (x5 ^ ~x6));
  assign n3698 = (x3 | n3699) & (x1 | (~n2114 & ~n3700));
  assign n3699 = (x1 | ~x2 | ((x6 | x7) & (x4 | ~x6 | ~x7))) & (x2 | ((x1 | x4 | x6 | ~x7) & (~x1 | ~x6 | (x4 & ~x7))));
  assign n3700 = ~x6 & ((n339 & n1422) | (n493 & ~n766));
  assign z197 = n3705 | ~n3707 | (~x2 & (n3702 | n3704));
  assign n3702 = x0 & (n3703 | (x6 & n910 & n1876));
  assign n3703 = ~x7 & ((n625 & n764) | (~x1 & ~n2903));
  assign n3704 = n285 & n450 & ((x4 & ~x6) | (~x1 & ~x4 & x6));
  assign n3705 = ~n998 & ((n659 & n886) | (n341 & ~n3706));
  assign n3706 = (x5 & (~x3 | (~x0 & ~x1))) | (x0 & x1) | (x3 & ~x5);
  assign n3707 = n3708 & ~n3712 & n3713 & (n453 | n2555);
  assign n3708 = ~n3709 & ~n3711 & (~x3 | ~n782 | ~n1863);
  assign n3709 = ~n3710 & ~x4 & n857;
  assign n3710 = (~x1 | x2 | ~x5 | x7) & (x1 | ~x2 | (x5 ^ x7));
  assign n3711 = ~x0 & ((n1986 & n662) | (n1658 & n1187));
  assign n3712 = n339 & ((x4 & n786) | (x0 & ~x4 & n450));
  assign n3713 = n3714 & (~n425 | ~n521 | ~n426 | n470);
  assign n3714 = (~x4 | x7 | x2 | ~x3) & (~x2 | x3 | x4 | ~x7);
  assign z198 = ~n3719 | n3716 | (x5 & ~n310 & ~n3718);
  assign n3716 = x0 & ((~x6 & ~n3717) | (n725 & n1704));
  assign n3717 = (~x1 | x2 | (x3 ? (x4 ^ x5) : (~x4 | x5))) & (x1 | ~x2 | x3 | x4 | ~x5);
  assign n3718 = (x0 | ((x4 | x6) & (~x1 | ~x4 | ~x6))) & (~x4 | ~x6 | ~x1 | x2) & (x1 | ((x2 | x4 | x6) & (~x0 | ~x4 | ~x6)));
  assign n3719 = ~n3723 & ~n3722 & ~n3721 & ~n1420 & ~n3720;
  assign n3720 = x5 & x4 & x3 & ~x0 & ~x1;
  assign n3721 = ~n470 & ((n587 & n588) | (~x3 & ~n673));
  assign n3722 = ~x4 & ((x0 & x1 & ~x3 & x5) | (x3 & ~x5 & (~x0 | ~x1)));
  assign n3723 = ~n1331 & n588 & x5 & ~x6;
  assign z199 = ~n3729 | (x0 & ~n3725) | (x5 & ~n3727);
  assign n3725 = (x7 | n3726) & (x3 | ~n282 | ~n633);
  assign n3726 = (x1 | x2 | ~x3 | ~n320) & (~x1 | ~x2 | x3 | ~n2085);
  assign n3727 = (x0 & ((x2 & ~n1147) | (x1 & (x2 | ~n1147)))) | (~n3728 & (~n1147 | (~x0 & ~x1)));
  assign n3728 = ~x6 & (x4 ^ ~x7);
  assign n3729 = ~n3730 & (~n441 | ~n301) & (~n2085 | n2575);
  assign n3730 = ~n271 & ((n1039 & n559) | n2085);
  assign z200 = ~n3734 | (~n1291 & (n2777 | ~n3732 | n3733));
  assign n3732 = x0 ? ((x1 & x2) | ~x6) : (x6 & (~x1 | (~x2 & ~n590)));
  assign n3733 = ~x2 & ((x3 & x6 & ~x0 & x1) | (~x3 & ~x6 & x0 & ~x1));
  assign n3734 = n3737 & (~n1921 | ~n2778) & (n3735 | ~n3736);
  assign n3735 = (~x0 | ~x2 | ~x4 | x5 | x6) & (x0 | x2 | x4 | ~x5 | ~x6);
  assign n3736 = ~x7 & x1 & ~x3;
  assign n3737 = (x0 | x1 | ~x5 | ~x6) & (~x0 | x5 | x6 | (x1 ^ ~x2));
  assign z201 = ~n3744 | n3743 | n3742 | n3739 | ~n3741;
  assign n3739 = ~x2 & ((n2131 & n728) | n3740);
  assign n3740 = n955 & (x0 ? (x3 & ~n1254) : (~x3 & n700));
  assign n3741 = (~x0 & (x6 | x7)) | (x1 & x2) | (x6 & x7) | (~x7 & ((~x1 & ~x2) | (x0 & ~x6)));
  assign n3742 = n1837 & ((n363 & n3607) | (n659 & ~n1486));
  assign n3743 = n1747 & ~x3 & n1179;
  assign n3744 = ~n3745 & (~n579 | ~n606 | n3746);
  assign n3745 = ~x0 & (x1 ? (x2 & ~x6) : (x6 & x7));
  assign n3746 = (x1 | ~x5 | x6 | x7) & (~x1 | ~x7 | (x5 ^ ~x6));
  assign z202 = ~n3753 | n3751 | ~n3748 | n3750;
  assign n3748 = ~n3749 & (~n295 | ~n1473) & (~n387 | ~n3141);
  assign n3749 = ~x2 & ~x7 & (x0 ? (~x1 & ~x3) : (x1 & x3));
  assign n3750 = n625 & ((n324 & n760) | (n579 & n1074));
  assign n3751 = ~n3752 & n366 & n327;
  assign n3752 = (~x0 | x1 | ~x3 | ~x7) & (x0 | ~x1 | x3 | x7);
  assign n3753 = (~x7 | ~n441) & (~x0 | (~n3754 & (~x7 | n271)));
  assign n3754 = ~x1 & ~x2 & x3 & (~x4 ^ x7);
  assign z203 = n3756 | n3759 | ~n3760 | (~x2 & ~n3758);
  assign n3756 = ~x7 & ((n295 & n1161) | n3757);
  assign n3757 = x0 & ((n272 & n494) | (n764 & n1127));
  assign n3758 = (x0 | ((~x4 | ~x5 | x1 | ~x3) & (x4 | x5 | ~x1 | x3))) & (~x0 | x1 | ~x3 | x4 | x5);
  assign n3759 = x5 & ((n3297 & n428) | (n514 & n590));
  assign n3760 = x0 ? ((x2 | x3) & (~x1 | (x2 & (x3 | x4)))) : (~x2 | (x1 & ~x3));
  assign z204 = ~n3771 | n3770 | n3769 | ~n3762 | n3767;
  assign n3762 = (~n3763 | n3764) & (~n423 | (n3765 & n3766));
  assign n3763 = x6 & ~x4 & ~x1 & ~x2;
  assign n3764 = (x0 | x3 | ~x5 | ~x7) & (~x0 | (x3 ? (~x5 | x7) : (x5 | ~x7)));
  assign n3765 = (~x0 | x1 | x4 | x5) & (x0 | ~x4 | (~x1 ^ ~x5));
  assign n3766 = (~x0 | x4 | ~x5 | (~x1 ^ ~x6)) & (x0 | ~x1 | ~x4 | x5 | ~x6);
  assign n3767 = n3440 & (x0 ? ~n3768 : (~x2 & ~n1861));
  assign n3768 = (~x2 | x3 | ~x4 | x5 | x7) & (x2 | ~x3 | x4 | ~x5 | ~x7);
  assign n3769 = ~x0 & ((~x1 & ((x3 & ~x4) | (~x2 & ~x3 & x4))) | (x2 & (x1 ? (~x3 & ~x4) : x3)));
  assign n3770 = x0 & (x1 ? (x2 ? (~x3 & ~x4) : (x3 & x4)) : (x2 ? x3 : (~x3 & x4)));
  assign n3771 = (~n514 | ~n2289) & (x3 | n1011 | n868);
  assign z205 = n3775 | n3777 | ~n3780 | (~n1274 & ~n3773);
  assign n3773 = x2 ? (x1 | (~x4 & ~n494)) : n3774;
  assign n3774 = (~x1 | ((x4 | x6 | x7) & (~x4 | ~x5 | ~x6 | ~x7))) & (x4 | ((x1 | (~x6 ^ x7)) & (~x5 | x6 | x7) & (x5 | (~x6 & ~x7))));
  assign n3775 = ~x1 & ((~x5 & ~n3776) | (n301 & n661));
  assign n3776 = (x0 | ~x2 | ~x3 | ~x4 | ~x6) & (x4 | ((x0 | x2 | ~x3 | ~x6) & (~x0 | x3 | (~x2 ^ ~x6))));
  assign n3777 = ~x5 & (n3779 | (n647 & n709 & ~n3778));
  assign n3778 = x1 ? (~x4 | ~x7) : (x4 | x7);
  assign n3779 = ~x6 & (n2878 | (x3 & n342 & n428));
  assign n3780 = ~n3782 & ~n3783 & n3784 & (~x1 | n3781);
  assign n3781 = x0 ? (x3 | (x2 ? x4 : (~x4 | ~x5))) : (~x3 | (~x2 ^ ~x4));
  assign n3782 = ~n614 & ((n363 & n426) | (~x0 & ~n1516));
  assign n3783 = n594 & n308 & n284;
  assign n3784 = (~n514 | ~n2289) & (~n300 | ~n612);
  assign z206 = ~n3796 | ~n3793 | n3786 | ~n3789;
  assign n3786 = ~x3 & ((n364 & n1145) | n3787);
  assign n3787 = ~x7 & ((n359 & n494) | (n1921 & ~n3788));
  assign n3788 = (x1 | ~x2 | x4 | x6) & (~x1 | ~x4 | (~x2 ^ x6));
  assign n3789 = n3790 & ~n3791 & (n1254 | n1274 | n3792);
  assign n3790 = (n673 | n1652) & (n498 | n755);
  assign n3791 = n659 & n327 & (x1 ? x4 : (~x2 & ~x4));
  assign n3792 = (x5 | ~x7 | x1 | ~x2) & (~x1 | x2 | ~x5 | x7);
  assign n3793 = n3795 & (n822 | n3794) & (n976 | n3338);
  assign n3794 = (x0 | ~x1 | ~x2 | x5 | ~x7) & (~x0 | x1 | x2 | ~x5 | x7);
  assign n3795 = ~n408 | (x0 ? (~n606 | ~n328) : ~n609);
  assign n3796 = (n2158 | n3798) & (n377 | n3797);
  assign n3797 = x0 ? (~x3 | (x1 ? (x2 | ~x4) : x4)) : (x3 | (~x1 ^ ~x4));
  assign n3798 = (~x0 | x1 | x3 | x4 | ~x6) & (x0 | ~x3 | x6 | (~x1 ^ ~x4));
  assign z207 = ~n3800 | (x5 ? ~n3813 : (n3808 | ~n3810));
  assign n3800 = ~n3804 & (x1 | (~n3801 & n3802));
  assign n3801 = ~n1254 & ((~x0 & ~x2 & x3 & ~x7) | ((x2 ^ x7) & (x0 | ~x3)));
  assign n3802 = (~n413 | ~n2131) & (~x6 | n3803);
  assign n3803 = (x0 | x2 | ~x3 | ~x4 | ~x7) & (~x0 | x3 | (x2 ? (~x4 | ~x7) : (x4 | x7)));
  assign n3804 = x1 & (n3806 | n3807 | (~x2 & ~n3805));
  assign n3805 = (x0 | ~x3 | x4 | ~x6 | ~x7) & (~x4 | (x0 ? (x3 | (~x6 ^ x7)) : (x6 | x7)));
  assign n3806 = ~n836 & ((x0 & ~x2 & x3 & x7) | (~x0 & ~x3 & (x2 ^ x7)));
  assign n3807 = x6 & n624 & ((~x3 & x7) | (~x0 & x3 & ~x7));
  assign n3808 = ~x0 & ((~x2 & ~n3809) | (n1114 & n634));
  assign n3809 = (~x6 | x7 | ~x1 | x4) & (x1 | ~x4 | (x3 ? (x6 | ~x7) : (~x6 | x7)));
  assign n3810 = n3812 & (n836 | n3811) & (n485 | n1652);
  assign n3811 = (x0 | x1 | ~x2 | x3 | ~x7) & (~x0 | ((~x3 | ~x7 | x1 | ~x2) & (~x1 | x7 | (x2 ^ ~x3))));
  assign n3812 = ~n2450 & (~n308 | ~n356 | ~n394);
  assign n3813 = n3818 & (x2 ? n3814 : (~n3816 & ~n3817));
  assign n3814 = (~n2131 | ~n728) & (x1 | n3815);
  assign n3815 = (x0 | ~x3 | ~x4 | ~x6 | ~x7) & (~x0 | x3 | x4 | (~x6 ^ x7));
  assign n3816 = x1 & ((n659 & n2131) | (n1064 & ~n975));
  assign n3817 = n473 & ((x0 & x3 & x6 & ~x7) | (~x0 & (x3 ? (~x6 & x7) : ~x7)));
  assign n3818 = (n1254 | n3820) & (n485 | n3819);
  assign n3819 = (x0 | ~x1 | ~x2 | ~x3) & (~x0 | x1 | x2 | x3);
  assign n3820 = (x0 | x1 | ~x2 | ~x3 | x7) & ((x1 ? (x2 | x7) : (~x2 | ~x7)) | (~x0 ^ ~x3));
  assign z208 = ~n3836 | n3834 | ~n3830 | n3822 | n3825;
  assign n3822 = ~n703 & (n3824 | (~x5 & ~n3823));
  assign n3823 = (x0 | x2 | ~x7 | (x3 ^ x6)) & (x7 | ((x3 | ((~x0 | x2 | ~x6) & (~x2 | x6))) & (x0 | (x2 ? ~x6 : (~x3 | x6)))));
  assign n3824 = x7 & n730 & (x2 ^ (x3 & ~x6));
  assign n3825 = ~n1291 & (n3827 | ~n3828 | (x3 & ~n3826));
  assign n3826 = (x0 | x1 | ~x2 | x6) & (x2 | ((x0 | ~x1 | x4 | ~x6) & (~x0 | (x1 ? (~x4 | x6) : (x4 | ~x6)))));
  assign n3827 = ~x2 & (x0 ? (x3 ? (~x4 ^ x6) : (x4 & ~x6)) : (~x3 & x6));
  assign n3828 = ~n3829 & (x4 | x6 | ~n339 | n1331);
  assign n3829 = x6 & ~x4 & ~x3 & x0 & x2;
  assign n3830 = ~n3833 & (x3 | (x1 & n3832) | (~x1 & n3831));
  assign n3831 = x0 ? (~x6 | (x2 ? (~x4 | x5) : (x4 | ~x5))) : (~x4 | x6 | (~x2 ^ ~x5));
  assign n3832 = (~x0 | ((~x5 | ~x6 | x2 | ~x4) & (x5 | x6 | ~x2 | x4))) & (x0 | ~x2 | x4 | x5 | ~x6);
  assign n3833 = n3347 & ((n700 & n363) | (~x0 & ~n770));
  assign n3834 = n327 & ((n514 & n2006) | (~x2 & ~n3835));
  assign n3835 = (x0 | x1 | ~x3 | ~x4 | ~x7) & (~x0 | x7 | (x1 ? (~x3 | x4) : (x3 | ~x4)));
  assign n3836 = ~n3839 & (n570 | (x2 & n3838) | (~x2 & n3837));
  assign n3837 = (x0 | x1 | ~x3 | ~x4 | x6) & (~x0 | ~x1 | x3 | x4 | ~x6);
  assign n3838 = x0 ? (x1 | (~x3 ^ (x4 & ~x6))) : ((~x4 | ~x6 | x1 | x3) & (~x1 | x4 | (x3 ^ x6)));
  assign n3839 = ~x6 & (x2 ? ~n3840 : (x5 & ~n3841));
  assign n3840 = (~n363 | n2979) & (x7 | ~n380 | n677);
  assign n3841 = (~x0 | ~x1 | x3 | x4 | x7) & (x0 | ~x7 | (x1 ? (~x3 | x4) : (x3 | ~x4)));
  assign z209 = n3847 | ~n3856 | (x3 ? ~n3851 : ~n3843);
  assign n3843 = x2 ? n3846 : (~n3845 & (x5 | n3844));
  assign n3844 = (x0 | ~x1 | x4 | x6 | x7) & (x1 | ~x4 | ((~x6 | ~x7) & (~x0 | x6 | x7)));
  assign n3845 = n981 & (x1 ? (x4 & n717) : (~x4 & ~n542));
  assign n3846 = (~n601 | ~n921) & (n542 | (~n896 & ~n1483));
  assign n3847 = ~n565 & (~n3849 | (~x3 & ~n3848));
  assign n3848 = (x0 | x1 | ~x2 | x4 | ~x5) & (x2 | ((~x0 | ~x1 | x4 | x5) & (x0 | ~x4 | (~x1 ^ ~x5))));
  assign n3849 = ~n2793 & ~n3850 & (~x3 | n1011 | n868);
  assign n3850 = ~x0 & ((x1 & x2 & x3 & ~x4) | (~x1 & ~x3 & (~x2 ^ x4)));
  assign n3851 = ~n3852 & n3853 & (n542 | n614 | ~n1241);
  assign n3852 = ~n1091 & ((n363 & n635) | (n387 & n1370));
  assign n3853 = n3855 & (n3854 | (x1 ? (x4 | x5) : (~x4 | ~x5)));
  assign n3854 = (~x0 | x2 | ~x6 | ~x7) & (x0 | ~x2 | x6 | x7);
  assign n3855 = (~n364 | ~n635) & (~n300 | ~n1370);
  assign n3856 = ~n3859 & n3860 & (x0 | (~n3857 & ~n3858));
  assign n3857 = x2 & ((n301 & n620) | (n276 & n458));
  assign n3858 = n408 & ((n327 & n356) | (x3 & ~n2519));
  assign n3859 = ~x2 & n363 & (n757 | (~x3 & ~n2519));
  assign n3860 = ~n3862 & (n614 | n3861) & (~x0 | n1878);
  assign n3861 = x0 ? ((~x1 | x2 | x3 | ~x6) & (x1 | ~x2 | ~x3 | x6)) : (~x1 | x2 | (x3 ^ x6));
  assign n3862 = n782 & ((n700 & n625) | (n1683 & n923));
  assign z210 = n3864 | ~n3867 | (x5 ? ~n3877 : ~n3873);
  assign n3864 = ~x0 & (x1 ? ~n3865 : ~n3866);
  assign n3865 = x2 ? ((x5 | ~x7 | x3 | x4) & (~x3 | ~x4 | ~x5 | x7)) : ((x3 | ~x5 | (x4 ^ x7)) & (x5 | ((~x4 | x7) & (~x3 | x4 | ~x7))));
  assign n3866 = (x2 | ~x3 | ~x7 | (x4 ^ ~x5)) & (x7 | ((~x2 | x3 | x4 | x5) & (x2 | (x3 ? (x4 | x5) : (~x4 | ~x5)))));
  assign n3867 = ~n3868 & (x2 ? n3872 : n3871);
  assign n3868 = x0 & ((~x1 & ~n3869) | (n725 & ~n3870));
  assign n3869 = x2 ? (~x3 | (x4 ? (x5 ^ x7) : (~x5 | x7))) : (x4 ? (x5 | ~x7) : ((x5 | x7) & (x3 | ~x5 | ~x7)));
  assign n3870 = (x4 | x5 | ~x7) & (x3 | x7 | (x4 ^ ~x5));
  assign n3871 = (x0 | x1 | x3 | x4 | ~x7) & (~x0 | ~x1 | ~x3 | ~x4 | x7);
  assign n3872 = x4 ? ((x1 | x3 | ~x7) & (x0 | (x1 ? (x3 | x7) : ~x7))) : ((~x1 ^ ~x7) | (x0 ^ ~x3));
  assign n3873 = ~n3874 & (~n514 | ~n2492) & (n565 | n3876);
  assign n3874 = ~x1 & ((n413 & n634) | (x7 & ~n3875));
  assign n3875 = (x0 | x2 | x3 | ~x4 | x6) & (~x0 | ~x6 | (x2 ? (~x3 | ~x4) : (x3 | x4)));
  assign n3876 = (~x0 | x1 | ~x2 | ~x3 | x4) & (x0 | ~x1 | (x2 ? (~x3 | ~x4) : (x3 | x4)));
  assign n3877 = ~n3879 & ~n3880 & (n542 | n3878);
  assign n3878 = (x0 | x1 | ~x2 | x3 | x4) & (x2 | ((~x3 | ~x4 | x0 | ~x1) & (~x0 | (x1 ? (x3 | ~x4) : (~x3 | x4)))));
  assign n3879 = ~x3 & ((n428 & n622) | (n345 & n514));
  assign n3880 = n423 & ~n1016 & (x0 ? n308 : n521);
  assign z211 = n3882 | ~n3887 | n3895 | (x0 & ~n3898);
  assign n3882 = ~n350 & (n3883 | ~n3885 | (~x0 & ~n3884));
  assign n3883 = x0 & ((~x1 & x2 & ~x3 & x5) | (~x2 & ((~x3 & ~x5) | (x1 & x3 & x5))));
  assign n3884 = (~x1 | x5 | x6 | (x2 ^ x3)) & (~x5 | ~x6 | ((~x2 | ~x3) & (x1 | x2 | x3)));
  assign n3885 = ~n3886 & (x0 ? (~n438 | ~n807) : n1116);
  assign n3886 = ~n377 & (n2786 | (~x0 & (n628 | n1114)));
  assign n3887 = n3890 & (x0 | (n3889 & (~n346 | n3888)));
  assign n3888 = (~x2 | ((~x6 | ~x7 | x3 | x4) & (~x3 | ~x4 | x6 | x7))) & (x2 | x3 | ~x4 | x6 | ~x7);
  assign n3889 = (~n1127 | ~n1145) & (n310 | n1254 | n1119);
  assign n3890 = x2 ? (n3892 & (~x1 | x5 | n3891)) : (~x5 | n3891);
  assign n3891 = (~x0 | x3 | ~x4 | x6 | x7) & (x0 | ((~x6 | ~x7 | x3 | x4) & (~x3 | ~x4 | x6 | x7)));
  assign n3892 = x1 ? (~x5 | n3894) : n3893;
  assign n3893 = x0 ? ((~x5 | ~x7 | x3 | x4) & (~x3 | ~x4 | x5 | x7)) : (~x5 | (x3 ? (x4 | ~x7) : (~x4 | x7)));
  assign n3894 = (~x0 | x3 | x4 | ~x7) & (x0 | (x3 ? (x4 | ~x7) : (~x4 | x7)));
  assign n3895 = ~x2 & (~n3897 | (~x5 & ~n3896));
  assign n3896 = (~x0 | ~x1 | x3 | x4 | ~x7) & (x1 | ((~x4 | x7 | x0 | ~x3) & (~x0 | (x3 ? (x4 | ~x7) : (~x4 | x7)))));
  assign n3897 = (~x0 | ~x3 | ~x4 | ~x5 | x7) & (x0 | x5 | (x3 ? (x4 | ~x7) : (~x4 | x7)));
  assign n3898 = ~n3899 & (x4 | (~n3901 & (~x6 | n3900)));
  assign n3899 = ~n1597 & ((n725 & ~n555) | (n438 & n556));
  assign n3900 = (x1 | ~x2 | ~x3 | ~x5 | ~x7) & (~x1 | ((x2 | ~x3 | x5 | ~x7) & (~x2 | x3 | ~x5 | x7)));
  assign n3901 = x7 & n3596 & (x2 ? (x3 & ~x5) : (~x3 ^ x5));
  assign z212 = ~n3903 | n3915 | n3920 | (~x1 & ~n3918);
  assign n3903 = ~n3904 & ~n3907 & n3910 & (n485 | n3906);
  assign n3904 = x1 & ((~x2 & ~n3905) | (n458 & n720));
  assign n3905 = (x0 | ~x3 | ~x4 | ~x5 | x6) & (x4 | x5 | (x0 ? (~x3 ^ x6) : (x3 | x6)));
  assign n3906 = (x0 | x1 | ~x2 | ~x3 | ~x5) & (~x1 | ((x0 | x2 | ~x3 | x5) & (~x0 | x3 | (~x2 ^ x5))));
  assign n3907 = ~n542 & (n3909 | (~x3 & n647 & n3908));
  assign n3908 = x4 & (~x1 ^ ~x5);
  assign n3909 = ~n1016 & ((n324 & n314) | (n659 & ~n1091));
  assign n3910 = ~n3914 & (~x2 | (~n3911 & ~n3912 & n3913));
  assign n3911 = ~n753 & ((n363 & n341) | (n387 & n342));
  assign n3912 = n2653 & ((~x1 & n308) | (n521 & n620));
  assign n3913 = (x0 | x1 | x3 | x4 | x6) & ((~x3 ^ x6) | (x0 ? (x1 | x4) : (~x1 | ~x4)));
  assign n3914 = n740 & ((x0 & x1 & x3 & x4) | (~x0 & (x1 ? (~x3 & x4) : (x3 & ~x4))));
  assign n3915 = ~x2 & ((n1008 & n1755) | n3916);
  assign n3916 = x4 & ((~x5 & ~n3917) | (n656 & n457));
  assign n3917 = (~x7 | ((~x1 | ~x3 | x6) & (x0 | (x1 ? x6 : (~x3 | ~x6))))) & (x1 | ~x6 | x7 | (~x0 ^ ~x3));
  assign n3918 = (~x6 | n3919) & (x2 | x6 | n614 | n1274);
  assign n3919 = (~x0 | x2 | x3 | (~x4 ^ x5)) & (~x2 | ((~x4 | ~x5 | ~x0 | ~x3) & (x0 | (x3 ? (x4 | x5) : (~x4 | ~x5)))));
  assign n3920 = ~n565 & ((n857 & ~n1803) | (~x3 & ~n3921));
  assign n3921 = (x0 | ~x1 | x4 | ~x5) & (x1 | ((x4 | x5 | ~x0 | x2) & (x0 | ~x4 | (~x2 ^ x5))));
  assign z213 = ~n3931 | (~x3 & ~n3928) | (~x7 & ~n3923);
  assign n3923 = ~n3926 & (x1 | (~n3925 & (x2 | n3924)));
  assign n3924 = (~x0 | x3 | x4 | ~x5 | x6) & (x0 | x5 | ~x6 | (x3 ^ x4));
  assign n3925 = n278 & ((n659 & n1039) | (x0 & ~n753));
  assign n3926 = n625 & ~n3927;
  assign n3927 = (~x2 | x5 | ((x4 | ~x6) & (~x0 | ~x4 | x6))) & (~x0 | x2 | ~x5 | (~x4 ^ x6));
  assign n3928 = ~n3930 & (~n394 | ~n1183) & (~x1 | n3929);
  assign n3929 = (~x0 | x2 | ~x4 | ~x5 | ~x7) & (~x2 | ((x4 | ~x5 | x7) & (x5 | ~x7 | x0 | ~x4)));
  assign n3930 = ~n688 & ((~x2 & ~n1417) | (n438 & ~n566));
  assign n3931 = ~n3933 & ~n3935 & ~n3938 & (n350 | n3932);
  assign n3932 = (~x0 | x1 | x2 | x3 | x5) & (~x1 | ((x2 | ~x3 | ~x5) & (x0 | (x2 ? (~x3 | x5) : ~x5))));
  assign n3933 = ~n3934 & (n834 | (~x2 & n2085));
  assign n3934 = (~x0 | x1 | ~x3 | ~x7) & (x0 | (x1 ? (~x3 | x7) : (x3 | ~x7)));
  assign n3935 = x3 & ((n428 & n662) | n3936 | n3937);
  assign n3936 = n2773 & ((n725 & n425) | (~x1 & ~n2933));
  assign n3937 = ~n688 & ((n484 & n480) | (~x1 & ~n1091));
  assign n3938 = ~n1486 & (x5 ? (n782 & ~n822) : ~n3939);
  assign n3939 = x0 ? ((~x4 | ~x6 | x2 | ~x3) & (x4 | x6 | ~x2 | x3)) : (x2 | (x3 ? (x4 | x6) : (~x4 | ~x6)));
  assign z214 = n3946 | ~n3950 | (x0 ? ~n3948 : ~n3941);
  assign n3941 = x2 ? (x1 ? n3942 : n3943) : n3944;
  assign n3942 = x3 ? ((~x4 | ~x5 | x6 | ~x7) & (~x6 | x7 | x4 | x5)) : ((x6 | ~x7 | x4 | x5) & (~x4 | ~x6 | (x5 ^ x7)));
  assign n3943 = x3 ? (x6 | ((~x5 | ~x7) & (~x4 | x5 | x7))) : (~x6 | ((x5 | x7) & (x4 | ~x5 | ~x7)));
  assign n3944 = n3945 & (n1291 | n703 | n1163);
  assign n3945 = (x1 | ~x3 | ~x4 | ~n294) & (~x1 | x3 | x4 | ~n556);
  assign n3946 = x3 & ((n295 & n971) | (~x1 & ~n3947));
  assign n3947 = (x0 | ~x2 | x4 | x5 | x6) & (~x0 | ~x5 | (x2 ? (~x4 | ~x6) : (x4 | x6)));
  assign n3948 = ~n3949 & (n1262 | n2925) & (~n269 | ~n1476);
  assign n3949 = ~n731 & (~n791 | (n408 & n424));
  assign n3950 = n3953 & (x3 | ((~n441 | ~n3951) & n3952));
  assign n3951 = x5 & (x2 ? (x4 & x6) : (~x4 & ~x6));
  assign n3952 = (~n364 | ~n458) & (n836 | n581);
  assign n3953 = ~n3955 & (n791 | n3954) & (n377 | n3956);
  assign n3954 = x0 ? (x3 ^ ~x6) : (x3 | x6);
  assign n3955 = n659 & ((~x1 & ~x2 & ~x5 & x6) | (x2 & ((x5 & x6) | (x1 & ~x5 & ~x6))));
  assign n3956 = x0 ? ((~x3 | ~x4 | x1 | x2) & (~x1 | ~x2 | x3 | x4)) : (x2 | (x1 ? (~x3 | x4) : (x3 | ~x4)));
  assign z215 = n3962 | ~n3968 | (x5 ? ~n3958 : ~n3965);
  assign n3958 = n3960 & (x0 | (~n3959 & (~x7 | n3389)));
  assign n3959 = n955 & ((n426 & n1964) | (n1837 & ~n436));
  assign n3960 = (n506 | n3961) & (~n717 | ~n356 | ~n428);
  assign n3961 = (x0 | ~x1 | ~x2 | x4 | x7) & (~x0 | ((~x1 | x2 | x4 | ~x7) & (x1 | ~x2 | ~x4 | x7)));
  assign n3962 = x7 & ((~x6 & ~n3963) | (n3222 & ~n3964));
  assign n3963 = (x0 | x1 | x2 | ~x3 | x4) & (x3 | ((x0 | ~x1 | ~x2 | x4) & (~x0 | ~x4 | (x1 ^ ~x2))));
  assign n3964 = (~x0 | x1 | ~x3 | ~x4) & (x0 | (x1 ? (~x3 | x4) : (x3 | ~x4)));
  assign n3965 = ~n3966 & (n688 | n3967) & (~n428 | ~n996);
  assign n3966 = n3691 & ((n308 & n356) | (x3 & ~n975));
  assign n3967 = x0 ? ((~x1 | x2 | x3 | ~x6) & (x1 | ~x2 | ~x3 | x6)) : (x1 | ~x2 | (x3 ^ x6));
  assign n3968 = n3971 & (n1163 | n3970) & (x2 | n3969);
  assign n3969 = ((x3 ^ x6) | (x0 ? (x1 | ~x4) : (~x1 | x4))) & (~x0 | ~x1 | ~x3 | x4 | x6) & (x0 | x1 | x3 | ~x4 | ~x6);
  assign n3970 = (~x0 | x1 | ~x2 | x4 | x7) & (x0 | ~x1 | x2 | ~x4 | ~x7);
  assign n3971 = ~n3975 & ~n3974 & ~n3972 & n3973;
  assign n3972 = ~n580 & ((x0 & x1 & ~x2 & ~x7) | (~x0 & ~x1 & x7));
  assign n3973 = (~n1498 | ~n1063) & (~n1761 | ~n742);
  assign n3974 = ~n506 & ((n363 & n760) | (n387 & n1074));
  assign n3975 = ~n1028 & ((n717 & n910) | (n382 & n473));
  assign z216 = n3977 | ~n3982 | ~n3987 | (x1 & ~n3980);
  assign n3977 = ~x1 & (x2 ? ~n3979 : ~n3978);
  assign n3978 = (~x0 | x3 | x4 | x5 | ~x7) & (x0 | ~x3 | ~x4 | ~x5 | x7);
  assign n3979 = (x0 & ~x3 & (~x5 | x7)) | (x4 & (~x5 ^ x7)) | (~x4 & (x5 ^ x7)) | (~x0 & x3 & x5 & ~x7);
  assign n3980 = n3981 & (~n663 | (~n790 & (~x3 | ~n789)));
  assign n3981 = (~n629 | ~n661) & (n570 | (~n1416 & ~n898));
  assign n3982 = ~n3985 & (x4 ? (x2 | n3986) : n3983);
  assign n3983 = (n581 | ~n3984) & (x7 | n605 | ~n1907);
  assign n3984 = ~x3 & (~x6 ^ ~x7);
  assign n3985 = ~x4 & ~n1318 & ((x0 & x2 & ~x3) | (~x2 & (~x0 | x3)));
  assign n3986 = x7 ? (~x1 | (x0 & ~x3)) : (x1 | (~x0 & x3));
  assign n3987 = (n791 | n3988) & (~x4 | (~n3989 & ~n3990));
  assign n3988 = (x0 | x3 | x4 | ~x6 | ~x7) & (~x0 | ((~x6 | ~x7 | ~x3 | x4) & (x3 | (x4 ? (~x6 ^ x7) : (x6 | x7)))));
  assign n3989 = ~x3 & (x0 ? ~n2927 : (n282 & n313));
  assign n3990 = n659 & ~n605 & (x1 ? (~x6 & ~x7) : (~x6 ^ ~x7));
  assign z217 = n3992 | ~n3996 | ~n4000 | (~n570 & ~n1356);
  assign n3992 = ~x1 & ((n2514 & n1476) | n3993 | n3995);
  assign n3993 = ~x4 & ((~x5 & ~n3994) | (n921 & n2514));
  assign n3994 = (x0 | x2 | x3 | ~x6 | x7) & (~x7 | ((x0 | x2 | x3 | x6) & (~x0 | ~x2 | (x3 ^ x6))));
  assign n3995 = ~n761 & (n3293 | (n790 & n559));
  assign n3996 = ~n3998 & ((x5 & (~x6 | n3999)) | (n3997 & (n3999 | (~x5 & x6))));
  assign n3997 = (~x0 | ~x1 | ~x2 | x3 | x4) & (x2 | ((x0 | x3 | ~x4) & (~x3 | (~x0 ^ (x1 & ~x4)))));
  assign n3998 = n483 & ((~x1 & ~n1274) | (~x0 & x1 & ~n1597));
  assign n3999 = (x0 | x1 | ~x2 | ~x3 | ~x4) & (~x0 | x2 | x3 | (~x1 ^ ~x4));
  assign n4000 = n4004 & (x0 | n4002) & (n377 | n4001);
  assign n4001 = (~x0 | x1 | ~x2 | x3) & (x0 | ((x2 | ~x3 | ~x4) & (~x1 | ~x2 | x3 | x4)));
  assign n4002 = (x4 | ~n3342 | x1 | ~x3) & (~x1 | n4003);
  assign n4003 = (~x2 | ~x3 | ~x4 | ~x5 | ~x6) & (x2 | x3 | x4 | x5 | x6);
  assign n4004 = (~n647 | n4005) & (~x1 | n4006);
  assign n4005 = (x1 | x3 | ~x4 | x5 | x6) & (~x1 | x4 | (x3 ? (x5 | x6) : (~x5 | ~x6)));
  assign n4006 = x0 ? (~n426 | ~n595) : (n574 | n761);
  assign z218 = n4023 | n4020 | ~n4016 | n4008 | ~n4011;
  assign n4008 = ~n565 & (x1 ? ~n4010 : ~n4009);
  assign n4009 = x0 ? ((x4 | x5 | ~x2 | x3) & (~x3 | ~x4 | (x2 & ~x5))) : ((~x3 | x4) & (~x4 | ~x5 | x2 | x3));
  assign n4010 = x0 ? (x3 | x4) : (~x3 | ((x2 | x4 | ~x5) & (~x4 | (~x2 & x5))));
  assign n4011 = n4012 & (n605 | n4015) & (~x1 | n4014);
  assign n4012 = (~n875 | ~n1471) & (x1 | n4013);
  assign n4013 = x0 ? (x2 | x4 | (~x3 ^ x6)) : (~x2 | ~x4 | (x3 ^ x6));
  assign n4014 = (x0 | ~x2 | ~x3 | x4 | x6) & (~x0 | x2 | ~x4 | (~x3 ^ x6));
  assign n4015 = (~x0 | x1 | ~x3 | ~n634) & (x0 | ~x1 | x3 | (~n633 & ~n634));
  assign n4016 = ~n4018 & (x1 | ((~n971 | ~n2514) & ~n4017));
  assign n4017 = ~n614 & ((~x0 & ~x2 & ~x3 & ~x6) | (x0 & x2 & (~x3 ^ ~x6)));
  assign n4018 = n387 & ~n4019;
  assign n4019 = (~x2 | x3 | x4 | x5 | ~x6) & (x2 | ((~x3 | (x4 ? (~x5 | ~x6) : (x5 | x6))) & (x3 | ~x4 | ~x5 | x6)));
  assign n4020 = ~n542 & (n4022 | (~x3 & ~n4021));
  assign n4021 = (x1 | ((x4 | x5 | x0 | ~x2) & (~x0 | ~x4 | (x2 & ~x5)))) & (x0 | ~x1 | (x2 ? (~x4 | x5) : (x4 | ~x5)));
  assign n4022 = ~x4 & n857 & (x1 ? ~x2 : (x2 & ~x5));
  assign n4023 = ~x3 & ((n296 & n359) | n4024);
  assign n4024 = ~x4 & ((n480 & ~n2624) | (~x1 & ~n4025));
  assign n4025 = (~x0 | ~x2 | x5 | ~x6 | ~x7) & (x0 | ((~x6 | ~x7 | x2 | x5) & (~x2 | ~x5 | x6 | x7)));
  assign z219 = ~n4035 | n4033 | n4027 | n4029;
  assign n4027 = n1074 & ((n2431 & n514) | (~x1 & ~n4028));
  assign n4028 = (x0 | x2 | ~x5 | x6) & (~x3 | ((~x0 | x6 | (~x2 ^ ~x5)) & (x0 | ~x2 | x5 | ~x6)));
  assign n4029 = ~x4 & ((n1151 & ~n4032) | (x2 & ~n4030));
  assign n4030 = (x5 | x6 | n1318 | ~n1064) & (~x5 | n4031);
  assign n4031 = (~x0 | x1 | ~x3 | ~x6 | x7) & (x0 | ~x7 | (x1 ? (~x3 | ~x6) : (x3 | x6)));
  assign n4032 = (~x0 | ~x1 | x3 | ~x5 | x6) & (x0 | ((~x1 | x5 | ~x6) & (x1 | ~x3 | ~x5 | x6)));
  assign n4033 = ~n350 & ((n352 & n514) | (~x2 & ~n4034));
  assign n4034 = (x0 | ~x1 | x3 | x5 | x6) & (~x6 | ((x0 | x1 | ~x3 | ~x5) & (~x0 | (x1 ? (x3 | ~x5) : (~x3 | x5)))));
  assign n4035 = ~n4036 & n4040 & (~x5 | ~n387 | n4039);
  assign n4036 = ~x1 & (n4038 | (x3 & ~n4037));
  assign n4037 = (~x0 | ~x2 | ~x4 | ~x5 | ~x7) & (x5 | (~x0 ^ ~x2) | (~x4 ^ x7));
  assign n4038 = ~x5 & n285 & ((~x4 & x7) | (~x2 & x4 & ~x7));
  assign n4039 = (x2 | ~x4 | x7) & (x3 | x4 | ~x7);
  assign n4040 = ~n4042 & ~n4043 & n4044 & (~x0 | ~n4041);
  assign n4041 = x1 & ((x2 & ~x3 & ~x4 & x7) | (~x2 & x3 & x4 & ~x7));
  assign n4042 = ~n350 & ((n441 & n2106) | (~n388 & ~n868));
  assign n4043 = ~n2004 & ((n725 & n760) | (n438 & n1074));
  assign n4044 = x4 ? ((~x7 | n3819) & (x3 | x7 | n420)) : ((x7 | n3819) & (~x3 | ~x7 | n420));
  assign z220 = ~n4046 | (x6 ? ~n4056 : (n4060 | n4062));
  assign n4046 = ~n4047 & n4050 & (~n363 | n4049);
  assign n4047 = ~x0 & ((~x5 & ~n4048) | (n483 & ~n1511));
  assign n4048 = (x1 | x2 | x3 | x6 | ~x7) & (~x1 | ((x2 | ~x3 | ~x6 | x7) & (~x2 | ~x7 | (x3 ^ x6))));
  assign n4049 = (x2 | ~x5 | (x3 ? (~x6 | x7) : (x6 | ~x7))) & (x5 | ((x6 | x7 | x2 | ~x3) & (~x2 | (x3 ? (x6 | ~x7) : (~x6 | x7)))));
  assign n4050 = n4052 & ~n4054 & ~n4055 & (x2 | n4051);
  assign n4051 = (x0 | x5 | (~x1 ^ x6)) & (~x5 | ((~x0 | (x1 ? (~x3 | x6) : (x3 | ~x6))) & (x0 | x1 | ~x3 | x6)));
  assign n4052 = (n1243 | ~n1268) & (~n387 | (~n4053 & (~n314 | n1243)));
  assign n4053 = x2 & (x3 ? (x5 & ~x6) : (~x5 & x6));
  assign n4054 = ~n506 & ((n483 & n441) | (x0 & ~n791));
  assign n4055 = ~n1402 & ((n340 & n662) | (~x2 & ~n1861));
  assign n4056 = ~n4059 & (~x1 | (~n4058 & (~x4 | n4057)));
  assign n4057 = (~x0 | x2 | x3 | ~x5 | x7) & (x0 | ((~x2 | ~x3 | ~x5 | ~x7) & (x5 | x7 | x2 | x3)));
  assign n4058 = n330 & (x2 ? (~x3 & x5) : (~x5 & (x3 ^ ~x7)));
  assign n4059 = n438 & n403 & (x0 ? (~x4 ^ ~x5) : (~x4 ^ x5));
  assign n4060 = ~x3 & ((n359 & n1422) | (x5 & ~n4061));
  assign n4061 = (~x0 | ~x1 | ~x2 | x4 | ~x7) & (x0 | ~x4 | (x1 ? (~x2 | ~x7) : (x2 | x7)));
  assign n4062 = ~n1279 & n441 & n400;
  assign z221 = n4064 | ~n4068 | (~n542 & ~n4067);
  assign n4064 = x4 & (x0 ? ~n4066 : ~n4065);
  assign n4065 = x1 ? ((~x3 | ~x5 | ~x6) & (x2 | (x3 ? ~x6 : (x5 | x6)))) : ((x2 | ~x3 | x6) & (~x2 | x3 | x5 | ~x6));
  assign n4066 = (x1 | ~x2 | x3 | x5 | ~x6) & (x2 | (x1 ? (x3 ? ~x6 : (x5 | x6)) : (~x3 | x6)));
  assign n4067 = (~x1 | ~x2 | x3 | x4) & (x1 | ((~x4 | ~x5 | x2 | x3) & (~x3 | (x2 ? (~x4 ^ x5) : (x4 | x5)))));
  assign n4068 = ~n4070 & ~n4071 & n4072 & (~x4 | n4069);
  assign n4069 = (~n1658 | ~n921) & (n998 | n1318 | ~n465);
  assign n4070 = (n974 | n2821) & ((~x1 & x6) | (~x0 & x1 & ~x6));
  assign n4071 = n592 & ((n308 & n284) | (~n565 & ~n614));
  assign n4072 = (n565 | n4074) & (~n366 | n4073);
  assign n4073 = (x1 | ~x3 | ~x5 | x6) & (~x1 | ((~x3 | ~x5 | ~x6) & (~x0 | x3 | x6)));
  assign n4074 = (x1 | ~x2 | x3 | x4) & (~x1 | x2 | (x3 ? (x4 | x5) : (~x4 | ~x5)));
  assign z222 = ~n4081 | ~n4077 | (x2 & n363 & ~n4076);
  assign n4076 = (x3 | (x4 ? (~x5 | ~x7) : (x5 | x7))) & (~x3 | x4 | ~x5 | x7);
  assign n4077 = ~n4078 & n4079 & (x7 | ~n324 | n357);
  assign n4078 = ~n453 & (n1037 | (~n736 & ~n470));
  assign n4079 = ~n4080 & (~n647 | ~n2006) & (~n720 | ~n1187);
  assign n4080 = ~x0 & ((~x4 & x7 & ~x2 & ~x3) | (x2 & x3 & x4 & ~x7));
  assign n4081 = x4 ? n4083 : n4082;
  assign n4082 = (~x5 | ~x7 | x2 | ~x3) & (x7 | ((x2 | ~x3 | x5) & (x0 | ~x2 | (x3 ^ x5))));
  assign n4083 = (~n1876 | n4084) & (x3 | ~n2398);
  assign n4084 = x6 ? (~x2 | (x0 & x1)) : x2;
  assign z223 = ~n4090 | n4089 | n4088 | n4086 | n4087;
  assign n4086 = ~x4 & ~n2832;
  assign n4087 = n2569 & (x3 ? (x4 ? (~x5 & ~x6) : x5) : (x4 & (~x5 ^ ~x6)));
  assign n4088 = ~n2755 & ~n487 & x6 & n284;
  assign n4089 = x4 & ~n470 & (x3 ? (~x5 & ~x6) : (~x5 ^ ~x6));
  assign n4090 = (~n300 | ~n606 | ~n328) & (~n270 | ~n2076);
  assign z224 = n4094 | ~n4095 | (~x4 & ~n4092);
  assign n4092 = (~n410 | n4093) & (~n382 | ~n359 | ~n400);
  assign n4093 = x6 & (~x5 | x7);
  assign n4094 = n2569 & (n971 | n1019 | (x5 & n3662));
  assign n4095 = n4096 & n4097 & (n1331 | (~n971 & ~n1019));
  assign n4096 = x0 | ((~n294 | ~n473) & (~n438 | ~n1755));
  assign n4097 = (x1 | ~n327 | n350) & (x0 | ((x1 | n534) & (~n327 | n350)));
  assign z225 = ~n4099 & (~n470 | (n480 & (~x2 | n1383)));
  assign n4099 = ~x5 ^ (x6 & ~x7);
  assign z226 = n4103 | (~n542 & ~n4101);
  assign n4101 = n4102 & (x3 | ((~n424 | ~n359) & n2234));
  assign n4102 = (x0 & x1 & x2) | (~x0 & ~x1 & ~x2 & ~x3);
  assign n4103 = n465 & ((n634 & n742) | (n359 & n633));
  assign z227 = ~x7 & (~n4101 | (n465 & ~n3271));
  assign z228 = n1241 & ~n4106;
  assign n4106 = (~x3 & ~x4 & ~x5 & ~x6 & ~x7) | (x3 & (x4 | (x5 & (x6 | x7))));
  assign z229 = ~x0 & (~n4110 | (n464 & (~n4108 | ~n4109)));
  assign n4108 = (x1 | x2 | x4 | x6 | ~x7) & (~x1 | ~x2 | ~x4 | ~x6 | x7);
  assign n4109 = (~x1 | ~x2 | ~x4 | x6) & (x1 | x2 | x4 | ~x6);
  assign n4110 = (x1 & x2 & x3 & x4 & x5) | (~x1 & ~x2 & (~x3 | ~x4));
  assign z230 = n4113 | n4114 | ~n4116 | (n579 & ~n4112);
  assign n4112 = (~x1 | x3 | ~x4 | x5 | x6) & (x1 | ~x3 | x4 | ~x5 | ~x6);
  assign n4113 = ~x1 & (x2 ? (~x0 | ~x3) : (x0 | (x3 & x4)));
  assign n4114 = ~n4115 & n659 & n786;
  assign n4115 = (~x1 | ~x2 | ~x4 | ~x6) & (x1 | x2 | x4 | x6);
  assign n4116 = (~n387 | ~n974) & (~n394 | ~n1270);
  assign z231 = n4120 | n4122 | ~n4123 | (x5 & ~n4118);
  assign n4118 = (~n1964 | n4119) & (~n308 | ~n443 | ~n359);
  assign n4119 = (x0 | ~x2 | (x1 ? (~x3 | ~x7) : (x3 | x7))) & (~x0 | ~x1 | x2 | x3 | x7);
  assign n4120 = ~x2 & ((n494 & n1063) | (x4 & ~n4121));
  assign n4121 = (x0 | ~x1 | x3 | x5 | ~x6) & (~x0 | x6 | (x1 ? (x3 | ~x5) : (~x3 | x5)));
  assign n4122 = ~x1 & (x0 ? (~x2 ^ (x3 & x4)) : (x2 ? (~x3 & ~x4) : (x3 & x4)));
  assign n4123 = ~n4124 & ~n4125 & ~n4126 & (~n300 | ~n2289);
  assign n4124 = n285 & ((n438 & n425) | (x1 & ~n1012));
  assign n4125 = x0 & ((n725 & n1265) | (n438 & n547));
  assign n4126 = x1 & ~x2 & (x0 ? (~x3 & ~x4) : x3);
  assign z232 = ~n4130 | (x5 & (n4128 | (~n1279 & n1907)));
  assign n4128 = x6 & ((n380 & ~n2563) | (~x3 & ~n4129));
  assign n4129 = x0 ? ((x4 | x7 | x1 | ~x2) & (~x4 | ~x7 | ~x1 | x2)) : (x1 | (x2 ? (~x4 | ~x7) : (x4 | x7)));
  assign n4130 = n4133 & (x2 | (~n4132 & (x5 | n4131)));
  assign n4131 = x0 ? ((~x4 | ~x6 | x1 | ~x3) & (x4 | x6 | ~x1 | x3)) : (x3 | ~x6 | (~x1 ^ ~x4));
  assign n4132 = x5 & n601 & (x1 ? (x3 & ~x6) : (x3 ^ ~x6));
  assign n4133 = n4137 & ~n4136 & ~n4135 & ~n3284 & ~n4134;
  assign n4134 = ~x0 & ((x2 & ~n2345) | (x1 & ~x2 & ~n766));
  assign n4135 = ~x1 & (x0 ? (x2 ? (x3 & x4) : (~x3 & ~x4)) : (x3 & (x2 ^ x4)));
  assign n4136 = x1 & ((x3 & ~x4 & x0 & ~x2) | (~x3 & x4 & ~x0 & x2));
  assign n4137 = (x6 | ~n624 | n4139) & (~x0 | n4138);
  assign n4138 = (~x1 | x2 | ~x3 | ~x4 | x5) & (x1 | (~x2 ^ x4) | (x3 ^ x5));
  assign n4139 = (~x0 | x1 | x3 | ~x5) & (x0 | x5 | (x1 ^ x3));
  assign z233 = n4141 | n4145 | ~n4149 | (n343 & ~n4147);
  assign n4141 = ~x0 & ((n628 & n1755) | n4142 | n4144);
  assign n4142 = ~x1 & (x2 ? (n356 & n875) : ~n4143);
  assign n4143 = (~x3 | ((x4 | ~x5 | x6 | ~x7) & (~x4 | x5 | ~x6 | x7))) & (x3 | x4 | ~x5 | ~x6 | ~x7);
  assign n4144 = ~n1870 & ((x4 & ~x6 & ~x1 & x2) | (x1 & x6 & (~x2 ^ x4)));
  assign n4145 = x3 & ((~x5 & ~n4146) | (n394 & n512));
  assign n4146 = x0 ? (x1 | (x2 ? (~x4 | x6) : (x4 ^ x6))) : ((~x1 | ~x2 | x4 | ~x6) & (~x4 | x6 | x1 | x2));
  assign n4147 = (x3 | n4148) & (~n450 | n1011 | x1 | ~x3);
  assign n4148 = (~x1 | ((~x5 | ~x7 | x2 | ~x4) & (x5 | x7 | ~x2 | x4))) & (x1 | ~x2 | x4 | ~x5 | ~x7);
  assign n4149 = ~n4151 & n4154 & (x5 ? n4150 : n4153);
  assign n4150 = x0 ? (x2 | ((~x1 | x3 | x4) & (~x4 | (x1 & ~x3)))) : ((~x2 | x3 | x4) & (~x1 | (x2 ? x4 : (x3 | ~x4))));
  assign n4151 = ~n753 & ((n366 & n480) | (~x0 & ~n4152));
  assign n4152 = x1 ? (x2 | ~x4) : (~x2 | x4);
  assign n4153 = (x2 | (~x1 ^ ~x3) | (x0 ^ ~x4)) & (x1 | ~x2 | (x0 ? (x3 | ~x4) : (~x3 | x4)));
  assign n4154 = ((~x0 ^ ~x2) | (x4 ? ~n4156 : n4155)) & (~x4 | n4155 | x0 | ~x2) & (~x0 | x2 | x4 | ~n4156);
  assign n4155 = (x1 | ~x3 | ~x5 | ~x6) & (~x1 | x3 | x5 | x6);
  assign n4156 = ~x6 & x5 & ~x1 & ~x3;
  assign z234 = ~n4169 | n4166 | n4158 | n4163;
  assign n4158 = ~x2 & (n4159 | (n730 & ~n4162));
  assign n4159 = ~x5 & ((~x1 & ~n4160) | (n387 & ~n4161));
  assign n4160 = x0 ? ((x6 | x7 | x3 | ~x4) & (~x6 | ~x7 | ~x3 | x4)) : ((x3 | (x4 ? (~x6 | x7) : (x6 | ~x7))) & (~x3 | ~x4 | ~x6 | ~x7));
  assign n4161 = (x3 | x4 | ~x6 | ~x7) & (~x3 | (x4 ? (~x6 | x7) : (x6 | ~x7)));
  assign n4162 = (x1 | ~x3 | ~x4 | ~x6 | x7) & (x4 | ((x1 | ~x3 | x6 | ~x7) & (~x1 | ~x6 | (~x3 ^ ~x7))));
  assign n4163 = n782 & (x3 ? ~n4164 : (~x6 & ~n4165));
  assign n4164 = (x1 | x4 | x5 | ~x6 | x7) & (~x5 | ((x1 | ~x4 | x6 | ~x7) & (~x1 | (x4 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n4165 = (~x1 | x4 | x5 | x7) & (x1 | (x4 ? (x5 | ~x7) : (~x5 | x7)));
  assign n4166 = ~x0 & ((~x2 & ~n4167) | (n3222 & ~n4168));
  assign n4167 = (x1 | ~x3 | ~x4 | ~x5 | x6) & (x4 | (x1 ? (x3 ? (x5 | ~x6) : (~x5 | x6)) : (~x6 | (~x3 ^ ~x5))));
  assign n4168 = (~x1 | ~x3 | x4 | x5) & (x1 | (x3 ? (~x4 | ~x5) : x5));
  assign n4169 = ~n4170 & ~n4172 & n4173 & (~n428 | ~n1259);
  assign n4170 = x1 & ~n4171;
  assign n4171 = (x0 | ~x2 | x3 | x4 | ~x5) & (~x4 | ((x0 | ~x2 | ~x3 | x5) & (~x0 | x2 | (x3 ^ x5))));
  assign n4172 = n363 & ((~x2 & ~x3 & x4 & x5) | (x2 & ~x4 & (x3 ^ ~x5)));
  assign n4173 = n4174 & (n379 | n4153) & (n1909 | n1504);
  assign n4174 = (n583 | n952) & (n1504 | n4175);
  assign n4175 = (~x2 | x5 | ~x6 | ~x7) & (x2 | ~x5 | x6 | x7);
  assign z235 = ~n4182 | n4177 | n4180;
  assign n4177 = ~x0 & ((n269 & n1022) | n4178);
  assign n4178 = ~x7 & (x6 ? ~n4179 : (n282 & ~n989));
  assign n4179 = (~x1 | ~x2 | x3 | ~x4 | ~x5) & (x1 | x2 | (x3 ? (x4 | x5) : (~x4 | ~x5)));
  assign n4180 = ~n542 & (~n4181 | (~n614 & ~n1405));
  assign n4181 = n611 & n1407 & (n420 | n766);
  assign n4182 = n4191 & n4188 & ~n4186 & ~n4183 & ~n4185;
  assign n4183 = ~n4184 & ((n363 & n3141) | (n387 & n1151));
  assign n4184 = (~x3 | ~x4 | ~x5 | ~x6) & (x3 | x4 | x5 | x6);
  assign n4185 = ~n987 & ((n521 & n387) | (n308 & n363));
  assign n4186 = ~n4187 & ((n624 & n327) | (n1207 & n328));
  assign n4187 = (~x0 | ~x1 | x3 | x7) & (x0 | x1 | ~x3 | ~x7);
  assign n4188 = n4189 & n4190 & (n421 | n731);
  assign n4189 = (~n714 | ~n2786) & (~n308 | ~n300 | ~n588);
  assign n4190 = (n405 | n653) & (n481 | n584);
  assign n4191 = ~n4192 & (n614 | n4195) & (~n366 | n4194);
  assign n4192 = ~n377 & ((n428 & n890) | (~n4152 & ~n4193));
  assign n4193 = x0 ? (~x3 | x7) : (x3 | ~x7);
  assign n4194 = (~x6 | x7 | ~x0 | x3) & (x0 | x1 | x6 | ~x7);
  assign n4195 = x3 ? (~n782 | n1897) : (~n308 | ~n364);
  assign z236 = ~n4200 | (x2 & (n4199 | (x3 & ~n4197)));
  assign n4197 = (x1 | n4198) & (x4 | ~n876 | x0 | ~x1);
  assign n4198 = (~x4 | x5 | x6 | ~x7) & (~x0 | x4 | ~x5 | ~x6 | x7);
  assign n4199 = ~n2360 & n363 & ~x3 & ~x4;
  assign n4200 = n4201 & ~n4209 & (n688 | (~n4207 & n4208));
  assign n4201 = ~n4206 & (n1291 | n4203) & (n3778 | n4202);
  assign n4202 = (~x5 | ~x6 | x2 | x3) & (x0 | ~x2 | (x3 ? (~x5 | ~x6) : (x5 | x6)));
  assign n4203 = ~n4204 & ~n4205 & (x3 | n1254 | ~n3691);
  assign n4204 = x1 & ((x2 & ~x3 & ~x4 & x6) | (~x2 & x3 & x4 & ~x6));
  assign n4205 = ~x1 & ((x3 & (x2 ? (~x4 ^ x6) : (~x4 & x6))) | (~x2 & ~x3 & (x4 | ~x6)));
  assign n4206 = ~n377 & ((n394 & n842) | (n423 & ~n3033));
  assign n4207 = n282 & ((n328 & n1064) | (~x0 & n2560));
  assign n4208 = (x1 | ~x2 | x3 | ~x5 | x6) & (x2 | ((x5 | x6 | x1 | ~x3) & (~x1 | ~x6 | (x3 ^ x5))));
  assign n4209 = ~n570 & (x3 ? ~n4211 : ~n4210);
  assign n4210 = (x0 | (x1 ? (~x4 | x6) : (x4 | ~x6))) & (~x1 | x2 | x6) & (x1 | ~x6 | (x2 ^ x4));
  assign n4211 = (x1 | x2 | (x4 ^ x6)) & (x0 | ~x1 | ~x2 | (~x4 ^ x6));
  assign z237 = ~n4215 | ~n4220 | (~x2 & ~n4213);
  assign n4213 = ~n4214 & (~n606 | (~x0 & ~n875) | (x0 & ~n2795));
  assign n4214 = x4 & ((~x6 & ~x7 & ~x3 & ~x5) | (x3 & (x5 ? (~x6 & ~x7) : (x6 & x7))));
  assign n4215 = ~n4219 & (n565 | n4217) & (x4 | n4216);
  assign n4216 = x2 ? (x6 | ((x3 | x5) & (x0 | ~x3 | ~x5))) : (~x6 | (x3 ^ x5));
  assign n4217 = n4218 & (~n278 | ~n363 | (~x3 & ~n465));
  assign n4218 = (x4 | x5 | x2 | ~x3) & (~x2 | ((x3 | x4 | ~x5) & (x0 | ~x4 | (~x3 & x5))));
  assign n4219 = x5 & n356 & ((~x2 & ~x6) | (~x0 & x2 & x6));
  assign n4220 = ~x2 | (x0 ? (x1 | n4222) : n4221);
  assign n4221 = x3 ? ((~x4 | ~x5 | ~x6 | ~x7) & (x5 | ((x6 | x7) & (x4 | ~x6 | ~x7)))) : ((x6 | x7 | x4 | ~x5) & (~x6 | ~x7 | ~x4 | x5));
  assign n4222 = (~x6 | ((~x3 | x4 | x5 | ~x7) & (~x4 | ((~x5 | ~x7) & (x3 | (~x5 & ~x7)))))) & (~x3 | x6 | (x5 ? x4 : x7));
  assign z238 = ~n4227 | (~x6 & (n4224 | n4226));
  assign n4224 = ~x7 & (x4 ? (~n467 & n2569) : ~n4225);
  assign n4225 = (x0 | ~x2 | (x1 ? (~x3 | ~x5) : (x3 | x5))) & (~x0 | ~x1 | x2 | ~x3 | ~x5);
  assign n4226 = n480 & n1151 & (x3 ? (~x4 ^ x5) : (x4 & ~x5));
  assign n4227 = ~n4228 & ~n4230 & n4233 & (n470 | n4232);
  assign n4228 = ~x4 & ((n728 & n876) | (x0 & ~n4229));
  assign n4229 = (x1 | ~x3 | ~x5 | x6 | x7) & (x3 | ((~x1 | (x5 ^ x7)) & (~x5 | ~x6 | ~x7) & (x5 | x6 | x7)));
  assign n4230 = ~n4231 & n480 & n740;
  assign n4231 = x3 ? ((x5 | ~x7) & (x4 | ~x5 | x7)) : (~x4 | (~x5 & x7));
  assign n4232 = (~x3 | x4 | x5 | ~x7) & (x3 | ((~x4 | ~x6 | x7) & (x4 | ~x5 | x6 | ~x7)));
  assign n4233 = (n498 | n470 | n481) & (n542 | n4234);
  assign n4234 = (x1 | ~x4 | (~x3 ^ x5)) & (x0 | (x3 ? (~x4 | x5) : ~x5));
  assign z239 = ~n4242 | (~x7 & (x5 ? ~n4239 : ~n4236));
  assign n4236 = ~n4237 & n4238 & (x3 | n836 | ~n1747);
  assign n4237 = ~x0 & ((~x4 & x6) | (~x1 & x4 & ~x6));
  assign n4238 = (x0 | ~x1 | x2 | ~x4 | x6) & (~x0 | x4 | (x1 & x2) | ~x6);
  assign n4239 = n4240 & (x0 | (~n1964 & (x1 | ~n1019)));
  assign n4240 = n4241 & (~n725 | (x0 ? (~x4 | ~x6) : (x4 | x6)));
  assign n4241 = (x3 | x4 | x6 | ~n514) & (~x4 | ~x6 | ~n363);
  assign n4242 = n4245 & ~n4243 & ~n4244;
  assign n4243 = ~n315 & ((n382 & n910) | (x7 & ~n836));
  assign n4244 = x7 & ~n836 & (n579 | n394);
  assign n4245 = (~n606 | ~n717 | ~n742) & (~n363 | ~n634);
  assign z240 = n4251 | n4250 | n4247 | ~n4248;
  assign n4247 = n725 & ((x5 & ~x7 & (x0 ^ ~x6)) | (x0 & ~x5 & (~x6 | x7)));
  assign n4248 = (x0 | ((x5 | ~x7) & (x1 | ~x5 | x7))) & ~n4249 & (x1 | x5 | ~x7);
  assign n4249 = ~n645 & n328 & ~x7 & n282;
  assign n4250 = ~x7 & ((~x0 & x1 & x5 & x6) | (x0 & ~x1 & (~x5 ^ x6)));
  assign n4251 = n3689 & (x0 ? (n789 | (x6 & n790)) : (~x6 & n790));
  assign z241 = ~n4255 | (~x3 & ((n359 & n634) | n4253));
  assign n4253 = n282 & ((n521 & n329) | (~x4 & ~n4254));
  assign n4254 = x0 ? (x6 ^ ~x7) : (x6 | x7);
  assign n4255 = n4257 & (~n659 | ~n4256) & (~n725 | n4254);
  assign n4256 = ~x7 & (x1 ? (x2 & x6) : (~x2 & ~x6));
  assign n4257 = ~n4259 & n4260 & (n4258 | ~n285 | ~n382);
  assign n4258 = (~x1 | ~x2 | ~x4 | x5) & (x1 | x2 | x4 | ~x5);
  assign n4259 = ~x1 & ((~x6 & x7) | (x0 & x6 & ~x7));
  assign n4260 = x0 | x6 | (x1 ? ~x7 : (~x2 | x7));
  assign z242 = ~n4263 | ~n4265 | (~x3 & ~n4262);
  assign n4262 = (~x0 | ~x1 | ~x2 | x4 | ~x7) & (x0 | ((~x4 | x7 | x1 | x2) & (~x1 | ~x2 | (x4 ^ x7))));
  assign n4263 = n4264 & (~n790 | ~n606 | ~n359);
  assign n4264 = (~x7 & (x0 | (~x1 & ~x2))) | (x1 & x2) | (~x0 & x7);
  assign n4265 = ~n4266 & (~n285 | ~n450 | n4109);
  assign n4266 = ~x0 & x3 & (x1 ? (x2 & x7) : (~x2 & ~x7));
  assign z243 = ~n4269 | n4268 | n3689 | n725 | n1658;
  assign n4268 = ~n1318 & n426 & x4 & n328;
  assign n4269 = (~n971 | ~n1114) & (~n438 | ~n609);
  assign z244 = ~n4271 | (~x6 & ~n478 & n1992);
  assign n4271 = (x2 & (x3 | x4)) | (~x3 & (x4 ? (~x5 & ~x6) : ~x2));
  assign z245 = n4273 | ~n4276 | ~n4278 | (n587 & ~n4275);
  assign n4273 = n328 & ((n359 & n2006) | (x4 & ~n4274));
  assign n4274 = x7 ? (~x3 | (x0 & x1 & x2)) : x3;
  assign n4275 = (x1 | ~x3 | ~x4) & (x0 | ((~x3 | ~x4) & (x1 | x3 | x4)));
  assign n4276 = n4277 & (~n606 | (~x0 & ~x5));
  assign n4277 = (~n300 | ~n606 | ~n328) & (~n387 | ~n613);
  assign n4278 = ~n4279 & (~n284 | ~n659) & (~n363 | ~n612);
  assign n4279 = x4 & n423 & n480 & (x5 | x6);
  assign z246 = ~n4281 & (n410 | ~n470 | n2569);
  assign n4281 = (~x4 & ~x5 & ~x6 & ~x7) | (x4 & (x5 | x6 | x7));
  assign z247 = ~n4284 | ~n4286 | (~n1331 & (n876 | n4283));
  assign n4283 = x5 & (x6 | x7);
  assign n4284 = n4285 & (x7 | ~n328 | (~n410 & ~n1471));
  assign n4285 = (~x0 | ~x1 | x2 | ~n327) & (x0 | x1 | ~n4283);
  assign n4286 = (x3 | n4288) & (x6 | n4287);
  assign n4287 = (x0 | x1 | ~x2 | x5 | x7) & (~x0 | ~x1 | x2 | (x5 ^ x7));
  assign n4288 = (~n359 | ~n411) & (~n624 | ~n480 | ~n4283);
  assign z040 = z037;
  assign z248 = z226;
  assign z249 = z227;
  assign z251 = z250;
  assign z252 = z250;
  assign z253 = z250;
  assign z254 = z250;
  assign z255 = z250;
  assign z256 = z250;
  assign z257 = z250;
endmodule


