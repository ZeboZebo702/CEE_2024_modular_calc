// Benchmark "X_4_64" written by ABC on Thu Jun 22 01:46:37 2023

module X_4_64 ( 
    x0, x1, x2, x3,
    z0, z1, z2, z3, z4, z5, z6, z7, z8, z9  );
  input  x0, x1, x2, x3;
  output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9;
  assign z0 = x0;
  assign z1 = x1;
  assign z2 = x2;
  assign z3 = x3;
  assign z4 = 1'b0;
  assign z5 = 1'b0;
  assign z6 = 1'b0;
  assign z7 = 1'b0;
  assign z8 = 1'b0;
  assign z9 = 1'b0;
endmodule


