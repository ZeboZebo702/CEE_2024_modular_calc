module mult_const_513_bit_mod(
     a,
     r
    );

input [8:1] a;
output [513:1] r;

assign r = (a * 513'd16120775370736350823988927470013450923234256650088346836566427204342423293769121730733856444103918043715008116418812536136346390139704435182750200089763840) % 513'd16353286553968125114719537000830952619242443044080005685170750673635823629736945601850210142816955323191666887328699255407543693843642479920962943360289280;

endmodule