module x_200_mod_4051(
    input [200:1] X,
    output [12:1] R
    );

wire [12:1] r1,r2,r3,r4,r5,r6,r7,r8,r9,r10,r11,r12,r13,r14,r15,r16,r17,r18,r19,r20,
	r21,r22,r23,r24,r25,r26,r27,r28,r29,r30,r31,r32, r33;

X_2 label2 (.x0(X[12]),.x1(X[11]),.x2(X[10]),.x3(X[9]),.x4(X[8]),.x5(X[7]),
.z00(r1[12]),.z01(r1[11]),.z02(r1[10]),.z03(r1[9]),.z04(r1[8]),.z05(r1[7]),.z06(r1[6]),.z07(r1[5]),.z08(r1[4]),.z09(r1[3]),.z10(r1[2]),.z11(r1[1]));

X_3 label3 (.x0(X[18]),.x1(X[17]),.x2(X[16]),.x3(X[15]),.x4(X[14]),.x5(X[13]),
.z00(r2[12]),.z01(r2[11]),.z02(r2[10]),.z03(r2[9]),.z04(r2[8]),.z05(r2[7]),.z06(r2[6]),.z07(r2[5]),.z08(r2[4]),.z09(r2[3]),.z10(r2[2]),.z11(r2[1]));

X_4 label4 (.x0(X[24]),.x1(X[23]),.x2(X[22]),.x3(X[21]),.x4(X[20]),.x5(X[19]),
.z00(r3[12]),.z01(r3[11]),.z02(r3[10]),.z03(r3[9]),.z04(r3[8]),.z05(r3[7]),.z06(r3[6]),.z07(r3[5]),.z08(r3[4]),.z09(r3[3]),.z10(r3[2]),.z11(r3[1]));

X_5 label5 (.x0(X[30]),.x1(X[29]),.x2(X[28]),.x3(X[27]),.x4(X[26]),.x5(X[25]),
.z00(r4[12]),.z01(r4[11]),.z02(r4[10]),.z03(r4[9]),.z04(r4[8]),.z05(r4[7]),.z06(r4[6]),.z07(r4[5]),.z08(r4[4]),.z09(r4[3]),.z10(r4[2]),.z11(r4[1]));

X_6 label6 (.x0(X[36]),.x1(X[35]),.x2(X[34]),.x3(X[33]),.x4(X[32]),.x5(X[31]),
.z00(r5[12]),.z01(r5[11]),.z02(r5[10]),.z03(r5[9]),.z04(r5[8]),.z05(r5[7]),.z06(r5[6]),.z07(r5[5]),.z08(r5[4]),.z09(r5[3]),.z10(r5[2]),.z11(r5[1]));

X_7 label7 (.x0(X[42]),.x1(X[41]),.x2(X[40]),.x3(X[39]),.x4(X[38]),.x5(X[37]),
.z00(r6[12]),.z01(r6[11]),.z02(r6[10]),.z03(r6[9]),.z04(r6[8]),.z05(r6[7]),.z06(r6[6]),.z07(r6[5]),.z08(r6[4]),.z09(r6[3]),.z10(r6[2]),.z11(r6[1]));

X_8 label8 (.x0(X[48]),.x1(X[47]),.x2(X[46]),.x3(X[45]),.x4(X[44]),.x5(X[43]),
.z00(r7[12]),.z01(r7[11]),.z02(r7[10]),.z03(r7[9]),.z04(r7[8]),.z05(r7[7]),.z06(r7[6]),.z07(r7[5]),.z08(r7[4]),.z09(r7[3]),.z10(r7[2]),.z11(r7[1]));

X_9 label9 (.x0(X[54]),.x1(X[53]),.x2(X[52]),.x3(X[51]),.x4(X[50]),.x5(X[49]),
.z00(r8[12]),.z01(r8[11]),.z02(r8[10]),.z03(r8[9]),.z04(r8[8]),.z05(r8[7]),.z06(r8[6]),.z07(r8[5]),.z08(r8[4]),.z09(r8[3]),.z10(r8[2]),.z11(r8[1]));

X_10 label10 (.x0(X[60]),.x1(X[59]),.x2(X[58]),.x3(X[57]),.x4(X[56]),.x5(X[55]),
.z00(r9[12]),.z01(r9[11]),.z02(r9[10]),.z03(r9[9]),.z04(r9[8]),.z05(r9[7]),.z06(r9[6]),.z07(r9[5]),.z08(r9[4]),.z09(r9[3]),.z10(r9[2]),.z11(r9[1]));

X_11 label11 (.x0(X[66]),.x1(X[65]),.x2(X[64]),.x3(X[63]),.x4(X[62]),.x5(X[61]),
.z00(r10[12]),.z01(r10[11]),.z02(r10[10]),.z03(r10[9]),.z04(r10[8]),.z05(r10[7]),.z06(r10[6]),.z07(r10[5]),.z08(r10[4]),.z09(r10[3]),.z10(r10[2]),.z11(r10[1]));

X_12 label12 (.x0(X[72]),.x1(X[71]),.x2(X[70]),.x3(X[69]),.x4(X[68]),.x5(X[67]),
.z00(r11[12]),.z01(r11[11]),.z02(r11[10]),.z03(r11[9]),.z04(r11[8]),.z05(r11[7]),.z06(r11[6]),.z07(r11[5]),.z08(r11[4]),.z09(r11[3]),.z10(r11[2]),.z11(r11[1]));

X_13 label13 (.x0(X[78]),.x1(X[77]),.x2(X[76]),.x3(X[75]),.x4(X[74]),.x5(X[73]),
.z00(r12[12]),.z01(r12[11]),.z02(r12[10]),.z03(r12[9]),.z04(r12[8]),.z05(r12[7]),.z06(r12[6]),.z07(r12[5]),.z08(r12[4]),.z09(r12[3]),.z10(r12[2]),.z11(r12[1]));

X_14 label14 (.x0(X[84]),.x1(X[83]),.x2(X[82]),.x3(X[81]),.x4(X[80]),.x5(X[79]),
.z00(r13[12]),.z01(r13[11]),.z02(r13[10]),.z03(r13[9]),.z04(r13[8]),.z05(r13[7]),.z06(r13[6]),.z07(r13[5]),.z08(r13[4]),.z09(r13[3]),.z10(r13[2]),.z11(r13[1]));

X_15 label15 (.x0(X[90]),.x1(X[89]),.x2(X[88]),.x3(X[87]),.x4(X[86]),.x5(X[85]),
.z00(r14[12]),.z01(r14[11]),.z02(r14[10]),.z03(r14[9]),.z04(r14[8]),.z05(r14[7]),.z06(r14[6]),.z07(r14[5]),.z08(r14[4]),.z09(r14[3]),.z10(r14[2]),.z11(r14[1]));

X_16 label16 (.x0(X[96]),.x1(X[95]),.x2(X[94]),.x3(X[93]),.x4(X[92]),.x5(X[91]),
.z00(r15[12]),.z01(r15[11]),.z02(r15[10]),.z03(r15[9]),.z04(r15[8]),.z05(r15[7]),.z06(r15[6]),.z07(r15[5]),.z08(r15[4]),.z09(r15[3]),.z10(r15[2]),.z11(r15[1]));

X_17 label17 (.x0(X[102]),.x1(X[101]),.x2(X[100]),.x3(X[99]),.x4(X[98]),.x5(X[97]),
.z00(r16[12]),.z01(r16[11]),.z02(r16[10]),.z03(r16[9]),.z04(r16[8]),.z05(r16[7]),.z06(r16[6]),.z07(r16[5]),.z08(r16[4]),.z09(r16[3]),.z10(r16[2]),.z11(r16[1]));

X_18 label18 (.x0(X[108]),.x1(X[107]),.x2(X[106]),.x3(X[105]),.x4(X[104]),.x5(X[103]),
.z00(r17[12]),.z01(r17[11]),.z02(r17[10]),.z03(r17[9]),.z04(r17[8]),.z05(r17[7]),.z06(r17[6]),.z07(r17[5]),.z08(r17[4]),.z09(r17[3]),.z10(r17[2]),.z11(r17[1]));

X_19 label19 (.x0(X[114]),.x1(X[113]),.x2(X[112]),.x3(X[111]),.x4(X[110]),.x5(X[109]),
.z00(r18[12]),.z01(r18[11]),.z02(r18[10]),.z03(r18[9]),.z04(r18[8]),.z05(r18[7]),.z06(r18[6]),.z07(r18[5]),.z08(r18[4]),.z09(r18[3]),.z10(r18[2]),.z11(r18[1]));

X_20 label20 (.x0(X[120]),.x1(X[119]),.x2(X[118]),.x3(X[117]),.x4(X[116]),.x5(X[115]),
.z00(r19[12]),.z01(r19[11]),.z02(r19[10]),.z03(r19[9]),.z04(r19[8]),.z05(r19[7]),.z06(r19[6]),.z07(r19[5]),.z08(r19[4]),.z09(r19[3]),.z10(r19[2]),.z11(r19[1]));

X_21 label21 (.x0(X[126]),.x1(X[125]),.x2(X[124]),.x3(X[123]),.x4(X[122]),.x5(X[121]),
.z00(r20[12]),.z01(r20[11]),.z02(r20[10]),.z03(r20[9]),.z04(r20[8]),.z05(r20[7]),.z06(r20[6]),.z07(r20[5]),.z08(r20[4]),.z09(r20[3]),.z10(r20[2]),.z11(r20[1]));

X_22 label22 (.x0(X[132]),.x1(X[131]),.x2(X[130]),.x3(X[129]),.x4(X[128]),.x5(X[127]),
.z00(r21[12]),.z01(r21[11]),.z02(r21[10]),.z03(r21[9]),.z04(r21[8]),.z05(r21[7]),.z06(r21[6]),.z07(r21[5]),.z08(r21[4]),.z09(r21[3]),.z10(r21[2]),.z11(r21[1]));

X_23 label23 (.x0(X[138]),.x1(X[137]),.x2(X[136]),.x3(X[135]),.x4(X[134]),.x5(X[133]),
.z00(r22[12]),.z01(r22[11]),.z02(r22[10]),.z03(r22[9]),.z04(r22[8]),.z05(r22[7]),.z06(r22[6]),.z07(r22[5]),.z08(r22[4]),.z09(r22[3]),.z10(r22[2]),.z11(r22[1]));

X_24 label24 (.x0(X[144]),.x1(X[143]),.x2(X[142]),.x3(X[141]),.x4(X[140]),.x5(X[139]),
.z00(r23[12]),.z01(r23[11]),.z02(r23[10]),.z03(r23[9]),.z04(r23[8]),.z05(r23[7]),.z06(r23[6]),.z07(r23[5]),.z08(r23[4]),.z09(r23[3]),.z10(r23[2]),.z11(r23[1]));

X_25 label25 (.x0(X[150]),.x1(X[149]),.x2(X[148]),.x3(X[147]),.x4(X[146]),.x5(X[145]),
.z00(r24[12]),.z01(r24[11]),.z02(r24[10]),.z03(r24[9]),.z04(r24[8]),.z05(r24[7]),.z06(r24[6]),.z07(r24[5]),.z08(r24[4]),.z09(r24[3]),.z10(r24[2]),.z11(r24[1]));

X_26 label26 (.x0(X[156]),.x1(X[155]),.x2(X[154]),.x3(X[153]),.x4(X[152]),.x5(X[151]),
.z00(r25[12]),.z01(r25[11]),.z02(r25[10]),.z03(r25[9]),.z04(r25[8]),.z05(r25[7]),.z06(r25[6]),.z07(r25[5]),.z08(r25[4]),.z09(r25[3]),.z10(r25[2]),.z11(r25[1]));

X_27 label27 (.x0(X[162]),.x1(X[161]),.x2(X[160]),.x3(X[159]),.x4(X[158]),.x5(X[157]),
.z00(r26[12]),.z01(r26[11]),.z02(r26[10]),.z03(r26[9]),.z04(r26[8]),.z05(r26[7]),.z06(r26[6]),.z07(r26[5]),.z08(r26[4]),.z09(r26[3]),.z10(r26[2]),.z11(r26[1]));

X_28 label28 (.x0(X[168]),.x1(X[167]),.x2(X[166]),.x3(X[165]),.x4(X[164]),.x5(X[163]),
.z00(r27[12]),.z01(r27[11]),.z02(r27[10]),.z03(r27[9]),.z04(r27[8]),.z05(r27[7]),.z06(r27[6]),.z07(r27[5]),.z08(r27[4]),.z09(r27[3]),.z10(r27[2]),.z11(r27[1]));

X_29 label29 (.x0(X[174]),.x1(X[173]),.x2(X[172]),.x3(X[171]),.x4(X[170]),.x5(X[169]),
.z00(r28[12]),.z01(r28[11]),.z02(r28[10]),.z03(r28[9]),.z04(r28[8]),.z05(r28[7]),.z06(r28[6]),.z07(r28[5]),.z08(r28[4]),.z09(r28[3]),.z10(r28[2]),.z11(r28[1]));

X_30 label30 (.x0(X[180]),.x1(X[179]),.x2(X[178]),.x3(X[177]),.x4(X[176]),.x5(X[175]),
.z00(r29[12]),.z01(r29[11]),.z02(r29[10]),.z03(r29[9]),.z04(r29[8]),.z05(r29[7]),.z06(r29[6]),.z07(r29[5]),.z08(r29[4]),.z09(r29[3]),.z10(r29[2]),.z11(r29[1]));

X_31 label31 (.x0(X[186]),.x1(X[185]),.x2(X[184]),.x3(X[183]),.x4(X[182]),.x5(X[181]),
.z00(r30[12]),.z01(r30[11]),.z02(r30[10]),.z03(r30[9]),.z04(r30[8]),.z05(r30[7]),.z06(r30[6]),.z07(r30[5]),.z08(r30[4]),.z09(r30[3]),.z10(r30[2]),.z11(r30[1]));

X_32 label32 (.x0(X[192]),.x1(X[191]),.x2(X[190]),.x3(X[189]),.x4(X[188]),.x5(X[187]),
.z00(r31[12]),.z01(r31[11]),.z02(r31[10]),.z03(r31[9]),.z04(r31[8]),.z05(r31[7]),.z06(r31[6]),.z07(r31[5]),.z08(r31[4]),.z09(r31[3]),.z10(r31[2]),.z11(r31[1]));

X_33 label33 (.x0(X[198]),.x1(X[197]),.x2(X[196]),.x3(X[195]),.x4(X[194]),.x5(X[193]),
.z00(r32[12]),.z01(r32[11]),.z02(r32[10]),.z03(r32[9]),.z04(r32[8]),.z05(r32[7]),.z06(r32[6]),.z07(r32[5]),.z08(r32[4]),.z09(r32[3]),.z10(r32[2]),.z11(r32[1]));

X_34 label34 (.x0(X[200]),.x1(X[199]),
.z00(r33[12]),.z01(r33[11]),.z02(r33[10]),.z03(r33[9]),.z04(r33[8]),.z05(r33[7]),.z06(r33[6]),.z07(r33[5]),.z08(r33[4]),.z09(r33[3]),.z10(r33[2]),.z11(r33[1]));


wire [14:1] R_temp_1,R_temp_2,R_temp_3,R_temp_4,R_temp_5,R_temp_6,R_temp_7,R_temp_8,R_temp_9,R_temp_10;
wire [13:1] R_temp_11;

assign R_temp_1 = r1 + r2 + r3;
assign R_temp_2 = r4 + r5 + r6;
assign R_temp_3 = r7 + r8 + r9;
assign R_temp_4 = r10 + r11 + r12;
assign R_temp_5 = r13 + r14 + r15;
assign R_temp_6 = r16 + r17 + r18;
assign R_temp_7 = r19 + r20 + r21;
assign R_temp_8 = r22 + r23 + r24;
assign R_temp_9 = r25 + r26 + r27;
assign R_temp_10 =r28  + r29 + r30;
assign R_temp_11 = r31 + r32 + r33;

wire [15:1] R_temp_12,R_temp_13,R_temp_14,R_temp_15;

assign R_temp_12 = R_temp_1 + R_temp_2 + R_temp_3;
assign R_temp_13 = R_temp_4 + R_temp_5 + R_temp_6;
assign R_temp_14 = R_temp_7 + R_temp_8 + R_temp_9;
assign R_temp_15 = R_temp_10 + R_temp_11 + X[6:1];

wire [16:1] R_temp_16,R_temp_17;

assign R_temp_16 = R_temp_12 + R_temp_13;
assign R_temp_17 = R_temp_14 + R_temp_15;

wire [13:1] R_temp_18;

assign R_temp_18 = R_temp_16[6:1] + 64* R_temp_16[12:7] + 45* R_temp_16[16:13] + R_temp_17[6:1] + 64* R_temp_17[12:7] + 45* R_temp_17[16:13];



/// arch_4_6_LUT_add_4_2
/*wire [14:1] R_temp_1,R_temp_2,R_temp_3,R_temp_4,R_temp_5,R_temp_6,R_temp_7,R_temp_8;

assign R_temp_1 = r1 + r2 + r3 + r4;
assign R_temp_2 = r5 + r6 + r7 + r8;
assign R_temp_3 = r9 + r10 + r11 + r12;
assign R_temp_4 = r13 + r14 + r15 + r16;
assign R_temp_5 = r17 + r18 + r19 + r20;
assign R_temp_6 = r21 + r22 + r23 + r24;
assign R_temp_7 = r25 + r26 + r27 + r28;
assign R_temp_8 = r29 + r30 + r31 + r32;

wire [13:1] R_temp_9,R_temp_10,R_temp_11,R_temp_12,R_temp_13,R_temp_14;

assign R_temp_9 = R_temp_1 [6:1] + 64 * R_temp_1 [12:7] + 45 * R_temp_1 [14:13] + R_temp_7 [6:1];
assign R_temp_10 = R_temp_2 [6:1] + 64 * R_temp_2 [12:7] + 45 * R_temp_2 [14:13] + R_temp_8 [6:1];
assign R_temp_11 = R_temp_3 [6:1] + 64 * R_temp_3 [12:7] + 45 * R_temp_3 [14:13] + 64 * R_temp_7 [12:7];
assign R_temp_12 = R_temp_4 [6:1] + 64 * R_temp_4 [12:7] + 45 * R_temp_4 [14:13] + 64 * R_temp_8 [12:7];
assign R_temp_13 = R_temp_5 [6:1] + 64 * R_temp_5 [12:7] + 45 * R_temp_5 [14:13] + 45 * R_temp_7 [14:13];
assign R_temp_14 = R_temp_6 [6:1] + 64 * R_temp_1 [12:7] + 45 * R_temp_6 [14:13] + 45 * R_temp_8 [14:13];

wire [13:1] R_temp_15,R_temp_16,R_temp_17,R_temp_18;
//wire [12:1] R_temp_19;

assign R_temp_15 = R_temp_9 [6:1] + 64 * R_temp_9 [12:7] + 45 * R_temp_9 [13] + X [6:1];
assign R_temp_16 = R_temp_10 [6:1] + 64 * R_temp_10 [12:7] + 45 * R_temp_10 [13] + R_temp_14 [6:1];
assign R_temp_17 = R_temp_11 [6:1] + 64 * R_temp_11 [12:7] + 45 * R_temp_11 [13] + 64 * R_temp_14 [12:7];
assign R_temp_18 = R_temp_12 [6:1] + 64 * R_temp_12 [12:7] + 45 * R_temp_12 [13] + 45 * R_temp_14 [13];
//assign R_temp_19 = R_temp_13 [6:1] + 64 * R_temp_13 [12:7] + 45 * R_temp_13 [13];

wire [13:1] R_temp_20,R_temp_21,R_temp_22,R_temp_23;

assign R_temp_20 = R_temp_15 [6:1] + 64 * R_temp_15 [12:7] + 45 * R_temp_15 [13] + R_temp_18 [6:1];
assign R_temp_21 = R_temp_16 [6:1] + 64 * R_temp_16 [12:7] + 45 * R_temp_16 [13] + 64 * R_temp_18 [12:7] ;
assign R_temp_22 = R_temp_17 [6:1] + 64 * R_temp_17 [12:7] + 45 * R_temp_17 [13] + 64 * R_temp_13 [12:7];
assign R_temp_23 = r33[6:1] + 64 * r33 [12:7] + R_temp_13 [6:1] + 45 * R_temp_18 [13] + R_temp_13 [13];

wire [13:1] R_temp_24,R_temp_25,R_temp_26;

assign R_temp_24 = R_temp_20 [6:1] + 64 * R_temp_21 [12:7] + 45 * R_temp_20 [13] + R_temp_23 [6:1];
assign R_temp_25 = R_temp_21 [6:1] + 64 * R_temp_21 [12:7] + 45 * R_temp_21 [13] + 64 * R_temp_23 [12:7];
assign R_temp_26 = R_temp_22 [6:1] + 64 * R_temp_22 [12:7] + 45 * R_temp_22 [13] + 45 * R_temp_23 [13];

wire [13:1] R_temp_27, R_temp_28;

assign R_temp_27 = R_temp_24 [6:1] + 64 * R_temp_24 [12:7] + 45 * R_temp_24 [13] + R_temp_26 [6:1] + 45 * R_temp_26 [13];
assign R_temp_28 = R_temp_25 [6:1] + 64 * R_temp_25 [12:7] + 45 * R_temp_25 [13] + 64 * R_temp_26 [12:7];

wire [13:1] R_temp_29;

assign R_temp_29 = R_temp_27 + R_temp_28;*/

reg [12:1]  R_temp;

always @(R_temp_18)
begin
  if (R_temp_18 >= 12'b111111010011  )
    R_temp <= R_temp_18 - 12'b111111010011;
  else
    R_temp <= R_temp_18;
end

assign R = R_temp;

endmodule
