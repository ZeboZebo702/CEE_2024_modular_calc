// Benchmark "256_256_mod" written by ABC on Thu Dec 01 02:21:46 2022

module const_256_256_mod ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z000, z001, z002, z003, z004, z005, z006, z007, z008, z009, z010, z011,
    z012, z013, z014, z015, z016, z017, z018, z019, z020, z021, z022, z023,
    z024, z025, z026, z027, z028, z029, z030, z031, z032, z033, z034, z035,
    z036, z037, z038, z039, z040, z041, z042, z043, z044, z045, z046, z047,
    z048, z049, z050, z051, z052, z053, z054, z055, z056, z057, z058, z059,
    z060, z061, z062, z063, z064, z065, z066, z067, z068, z069, z070, z071,
    z072, z073, z074, z075, z076, z077, z078, z079, z080, z081, z082, z083,
    z084, z085, z086, z087, z088, z089, z090, z091, z092, z093, z094, z095,
    z096, z097, z098, z099, z100, z101, z102, z103, z104, z105, z106, z107,
    z108, z109, z110, z111, z112, z113, z114, z115, z116, z117, z118, z119,
    z120, z121, z122, z123, z124, z125, z126, z127, z128, z129, z130, z131,
    z132, z133, z134, z135, z136, z137, z138, z139, z140, z141, z142, z143,
    z144, z145, z146, z147, z148, z149, z150, z151, z152, z153, z154, z155,
    z156, z157, z158, z159, z160, z161, z162, z163, z164, z165, z166, z167,
    z168, z169, z170, z171, z172, z173, z174, z175, z176, z177, z178, z179,
    z180, z181, z182, z183, z184, z185, z186, z187, z188, z189, z190, z191,
    z192, z193, z194, z195, z196, z197, z198, z199, z200, z201, z202, z203,
    z204, z205, z206, z207, z208, z209, z210, z211, z212, z213, z214, z215,
    z216, z217, z218, z219, z220, z221, z222, z223, z224, z225, z226, z227,
    z228, z229, z230, z231, z232, z233, z234, z235, z236, z237, z238, z239,
    z240, z241, z242, z243, z244, z245, z246, z247, z248, z249, z250, z251,
    z252, z253, z254, z255, z256, z257, z258, z259, z260, z261, z262, z263,
    z264, z265, z266, z267, z268, z269, z270, z271, z272, z273, z274, z275,
    z276, z277, z278, z279, z280, z281, z282, z283, z284, z285, z286, z287,
    z288, z289, z290, z291, z292, z293, z294, z295, z296, z297, z298, z299,
    z300, z301, z302, z303, z304, z305, z306, z307, z308, z309, z310, z311,
    z312, z313, z314, z315, z316, z317, z318, z319, z320, z321, z322, z323,
    z324, z325, z326, z327, z328, z329, z330, z331, z332, z333, z334, z335,
    z336, z337, z338, z339, z340, z341, z342, z343, z344, z345, z346, z347,
    z348, z349, z350, z351, z352, z353, z354, z355, z356, z357, z358, z359,
    z360, z361, z362, z363, z364, z365, z366, z367, z368, z369, z370, z371,
    z372, z373, z374, z375, z376, z377, z378, z379, z380, z381, z382, z383,
    z384, z385, z386, z387, z388, z389, z390, z391, z392, z393, z394, z395,
    z396, z397, z398, z399, z400, z401, z402, z403, z404, z405, z406, z407,
    z408, z409, z410, z411, z412, z413, z414, z415, z416, z417, z418, z419,
    z420, z421, z422, z423, z424, z425, z426, z427, z428, z429, z430, z431,
    z432, z433, z434, z435, z436, z437, z438, z439, z440, z441, z442, z443,
    z444, z445, z446, z447, z448, z449, z450, z451, z452, z453, z454, z455,
    z456, z457, z458, z459, z460, z461, z462, z463, z464, z465, z466, z467,
    z468, z469, z470, z471, z472, z473, z474, z475, z476, z477, z478, z479,
    z480, z481, z482, z483, z484, z485, z486, z487, z488, z489, z490, z491,
    z492, z493, z494, z495, z496, z497, z498, z499, z500, z501, z502, z503,
    z504, z505, z506, z507, z508, z509, z510, z511, z512  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z000, z001, z002, z003, z004, z005, z006, z007, z008, z009, z010,
    z011, z012, z013, z014, z015, z016, z017, z018, z019, z020, z021, z022,
    z023, z024, z025, z026, z027, z028, z029, z030, z031, z032, z033, z034,
    z035, z036, z037, z038, z039, z040, z041, z042, z043, z044, z045, z046,
    z047, z048, z049, z050, z051, z052, z053, z054, z055, z056, z057, z058,
    z059, z060, z061, z062, z063, z064, z065, z066, z067, z068, z069, z070,
    z071, z072, z073, z074, z075, z076, z077, z078, z079, z080, z081, z082,
    z083, z084, z085, z086, z087, z088, z089, z090, z091, z092, z093, z094,
    z095, z096, z097, z098, z099, z100, z101, z102, z103, z104, z105, z106,
    z107, z108, z109, z110, z111, z112, z113, z114, z115, z116, z117, z118,
    z119, z120, z121, z122, z123, z124, z125, z126, z127, z128, z129, z130,
    z131, z132, z133, z134, z135, z136, z137, z138, z139, z140, z141, z142,
    z143, z144, z145, z146, z147, z148, z149, z150, z151, z152, z153, z154,
    z155, z156, z157, z158, z159, z160, z161, z162, z163, z164, z165, z166,
    z167, z168, z169, z170, z171, z172, z173, z174, z175, z176, z177, z178,
    z179, z180, z181, z182, z183, z184, z185, z186, z187, z188, z189, z190,
    z191, z192, z193, z194, z195, z196, z197, z198, z199, z200, z201, z202,
    z203, z204, z205, z206, z207, z208, z209, z210, z211, z212, z213, z214,
    z215, z216, z217, z218, z219, z220, z221, z222, z223, z224, z225, z226,
    z227, z228, z229, z230, z231, z232, z233, z234, z235, z236, z237, z238,
    z239, z240, z241, z242, z243, z244, z245, z246, z247, z248, z249, z250,
    z251, z252, z253, z254, z255, z256, z257, z258, z259, z260, z261, z262,
    z263, z264, z265, z266, z267, z268, z269, z270, z271, z272, z273, z274,
    z275, z276, z277, z278, z279, z280, z281, z282, z283, z284, z285, z286,
    z287, z288, z289, z290, z291, z292, z293, z294, z295, z296, z297, z298,
    z299, z300, z301, z302, z303, z304, z305, z306, z307, z308, z309, z310,
    z311, z312, z313, z314, z315, z316, z317, z318, z319, z320, z321, z322,
    z323, z324, z325, z326, z327, z328, z329, z330, z331, z332, z333, z334,
    z335, z336, z337, z338, z339, z340, z341, z342, z343, z344, z345, z346,
    z347, z348, z349, z350, z351, z352, z353, z354, z355, z356, z357, z358,
    z359, z360, z361, z362, z363, z364, z365, z366, z367, z368, z369, z370,
    z371, z372, z373, z374, z375, z376, z377, z378, z379, z380, z381, z382,
    z383, z384, z385, z386, z387, z388, z389, z390, z391, z392, z393, z394,
    z395, z396, z397, z398, z399, z400, z401, z402, z403, z404, z405, z406,
    z407, z408, z409, z410, z411, z412, z413, z414, z415, z416, z417, z418,
    z419, z420, z421, z422, z423, z424, z425, z426, z427, z428, z429, z430,
    z431, z432, z433, z434, z435, z436, z437, z438, z439, z440, z441, z442,
    z443, z444, z445, z446, z447, z448, z449, z450, z451, z452, z453, z454,
    z455, z456, z457, z458, z459, z460, z461, z462, z463, z464, z465, z466,
    z467, z468, z469, z470, z471, z472, z473, z474, z475, z476, z477, z478,
    z479, z480, z481, z482, z483, z484, z485, z486, z487, z488, z489, z490,
    z491, z492, z493, z494, z495, z496, z497, z498, z499, z500, z501, z502,
    z503, z504, z505, z506, z507, z508, z509, z510, z511, z512;
  wire n523, n524, n526, n527, n528, n529, n531, n532, n533, n534, n535,
    n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n561,
    n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
    n574, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
    n613, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n637, n638,
    n639, n640, n641, n642, n643, n644, n645, n646, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671, n672, n673, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684, n685, n686, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697, n698, n699, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n727, n728, n729,
    n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n741, n742,
    n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
    n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
    n768, n769, n770, n771, n772, n774, n775, n776, n777, n778, n780, n781,
    n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
    n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
    n807, n808, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
    n820, n821, n822, n824, n825, n826, n827, n828, n829, n830, n831, n832,
    n833, n834, n835, n836, n837, n838, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n863, n864, n865, n866, n867, n868, n869, n870, n871,
    n872, n873, n874, n875, n876, n877, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891, n892, n894, n895, n896, n897,
    n898, n899, n900, n901, n902, n903, n904, n906, n907, n908, n909, n910,
    n911, n912, n913, n914, n915, n916, n917, n918, n919, n921, n922, n923,
    n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n935, n936,
    n937, n938, n939, n940, n942, n943, n944, n945, n946, n947, n949, n950,
    n951, n952, n953, n955, n956, n957, n958, n959, n960, n961, n963, n964,
    n965, n966, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
    n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n991,
    n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
    n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1023, n1024,
    n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
    n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
    n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
    n1079, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1110, n1111,
    n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
    n1122, n1123, n1124, n1125, n1127, n1128, n1129, n1130, n1131, n1132,
    n1134, n1135, n1136, n1137, n1139, n1140, n1141, n1142, n1144, n1145,
    n1148, n1149, n1150, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
    n1159, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1170,
    n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
    n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1192,
    n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
    n1214, n1215, n1216, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1233, n1234, n1235,
    n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
    n1268, n1269, n1270, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
    n1279, n1280, n1281, n1282, n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1299, n1300,
    n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1316, n1317, n1318, n1319, n1320, n1321,
    n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1330, n1331, n1332,
    n1333, n1334, n1335, n1336, n1338, n1339, n1340, n1341, n1342, n1343,
    n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1353, n1354,
    n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
    n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1397,
    n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1435, n1436, n1437, n1438, n1439, n1440,
    n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
    n1452, n1453, n1454, n1455, n1456, n1458, n1459, n1460, n1461, n1462,
    n1463, n1464, n1465, n1466, n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1483, n1484,
    n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1493, n1494, n1495,
    n1496, n1497, n1498, n1499, n1500, n1501, n1503, n1504, n1505, n1506,
    n1507, n1508, n1509, n1510, n1511, n1513, n1514, n1515, n1516, n1517,
    n1518, n1519, n1520, n1521, n1522, n1524, n1525, n1526, n1527, n1528,
    n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
    n1572, n1573, n1574, n1575, n1577, n1578, n1579, n1580, n1581, n1582,
    n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
    n1593, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609, n1611, n1612, n1613, n1614,
    n1615, n1616, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
    n1626, n1627, n1628, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
    n1637, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
    n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
    n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
    n1681, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
    n1692, n1693, n1694, n1695, n1696, n1698, n1699, n1700, n1701, n1702,
    n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1723, n1724,
    n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1733, n1734, n1735,
    n1736, n1737, n1738, n1739, n1740, n1741, n1743, n1744, n1745, n1746,
    n1747, n1748, n1749, n1750, n1751, n1752, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1764, n1765, n1766, n1767, n1768,
    n1769, n1770, n1771, n1772, n1773, n1774, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1802,
    n1803, n1804, n1805, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
    n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1823, n1824, n1825,
    n1826, n1827, n1828, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
    n1837, n1838, n1839, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
    n1848, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1859,
    n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1870,
    n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1892,
    n1893, n1894, n1895, n1896, n1897, n1898, n1900, n1901, n1902, n1903,
    n1904, n1905, n1906, n1908, n1909, n1910, n1911, n1913, n1914, n1915,
    n1916, n1917, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1927,
    n1928, n1929, n1930, n1931, n1933, n1934, n1935, n1936, n1937, n1938,
    n1939, n1940, n1941, n1942, n1943, n1945, n1946, n1947, n1948, n1949,
    n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1960,
    n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1970, n1971,
    n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1981, n1982,
    n1983, n1984, n1985, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
    n1994, n1995, n1996, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
    n2005, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
    n2016, n2017, n2018, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
    n2027, n2028, n2029, n2030, n2032, n2033, n2034, n2035, n2036, n2037,
    n2038, n2039, n2040, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
    n2049, n2050, n2051, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2073, n2074, n2075, n2077, n2078, n2080, n2081, n2082, n2083,
    n2084, n2085, n2086, n2087, n2089, n2090, n2091, n2092, n2093, n2094,
    n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2104, n2105,
    n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2116,
    n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
    n2127, n2128, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
    n2138, n2140, n2141, n2142, n2143, n2144, n2145, n2147, n2148, n2149,
    n2150, n2151, n2152, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
    n2161, n2162, n2163, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
    n2172, n2173, n2174, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
    n2183, n2184, n2185, n2186, n2188, n2189, n2190, n2191, n2192, n2193,
    n2194, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
    n2205, n2206, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
    n2216, n2217, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
    n2227, n2228, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
    n2238, n2239, n2240, n2241, n2242, n2243, n2245, n2246, n2247, n2248,
    n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2269, n2270,
    n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
    n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
    n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2300, n2301, n2302,
    n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2313,
    n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
    n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2334,
    n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2344, n2345,
    n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
    n2367, n2368, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
    n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2389,
    n2390, n2391, n2392, n2393, n2394, n2395, n2397, n2398, n2399, n2400,
    n2401, n2402, n2403, n2404, n2405, n2407, n2408, n2409, n2410, n2411,
    n2412, n2413, n2414, n2415, n2416, n2417, n2419, n2420, n2421, n2422,
    n2423, n2424, n2425, n2426, n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2436, n2437, n2438, n2439, n2440, n2441, n2443, n2444, n2445,
    n2446, n2447, n2448, n2450, n2451, n2452, n2453, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2463, n2464, n2465, n2466, n2467, n2468,
    n2469, n2470, n2471, n2472, n2473, n2475, n2476, n2477, n2478, n2479,
    n2480, n2481, n2482, n2483, n2484, n2485, n2487, n2488, n2489, n2490,
    n2491, n2492, n2493, n2494, n2495, n2497, n2498, n2499, n2500, n2501,
    n2502, n2503, n2504, n2505, n2507, n2508, n2509, n2510, n2511, n2512,
    n2513, n2514, n2515, n2516, n2517, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2529, n2530, n2531, n2532, n2533, n2534,
    n2535, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2546,
    n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
    n2557, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
    n2568, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
    n2579, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
    n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
    n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2611, n2612,
    n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2621, n2622, n2623,
    n2624, n2625, n2626, n2627, n2628, n2629, n2631, n2632, n2633, n2634,
    n2635, n2636, n2637, n2638, n2639, n2640, n2642, n2643, n2644, n2645,
    n2646, n2647, n2648, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
    n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2665, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2688, n2689,
    n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2699, n2700,
    n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2711,
    n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2721, n2722,
    n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
    n2733, n2734, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
    n2744, n2745, n2746, n2747, n2748, n2750, n2751, n2752, n2753, n2754,
    n2755, n2756, n2757, n2758, n2759, n2760, n2762, n2763, n2764, n2765,
    n2766, n2767, n2768, n2769, n2770, n2771, n2773, n2774, n2775, n2776,
    n2777, n2778, n2779, n2780, n2781, n2783, n2784, n2785, n2786, n2787,
    n2788, n2789, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
    n2799, n2800, n2801, n2802, n2804, n2805, n2806, n2807, n2808, n2809,
    n2810, n2811, n2812, n2813, n2815, n2816, n2817, n2818, n2819, n2820,
    n2821, n2822, n2823, n2824, n2825, n2826, n2828, n2829, n2830, n2831,
    n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2841, n2842,
    n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2862, n2863, n2864,
    n2865, n2866, n2867, n2868, n2869, n2871, n2872, n2873, n2874, n2875,
    n2876, n2877, n2878, n2879, n2881, n2882, n2883, n2884, n2885, n2886,
    n2887, n2888, n2889, n2890, n2892, n2893, n2894, n2895, n2896, n2897,
    n2898, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2909,
    n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2919, n2920,
    n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2930, n2931,
    n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2941, n2942,
    n2943, n2944, n2945, n2946, n2947, n2948, n2950, n2951, n2952, n2953,
    n2954, n2955, n2956, n2957, n2958, n2959, n2961, n2963, n2964, n2965,
    n2966, n2967, n2968, n2970, n2971, n2973, n2974, n2975, n2976, n2977,
    n2978, n2980, n2981, n2984, n2985, n2986, n2988, n2989, n2991, n2992,
    n2993, n2994, n2995, n2997, n2998, n2999, n3000, n3001, n3002, n3004,
    n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
    n3015, n3016, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
    n3026, n3027, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
    n3037, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
    n3048, n3049, n3050, n3051, n3053, n3054, n3055, n3056, n3057, n3058,
    n3059, n3060, n3061, n3062, n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075, n3077, n3078, n3079, n3080,
    n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3089, n3090, n3091,
    n3092, n3093, n3094, n3095, n3097, n3098, n3099, n3100, n3101, n3102,
    n3103, n3105, n3106, n3107, n3109, n3110, n3111, n3112, n3114, n3115,
    n3116, n3118, n3119, n3120, n3121, n3122, n3123, n3125, n3126, n3127,
    n3128, n3129, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3139,
    n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
    n3150, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3161,
    n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
    n3172, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
    n3183, n3184, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
    n3194, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3204, n3205,
    n3206, n3207, n3208, n3209, n3210, n3212, n3213, n3214, n3215, n3216,
    n3217, n3218, n3219, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
    n3228, n3229, n3230, n3231, n3233, n3234, n3235, n3236, n3237, n3238,
    n3239, n3240, n3241, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
    n3250, n3251, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
    n3261, n3262, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
    n3272, n3273, n3274, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
    n3283, n3284, n3285, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
    n3294, n3295, n3296, n3297, n3299, n3300, n3301, n3302, n3303, n3304,
    n3305, n3306, n3307, n3309, n3310, n3311, n3312, n3313, n3314, n3316,
    n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
    n3328, n3329, n3330, n3331, n3332, n3334, n3335, n3336, n3337, n3338,
    n3340, n3341, n3342, n3343, n3345, n3346, n3347, n3349, n3350, n3351,
    n3352, n3354, n3355, n3356, n3357, n3358, n3360, n3361, n3362, n3363,
    n3364, n3365, n3366, n3367, n3368, n3369, n3371, n3372, n3373, n3374,
    n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3385,
    n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
    n3396, n3397, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
    n3407, n3408, n3409, n3410, n3412, n3413, n3414, n3415, n3416, n3417,
    n3418, n3419, n3420, n3421, n3423, n3424, n3425, n3426, n3427, n3428,
    n3429, n3430, n3431, n3432, n3433, n3434, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3450,
    n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
    n3461, n3462, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
    n3472, n3473, n3474, n3475, n3477, n3478, n3479, n3480, n3481, n3482,
    n3483, n3484, n3485, n3486, n3487, n3488, n3490, n3491, n3492, n3493,
    n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3504,
    n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3514, n3515,
    n3516, n3517, n3518, n3519, n3520, n3522, n3523, n3524, n3525, n3526,
    n3527, n3528, n3529, n3530, n3532, n3533, n3534, n3535, n3536, n3537,
    n3538, n3539, n3540, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
    n3560, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
    n3571, n3572, n3573, n3574, n3575, n3577, n3578, n3579, n3580, n3581,
    n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3591, n3592,
    n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3603,
    n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
    n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
    n3625, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
    n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
    n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3657, n3658,
    n3659, n3660, n3661, n3662, n3663, n3664, n3666, n3667, n3668, n3669,
    n3670, n3671, n3672, n3673, n3674, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3686, n3687, n3688, n3689, n3690, n3691,
    n3692, n3693, n3694, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
    n3703, n3704, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
    n3715, n3716, n3717, n3718, n3719, n3720, n3722, n3723, n3724, n3725,
    n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3735, n3736,
    n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3745, n3746, n3747,
    n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3757, n3758,
    n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3767, n3768, n3769,
    n3770, n3771, n3772, n3773, n3774, n3775, n3777, n3778, n3779, n3780,
    n3781, n3782, n3783, n3784, n3785, n3786, n3788, n3789, n3790, n3791,
    n3792, n3793, n3794, n3796, n3797, n3798, n3799, n3800, n3801, n3803,
    n3804, n3805, n3806, n3808, n3809, n3810, n3812, n3813, n3814, n3816,
    n3817, n3818, n3819, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
    n3828, n3830, n3831, n3832, n3833, n3834, n3835, n3837, n3838, n3839,
    n3840, n3841, n3842, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
    n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3861, n3862,
    n3863, n3864, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3874,
    n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3884, n3885,
    n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
    n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3907,
    n3908, n3909, n3910, n3911, n3912, n3913, n3915, n3916, n3917, n3918,
    n3919, n3920, n3921, n3922, n3924, n3925, n3926, n3927, n3928, n3929,
    n3930, n3931, n3932, n3933, n3935, n3936, n3937, n3938, n3939, n3940,
    n3941, n3942, n3943, n3944, n3945, n3947, n3948, n3949, n3950, n3951,
    n3952, n3953, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
    n3963, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3974,
    n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3983, n3984, n3985,
    n3986, n3987, n3988, n3989, n3990, n3992, n3993, n3994, n3996, n3997,
    n3998, n3999, n4000, n4002, n4003, n4004, n4005, n4006, n4008, n4009,
    n4010, n4011, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
    n4022, n4023, n4024, n4025, n4026, n4027, n4029, n4030, n4031, n4032,
    n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4041, n4042, n4043,
    n4044, n4045, n4046, n4047, n4048, n4050, n4051, n4052, n4053, n4054,
    n4055, n4056, n4057, n4058, n4059, n4061, n4062, n4063, n4064, n4065,
    n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4074, n4075, n4076,
    n4077, n4078, n4079, n4080, n4082, n4083, n4084, n4085, n4086, n4087,
    n4088, n4089, n4090, n4091, n4093, n4094, n4095, n4096, n4097, n4098,
    n4099, n4100, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
    n4110, n4111, n4112, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
    n4121, n4122, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
    n4132, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
    n4143, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
    n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4165,
    n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4175, n4176,
    n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4185, n4186, n4187,
    n4188, n4189, n4190, n4191, n4193, n4194, n4195, n4196, n4197, n4198,
    n4199, n4200, n4201, n4202, n4204, n4205, n4206, n4207, n4208, n4209,
    n4210, n4211, n4212, n4213, n4214, n4216, n4217, n4218, n4219, n4220,
    n4221, n4222, n4223, n4224, n4225, n4227, n4228, n4229, n4230, n4231,
    n4232, n4234, n4235, n4236, n4237, n4239, n4240, n4241, n4242, n4243,
    n4244, n4245, n4246, n4247, n4249, n4250, n4251, n4252, n4253, n4254,
    n4255, n4256, n4258, n4259, n4260, n4261, n4262, n4263, n4265, n4266,
    n4267, n4269, n4270, n4271, n4272, n4273, n4274, n4276, n4277, n4278,
    n4279, n4280, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
    n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4299, n4300, n4301,
    n4302, n4303, n4304, n4305, n4307, n4308, n4309, n4310, n4311, n4312,
    n4313, n4314, n4315, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
    n4324, n4325, n4326, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
    n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
    n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4357,
    n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
    n4368, n4369, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4379,
    n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4389, n4390,
    n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4400, n4401,
    n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4410, n4411, n4412,
    n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4422, n4423,
    n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4433, n4434,
    n4435, n4436, n4437, n4438, n4439, n4440, n4442, n4443, n4444, n4445,
    n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4455, n4456,
    n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4465, n4466, n4467,
    n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4478,
    n4479, n4481, n4482, n4483, n4484, n4485, n4486, n4488, n4489, n4490,
    n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4501,
    n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4510, n4511, n4512,
    n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
    n4523, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
    n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4545,
    n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4555, n4556,
    n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
    n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
    n4578, n4580, n4581, n4582, n4583, n4584, n4585, n4587, n4588, n4589,
    n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4598, n4599, n4600,
    n4601, n4602, n4603, n4604, n4605, n4606, n4608, n4609, n4610, n4611,
    n4612, n4613, n4614, n4615, n4616, n4617, n4619, n4620, n4621, n4622,
    n4623, n4624, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
    n4635, n4636, n4637, n4638, n4639, n4640, n4642, n4643, n4644, n4645,
    n4647, n4648, n4649, n4650, n4651, n4653, n4654, n4655, n4658, n4659,
    n4660, n4662, n4663, n4664, n4666, n4667, n4668, n4669, n4671, n4672,
    n4673, n4674, n4675, n4676, n4677, n4679, n4680, n4681, n4682, n4684,
    n4685, n4686, n4688, n4689, n4690, n4691, n4692, n4694, n4695, n4696,
    n4698, n4699, n4700, n4701, n4702, n4704, n4705, n4706, n4707, n4708,
    n4709, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4720,
    n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
    n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4742,
    n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4753,
    n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
    n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4773, n4774, n4775,
    n4776, n4777, n4778, n4779, n4780, n4783, n4784, n4785, n4786, n4788,
    n4789, n4790, n4791, n4792, n4793, n4794, n4796, n4797, n4798, n4799,
    n4800, n4801, n4802, n4803, n4804, n4806, n4807, n4808, n4810, n4811,
    n4812, n4813, n4814, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
    n4823, n4824, n4825, n4826, n4827, n4829, n4830, n4831, n4832, n4833,
    n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4843, n4844,
    n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4853, n4854, n4855,
    n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4864, n4865, n4866,
    n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4875, n4876, n4877,
    n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4886, n4887, n4888,
    n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4898, n4899,
    n4900, n4901, n4902, n4903, n4904, n4905, n4907, n4908, n4909, n4910,
    n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4919, n4920, n4921,
    n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4931, n4932,
    n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
    n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
    n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
    n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4973, n4974, n4975,
    n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4985, n4986,
    n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4997,
    n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5007, n5008,
    n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5017, n5018, n5019,
    n5020, n5021, n5022, n5023, n5025, n5026, n5027, n5028, n5029, n5030,
    n5031, n5032, n5033, n5034, n5036, n5037, n5038, n5039, n5040, n5041,
    n5042, n5043, n5044, n5045, n5046, n5048, n5049, n5050, n5051, n5052,
    n5053, n5054, n5055, n5056, n5058, n5059, n5060, n5061, n5062, n5063,
    n5064, n5065, n5066, n5067, n5068, n5070, n5071, n5072, n5073, n5074,
    n5075, n5076, n5077, n5078, n5080, n5081, n5082, n5083, n5084, n5085,
    n5086, n5087, n5088, n5089, n5091, n5092, n5093, n5094, n5095, n5096,
    n5097, n5098, n5099, n5100, n5101, n5103, n5104, n5105, n5106, n5107,
    n5108, n5109, n5110, n5111, n5112, n5114, n5115, n5116, n5117, n5118,
    n5119, n5120, n5121, n5122, n5123, n5125, n5126, n5127, n5128, n5129,
    n5130, n5131, n5132, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
    n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
    n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5162, n5163,
    n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5174,
    n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
    n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5196,
    n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5205, n5206, n5207,
    n5208, n5209, n5210, n5211, n5212, n5213, n5215, n5216, n5217, n5218,
    n5219, n5220, n5221, n5222, n5224, n5225, n5226, n5227, n5228, n5229,
    n5230, n5231, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5241,
    n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5251, n5252,
    n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
    n5263, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5274,
    n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
    n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5296,
    n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5305, n5306, n5307,
    n5308, n5309, n5310, n5311, n5312, n5314, n5315, n5316, n5317, n5318,
    n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
    n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5340, n5341,
    n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5350, n5351, n5352,
    n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5361, n5362, n5363,
    n5364, n5365, n5366, n5367, n5368, n5369, n5371, n5372, n5373, n5374,
    n5375, n5376, n5377, n5378, n5379, n5381, n5382, n5383, n5384, n5385,
    n5386, n5387, n5388, n5389, n5390, n5391, n5393, n5394, n5395, n5396,
    n5397, n5398, n5399, n5400, n5401, n5403, n5404, n5405, n5406, n5407,
    n5408, n5409, n5410, n5412, n5413, n5414, n5415, n5416, n5417, n5418;
  assign z034 = 1'b0;
  assign z000 = ~x2 & (~n524 | (~x3 & ~n523));
  assign n523 = (x1 | x6 | ((x0 | (x4 ? (~x5 | x7) : (x5 | ~x7))) & (~x0 | ~x4 | ~x5 | ~x7))) & (x0 | ~x1 | x4 | ~x5 | ~x6 | ~x7);
  assign n524 = x0 ? (x1 | ((~x3 | (x4 & (x5 | x6))) & (~x5 | ~x6 | x3 | ~x4))) : ((~x1 | (x3 ? (x4 | x5) : ~x4)) & (x3 | ((x1 | (x5 ? x4 : ~x6)) & (~x4 | x5))));
  assign z001 = n527 | n528 | (~x1 & (~n526 | (x5 & ~n529)));
  assign n526 = x0 ? (~x3 | ((x5 | ~x6 | x2 | ~x4) & (~x2 | x4 | ~x5 | x6))) : (x3 | ~x4 | (x2 ? (x5 | x6) : (~x5 | ~x6)));
  assign n527 = ~x1 & (x2 ? ((~x3 & ~x4) | (x0 & (~x3 | (~x4 & ~x5)))) : (x3 & (~x0 | (x4 & x5))));
  assign n528 = ~x0 & x1 & (x2 ? ~x3 : (x3 & (x4 | x5)));
  assign n529 = (~x0 | ~x2 | ~x3 | x4 | ~x6 | x7) & (x0 | x2 | x3 | ~x4 | x6 | ~x7);
  assign z002 = ~n531 | ~n533 | (~x0 & ~n532);
  assign n531 = x3 ? ((~x4 | (x0 ? (x1 | (~x2 & ~x5)) : (x5 | (~x1 & x2)))) & (x0 | ((x4 | (x1 & ~x2)) & (~x1 | x2 | ~x5)))) : ((~x0 | x4 | (x1 ? (x2 | x5) : ~x2)) & (x0 | x1 | ~x2 | ~x4 | ~x5));
  assign n532 = (~x2 | ((~x1 | x6 | (x3 ? (~x4 | ~x5) : (x4 | x5))) & (~x4 | x5 | ~x6 | x1 | x3))) & (~x4 | ~x5 | ~x6 | x1 | x2 | x3);
  assign n533 = (~n534 | ~n535) & (~x5 | (~n536 & ~n542));
  assign n534 = ~x2 & x0 & ~x1;
  assign n535 = x6 & ~x5 & x3 & x4;
  assign n536 = n541 & (x3 ? (n537 & n538) : (n539 & n540));
  assign n537 = x6 & x7;
  assign n538 = ~x1 & x2;
  assign n539 = x1 & ~x2;
  assign n540 = ~x6 & ~x7;
  assign n541 = x0 & ~x4;
  assign n542 = n545 & ((~x3 & n543 & ~x1 & ~x2) | (x1 & x2 & x3 & n544));
  assign n543 = ~x6 & x7;
  assign n544 = x6 & ~x7;
  assign n545 = ~x0 & x4;
  assign z003 = n547 | ~n553 | (x0 ? ~n551 : ~n552);
  assign n547 = ~x3 & ((~n548 & n549) | (n544 & n538 & ~n550));
  assign n548 = (x4 | ((x0 | (x1 ? (~x5 | ~x6) : (x5 | x6))) & (~x5 | x6 | ~x0 | ~x1))) & (~x5 | x6 | x1 | ~x4);
  assign n549 = ~x2 & x7;
  assign n550 = x0 ? (~x4 | ~x5) : (x4 | x5);
  assign n551 = (x1 | ((x2 | (x4 ^ x6) | (~x3 ^ x5)) & (~x5 | x6 | ~x2 | ~x4))) & (~x1 | x2 | x3 | x4 | ~x5 | ~x6);
  assign n552 = (x5 | (x1 ? ((x4 | ~x6 | ~x2 | x3) & (~x4 | x6 | x2 | ~x3)) : (x3 | (x2 ? (x4 ^ x6) : (x4 | ~x6))))) & (x1 | x2 | x3 | ~x5 | (x4 ^ x6));
  assign n553 = ~n554 & ~n555 & (~n558 | ~n559) & (n556 | n557);
  assign n554 = ~x2 & (x3 ? ((~x1 & x4 & x5) | (~x0 & ~x4 & (~x1 ^ x5))) : (~x5 & ((x1 & x4) | (x0 & ~x1 & ~x4))));
  assign n555 = x2 & ((~x0 & (x1 ? (~x4 & (x3 | x5)) : (x4 & x5))) | (~x1 & x4 & ~x5 & (x0 | x3)));
  assign n556 = (~x2 | ((~x3 | ~x5 | ~x6 | ~x7) & (x3 | x5 | x6 | x7))) & (x2 | ~x3 | x5 | ~x6 | x7);
  assign n557 = x0 ? (x1 | x4) : (~x1 | ~x4);
  assign n558 = x3 & x2 & ~x0 & ~x1;
  assign n559 = ~x7 & ~x6 & ~x4 & ~x5;
  assign z004 = ~n569 | (x1 ? ~n566 : (~n562 | (~x7 & ~n561)));
  assign n561 = (~x2 | ((~x5 | ((~x0 | (x3 ? (~x4 | ~x6) : (x4 | x6))) & (x4 | x6 | x0 | ~x3))) & (x0 | ~x3 | ~x4 | x5 | x6))) & (~x4 | x5 | ~x6 | ~x0 | x2 | ~x3);
  assign n562 = (~x0 | ((~n563 | ~n565) & (~x5 | ~x7 | n564))) & (x0 | x5 | x7 | n564);
  assign n563 = ~x2 & ~x3;
  assign n564 = (x2 | x6 | (x3 ^ ~x4)) & (~x2 | x3 | ~x4 | ~x6);
  assign n565 = x7 & x6 & ~x4 & x5;
  assign n566 = x0 ? (~n563 | ~n568) : n567;
  assign n567 = (~x7 | (((x3 ? (~x4 | ~x6) : (x4 | x6)) | (~x2 ^ ~x5)) & (x2 | x3 | ~x4 | ~x5 | x6))) & (x2 | x3 | ~x6 | x7 | (~x4 ^ ~x5));
  assign n568 = ~x7 & ~x6 & x4 & x5;
  assign n569 = n574 & (n571 | n572) & (x2 ? n573 : n570);
  assign n570 = x1 ? (x3 | (x5 ? (~x7 | (~x0 ^ x6)) : (x6 | x7))) : (x0 ? ((~x3 | (x5 ? (x6 | x7) : (~x6 | ~x7))) & (x3 | ~x5 | ~x6 | x7)) : ((x6 | ~x7 | x3 | x5) & (~x6 | x7 | ~x3 | ~x5)));
  assign n571 = x3 ? (x4 | ~x6) : (~x4 | x6);
  assign n572 = (x0 | ((~x1 | (x2 ? (x5 | ~x7) : (~x5 | x7))) & (x1 | x2 | ~x5 | ~x7))) & (~x2 | x5 | x7 | ~x0 | x1);
  assign n573 = (x1 | ~x7 | (x0 ? (x3 ? (~x5 | ~x6) : (x5 | x6)) : (x5 | (~x3 ^ x6)))) & (x0 | ~x1 | x7 | (x3 ? (x5 | ~x6) : (~x5 | x6)));
  assign n574 = x2 ? ((x5 | (((~x3 ^ x6) | (x0 ^ ~x1)) & (~x3 | ~x6 | x0 | x1))) & (x3 | ~x5 | x6 | x0 | x1)) : ((x3 | ((~x0 | (x1 ? (~x5 | ~x6) : (x5 | x6))) & (~x5 | ~x6 | x0 | x1))) & (~x5 | x6 | x0 | ~x3));
  assign z005 = ~n578 | (~x3 & (x6 ? (~x7 & ~n577) : ~n576));
  assign n576 = (x4 | ((x1 | ((~x0 | (x2 ? (~x5 | ~x7) : (x5 | x7))) & (~x5 | x7 | x0 | ~x2))) & (x0 | ~x1 | x2 | ~x5 | x7))) & (~x1 | x2 | ~x4 | x5 | ~x7);
  assign n577 = (x0 | ~x2 | ~x5 | (~x1 ^ x4)) & (x1 | x2 | ~x4 | x5);
  assign n578 = n581 & n584 & (x6 ? (x7 ? n579 : n580) : (x7 ? n580 : n579));
  assign n579 = (~x3 | x4 | ~x5 | ~x0 | x1 | ~x2) & (x0 | ((x2 | ((~x1 | x4 | (x3 ^ x5)) & (~x4 | ~x5 | x1 | ~x3))) & (x1 | ~x2 | x3 | x4 | x5)));
  assign n580 = (x3 | (x0 ? (x4 | (x1 ? x2 : (~x2 | x5))) : (~x4 | (x1 ? ~x2 : (x2 | ~x5))))) & (x1 | ~x3 | ((x0 | x4 | (~x2 & x5)) & (~x4 | ~x5 | ~x0 | x2)));
  assign n581 = x2 ? n583 : n582;
  assign n582 = x1 ? ((x3 | ~x4 | ~x5 | x6) & (~x3 | ((x4 | x5 | x6) & (~x5 | ~x6 | x0 | ~x4)))) : ((~x6 | ((x3 | x4) & (~x0 | ((x4 | ~x5) & (~x3 | ~x4 | x5))))) & (x0 | ~x3 | x6 | (~x4 ^ x5)));
  assign n583 = (x1 | ((~x4 | (x0 ? (~x3 ^ ~x6) : (x3 ? x6 : (x5 | ~x6)))) & (x0 | x3 | x4 | ~x5 | ~x6))) & (x0 | ~x1 | x4 | (x3 ? x6 : (x5 | ~x6)));
  assign n584 = (~x3 | n585) & (~n587 | (~n586 & ~n588));
  assign n585 = (x5 | ((~x0 | x1 | x4 | (x6 ^ x7)) & (~x4 | ~x6 | ~x7 | x0 | ~x1))) & (x0 | ~x1 | ~x4 | x6 | x7);
  assign n586 = ~x3 & x0 & ~x1;
  assign n587 = x7 & x6 & x4 & x5;
  assign n588 = x3 & x2 & ~x0 & x1;
  assign z006 = ~n590 | n600 | (~x2 & (n596 | (x4 & ~n595)));
  assign n590 = n594 & (x0 | n591) & (n592 | n593);
  assign n591 = (~x3 | ((~x1 | ((~x2 | (x4 ^ x7)) & (~x7 | ((~x4 | x5) & (x2 | x4 | ~x5))))) & (x1 | x2 | ~x4 | x5 | x7))) & (~x1 | ~x2 | x5 | (x4 ^ x7));
  assign n592 = x4 ^ ~x7;
  assign n593 = (x1 | ((~x2 | (~x3 & x5)) & (~x0 | ~x3 | x5))) & (~x1 | x2 | x3 | ~x5);
  assign n594 = (x2 | ((~x5 | ~x7 | x1 | ~x4) & (x4 | (x1 ? (x5 | (~x3 ^ x7)) : (~x5 | x7))))) & (x1 | ~x2 | x3 | ~x4 | ~x5 | x7);
  assign n595 = (x7 | (x1 ? (~x6 | ((x3 | x5) & (x0 | ~x3 | ~x5))) : (x6 | ((x3 | x5) & (~x0 | ~x3 | ~x5))))) & (x3 | x5 | ~x7 | (~x1 ^ x6));
  assign n596 = n597 & (x3 ? (n543 & n598) : (~x7 & ~n599));
  assign n597 = ~x4 & ~x5;
  assign n598 = ~x0 & ~x1;
  assign n599 = x1 ^ ~x6;
  assign n600 = n601 & ((((~x1 & x6) | (~x0 & x1 & ~x6)) & (~x4 ^ x7)) | (~x4 & x7 & (x0 ? (~x1 & ~x6) : (x1 & x6))));
  assign n601 = x5 & x2 & ~x3;
  assign z007 = n606 | ~n609 | (~x0 & (n604 | (x1 & ~n603)));
  assign n603 = (~x6 | ((~x2 | ((~x5 | ~x7 | x3 | ~x4) & (~x3 | x4 | x5 | x7))) & (~x4 | ~x5 | x7 | x2 | x3))) & (x2 | ~x5 | x6 | (x3 ? (~x4 | ~x7) : (x4 | x7)));
  assign n604 = x5 & n605 & ((x2 & x7 & (~x4 ^ x6)) | (x6 & ~x7 & ~x2 & x4));
  assign n605 = ~x1 & ~x3;
  assign n606 = ~n607 & ~n608;
  assign n607 = x2 ^ ~x7;
  assign n608 = (x4 | x5 | ((x1 | x3 | x6) & (x0 | ((x3 | x6) & (x1 | ~x3 | ~x6))))) & (~x0 | x1 | ~x3 | ~x4 | ~x5 | x6);
  assign n609 = (~x2 | n613) & (~n610 | n611) & (x2 | n612);
  assign n610 = x0 & ~x3;
  assign n611 = (~x4 | ~x6 | ((x1 | ~x2 | (x5 ^ x7)) & (x2 | ~x5 | x7))) & (~x1 | x2 | x4 | x5 | x6 | ~x7);
  assign n612 = (x3 & ((x0 & (x1 | (x4 & ~x6))) | ~x5 | (x1 & x4 & ~x6))) | (~x5 & ~x6) | (~x3 & ((x5 & x6) | (~x0 & x1 & ~x4 & ~x6)));
  assign n613 = (~x3 & (x6 ? ~x5 : ~x4)) | (x5 & (x3 | x4)) | (x0 & x1) | (~x5 & x6 & ~x0 & ~x4);
  assign z008 = ~n632 | n628 | n626 | n615 | ~n619;
  assign n615 = ~x1 & ((x6 & ~n617) | (~x4 & n616 & n618));
  assign n616 = ~x0 & x2;
  assign n617 = (x5 | ((~x0 | ~x4 | (x2 ? (x3 | ~x7) : (~x3 | x7))) & (x0 | ~x2 | ~x3 | x4 | ~x7))) & (~x4 | ~x5 | ~x7 | ~x0 | x2 | x3);
  assign n618 = x5 & ~x6 & (x3 ^ x7);
  assign n619 = ~n621 & ~n623 & (n620 | n625) & (x2 | n624);
  assign n620 = x6 ^ ~x7;
  assign n621 = ~n622 & (x1 ? ((~x2 & ~x3 & ~x6) | (~x0 & ((~x3 & ~x6) | (x2 & x3 & x6)))) : ((~x0 & ~x2 & x3 & x6) | (x0 & x2 & ~x3 & ~x6)));
  assign n622 = x4 ? (~x5 | x7) : (x5 | ~x7);
  assign n623 = ~x1 & ((x4 & ~x6 & ~x0 & x3) | (x0 & ~x4 & (x2 ? (~x3 & x6) : (x3 & ~x6))));
  assign n624 = (~x0 | ~x4 | x5 | (x1 ? (x3 | ~x6) : (~x3 | x6))) & (x4 | ~x5 | x6 | x0 | x1 | ~x3);
  assign n625 = (x0 | ((~x1 | x2 | ~x3 | ~x4 | ~x5) & (x4 | x5 | x1 | x3))) & (x1 | ((~x4 | ~x5 | ~x0 | ~x3) & (x4 | x5 | x2 | x3)));
  assign n626 = ~n627 & ((~x0 & ((~x3 & x6) | (x1 & ~x2 & x3 & ~x6))) | (~x1 & ((~x2 & ~x3 & x6) | (x0 & x2 & x3 & ~x6))));
  assign n627 = x4 ^ ~x5;
  assign n628 = n631 & ((n544 & n629) | (~x2 & ~n630));
  assign n629 = x2 & ~x5;
  assign n630 = x5 ? (x6 | ~x7) : (~x6 | x7);
  assign n631 = ~x4 & ~x3 & ~x0 & x1;
  assign n632 = ~n634 & ((x0 & (x1 ^ ~x2)) | (n633 & (~x1 | ~x2 | ~n635)));
  assign n633 = (x5 | x6 | x7 | ~x3 | x4) & (~x5 | ~x6 | ~x7 | x3 | ~x4);
  assign n634 = x1 & ((x0 & ~x2 & ~x3 & ~x4 & x6) | (~x0 & x2 & x3 & x4 & ~x6));
  assign n635 = ~x6 & x5 & x3 & ~x4;
  assign z009 = (~x4 & ~n646) | (x4 & ~n645) | (~x0 & ~n637) | (x0 & ~n640);
  assign n637 = (~x7 | n638) & (~x5 | x7 | n639);
  assign n638 = (~x5 | ((x1 | ((~x2 | (x4 ^ x6)) & (~x3 | ~x4 | ~x6))) & (~x1 | x2 | x3 | x4 | x6))) & (~x1 | x2 | x5 | (x3 ? (x4 | x6) : (~x4 | ~x6)));
  assign n639 = (x1 | (x4 ? (x6 | (x2 & x3)) : ~x6)) & (~x1 | ~x2 | ~x3 | ~x4 | x6);
  assign n640 = (x1 | n643) & (~n644 | (~n642 & (x3 | ~n641)));
  assign n641 = x4 & x6;
  assign n642 = ~x4 & ~x6;
  assign n643 = (x7 | ((x5 | ((~x2 | ((x4 | ~x6) & (x3 | ~x4 | x6))) & (~x3 | ((x4 | ~x6) & (x2 | ~x4 | x6))))) & (x2 | x3 | ~x5 | (~x4 ^ x6)))) & (x5 | ~x7 | ((~x3 | ~x4 | ~x6) & (~x2 | (x4 ^ x6))));
  assign n644 = x7 & ~x5 & x1 & ~x2;
  assign n645 = (x7 | ((x0 | (x5 & (x1 | ~x2 | ~x3))) & (x5 | ((x2 | x3) & (x1 | ~x2 | ~x3))))) & (~x5 | ~x7 | ((x0 | ~x1) & (~x0 | x1) & (x2 | x3)));
  assign n646 = (x3 | ((x2 | ((x1 | x5 | ~x7) & (~x5 | x7 | ~x0 | ~x1))) & (x0 | x5 | ~x7))) & (~x5 | x7 | (~x2 & ~x3) | (x0 ^ ~x1)) & (x0 | x5 | ~x7 | (x1 & ~x2));
  assign z010 = n649 | (n648 & ~n656) | (x3 & ~n654) | (~x3 & ~n655);
  assign n648 = ~x1 & x4;
  assign n649 = x1 & ((n650 & n651 & n653) | (~x0 & ~n652));
  assign n650 = x3 & ~x4;
  assign n651 = x0 & ~x2;
  assign n652 = (x6 | (x2 ? (~x3 | x7 | (~x4 ^ ~x5)) : (x3 | (~x4 ^ x5)))) & (x2 | ((x5 | ((x3 | (x4 ? x7 : (~x6 | ~x7))) & (~x6 | ~x7 | ~x3 | ~x4))) & (x3 | x4 | ~x5 | x7)));
  assign n653 = ~x5 & (~x6 | ~x7);
  assign n654 = x0 ? (x1 | (x5 ? (~x6 | (x2 & ~x7)) : (x6 | (~x2 & x7)))) : ((x5 | ((~x1 | (x7 ? x6 : x2)) & (x2 | x6 | ~x7) & (~x6 | (x1 & ~x2)))) & (x1 | ~x5 | x6 | (~x2 & x7)));
  assign n655 = x2 ? ((x1 | (x0 ? (~x5 ^ ~x6) : (~x5 | x6))) & (x0 | x5 | (~x1 & ~x6))) : (x5 ? (x1 ? (~x6 | ~x7) : (x6 | x7)) : ((~x0 | (x7 ? x6 : ~x1)) & (x1 | (~x6 & ~x7))));
  assign n656 = (~x3 | (~x0 ^ x5) | (x2 ? (~x6 | x7) : (x6 | ~x7))) & (~x0 | x2 | x3 | ~x5 | (~x6 & ~x7));
  assign z011 = n659 | n661 | ~n663 | n668 | (n658 & ~n673);
  assign n658 = ~x1 & ~x6;
  assign n659 = ~n620 & ~n660;
  assign n660 = x1 ? (x2 | (x3 & (x4 | (x0 & x5)))) : (~x2 | ~x3 | ((~x4 | ~x5) & (~x0 | (~x4 & ~x5))));
  assign n661 = ~n662 & ((~x0 & x3 & (x1 ? (x2 & x4) : (~x2 & ~x4))) | (~x1 & ~x2 & ~x3 & (x0 | x4)));
  assign n662 = ~x6 ^ ~x7;
  assign n663 = ~n666 & ~n667 & (~n664 | ~n665 | ~n565);
  assign n664 = ~x0 & x1;
  assign n665 = ~x2 & x3;
  assign n666 = ~x0 & x2 & ((~x1 & ~x6 & (~x3 | ~x4)) | (~x4 & x6 & x1 & x3));
  assign n667 = (x2 ? ~x3 : (x3 & x4)) & (x0 ? (~x1 & ~x6) : (x1 & x6));
  assign n668 = n670 & ((n669 & n672) | (~x0 & ~n671));
  assign n669 = x0 & x3;
  assign n670 = ~x1 & ~x2;
  assign n671 = (~x3 | ~x4 | x6 | x7) & (x3 | x4 | ~x6 | ~x7);
  assign n672 = ~x7 & ~x4 & ~x6;
  assign n673 = (~x3 | (~x0 ^ x4) | (x2 ? x5 : (~x5 | ~x7))) & (x4 | ~x5 | x7 | x0 | x2 | x3);
  assign z012 = n680 | n681 | ~n682 | (x3 & (~n675 | ~n679));
  assign n675 = (x4 | n676) & (~n677 | ~n678);
  assign n676 = (~x7 | (~x2 ^ x6) | (x0 ? (x1 | x5) : (~x1 | ~x5))) & (~x0 | x1 | x2 | x5 | x6 | x7);
  assign n677 = ~x2 & ~x0 & ~x1;
  assign n678 = x7 & x6 & x4 & ~x5;
  assign n679 = (x4 | ((~x1 | x5 | (x0 ? (x2 | x7) : (~x2 | ~x7))) & (~x0 | x1 | ~x5 | (~x2 ^ x7)))) & (x0 | x1 | ~x4 | (x2 ? (~x5 ^ x7) : (x5 ^ x7)));
  assign n680 = (~x2 | (x3 ^ x7)) & (x2 | (~x3 ^ x7)) & (~x0 | ~x1) & (~x3 | x4) & (x0 | x1);
  assign n681 = ~x0 & x3 & ~x4 & ((~x2 & ~x7) | (~x1 & x2 & x7));
  assign n682 = (~n685 | ~n686) & (~n683 | ~n677) & (x3 | n684);
  assign n683 = ~x7 & x5 & ~x3 & ~x4;
  assign n684 = (x0 | x1 | (x2 ? ~x7 : (~x4 | x7))) & (~x0 | ~x1 | x2 | x7);
  assign n685 = ~x3 & ~x2 & ~x0 & ~x1;
  assign n686 = ~x7 & x6 & ~x4 & ~x5;
  assign z013 = n689 | n695 | ~n696 | (~x1 & ~n688);
  assign n688 = (x4 | ((~x0 | x2 | (x5 ? x3 : ~x6)) & (x0 | ~x2 | x3 | x5 | x6))) & (x0 | ~x2 | x3 | ~x4 | x5 | ~x6);
  assign n689 = x6 & ((~n692 & ~n693) | (n690 & n691 & n694));
  assign n690 = ~x3 & ~x4;
  assign n691 = ~x5 & ~x7;
  assign n692 = ~x3 ^ ~x7;
  assign n693 = (~x2 | x4 | x5 | ~x0 | x1) & (x0 | ((x1 | x2 | ~x4 | x5) & (~x1 | x4 | ~x5)));
  assign n694 = ~x2 & x0 & x1;
  assign n695 = ~x3 & ((~x0 & ((x1 & ~x4 & x5 & ~x6) | (~x1 & ~x5 & (x4 ^ x6)))) | (x0 & ~x1 & ~x4 & ~x5 & ~x6));
  assign n696 = n697 & ((x0 & (x1 | ~x3)) | (~x0 & ((x3 & ~x4) | (~x1 & ~x5))) | (~x3 & x4) | (~x4 & (x5 ? x1 : x3)));
  assign n697 = (~n698 | ~n685) & (~n694 | ~n699);
  assign n698 = x7 & ~x6 & ~x4 & ~x5;
  assign n699 = ~x6 & ~x5 & ~x3 & ~x4;
  assign z014 = n705 | ~n706 | ~n711 | (~x2 & (~n701 | ~n704));
  assign n701 = (x3 | n702) & (x0 | ~x3 | ~x6 | n703);
  assign n702 = x1 ? (~x6 | (~x4 ^ x7) | (~x0 ^ x5)) : ((~x4 | ((~x6 | ~x7 | x0 | x5) & (x6 | x7 | ~x0 | ~x5))) & (x0 | x4 | x5 | (~x6 ^ x7)));
  assign n703 = x1 ? (~x5 | (~x4 ^ x7)) : (x5 | (x4 ^ x7));
  assign n704 = (x6 | ((~x4 | (x0 ? (x5 | (x1 ^ ~x3)) : (~x1 | ~x5))) & (~x3 | x4 | x5 | x0 | x1))) & (~x0 | x1 | ~x3 | x4 | x5 | ~x6);
  assign n705 = x0 & ~x1 & ~x2 & (x3 ? (~x4 & x5) : (x4 & ~x5));
  assign n706 = (x1 | ((x0 | ((~x2 | x4 | x5) & (~x4 | ~x5))) & (~x0 | ~x2 | x4 | ~x5))) & ~n707 & (~x4 | x5 | x0 | ~x1);
  assign n707 = ~x6 & n710 & ((x0 & n709) | (n664 & n708));
  assign n708 = ~x3 & x5;
  assign n709 = ~x1 & ~x5;
  assign n710 = x2 & x4;
  assign n711 = ~n712 & (~x2 | ~x6 | n713);
  assign n712 = x1 & ((x0 & ~x2 & ~x3 & ~x4 & x5) | (~x0 & ((~x4 & ~x5 & ~x2 & ~x3) | (x4 & x5 & x2 & x3))));
  assign n713 = x0 ? (x1 | x5 | (~x4 ^ x7)) : (~x1 | ~x5 | ((x4 | ~x7) & (x3 | ~x4 | x7)));
  assign z015 = n717 | ~n718 | n722 | n725 | (~x2 & ~n715);
  assign n715 = (~x4 | n716) & (~x5 | ~n631 | (x6 & ~n544));
  assign n716 = x0 ? (x1 | ~x5 | (x3 ? (~x6 | x7) : (x6 | ~x7))) : (~x1 | x3 | x5 | (x6 & x7));
  assign n717 = ~x2 & ~x6 & ((x3 & ~x5 & ~x0 & x1) | (x0 & ~x1 & (x3 ^ ~x5)));
  assign n718 = (x0 | ~x2 | (x1 ? (x5 | x6) : ~x5)) & ~n719 & (~x0 | x1 | x2 | x5 | ~x6);
  assign n719 = (x5 | (x6 & x7)) & (n720 | (~x1 & ~n721)) & (~x5 | ~x6 | ~x7);
  assign n720 = ~x3 & ~x2 & x0 & x1;
  assign n721 = ~x0 ^ ~x2;
  assign n722 = n724 & ((n723 & (~x2 | ~x3)) | (n691 & (x2 | x3)));
  assign n723 = x5 & x7;
  assign n724 = x6 & ~x0 & x1;
  assign n725 = n588 & ~n627 & x6 & x7;
  assign z016 = (~x6 & (~n728 | (~x7 & ~n727))) | ~n729 | (x6 & x7 & ~n727);
  assign n727 = (~x0 & ((~x1 & x2) | (~x4 & ~x5 & ~x2 & ~x3))) | (x1 & x2 & x3 & x4) | (x0 & (x1 ? (x2 | x3) : (~x2 & (~x4 | ~x5))));
  assign n728 = (x1 | (x0 ? (x2 | x3 | (x4 & x5)) : (~x2 | (~x3 & ~x4 & ~x5)))) & (x0 | ((~x4 | ~x5 | ~x2 | ~x3) & (~x1 | x2 | x3 | x4 | x5)));
  assign n729 = ~n737 & ~n731 & (x7 | ~n730 | ~n616 | n739);
  assign n730 = ~x5 & ~x6;
  assign n731 = ~x2 & ((~n734 & n735) | (n732 & n733 & ~n736));
  assign n732 = ~x0 & ~x3;
  assign n733 = ~x4 & x7;
  assign n734 = (x4 | x5 | x6 | ~x1 | ~x3) & (x1 | x3 | ~x4 | ~x5 | ~x6);
  assign n735 = x0 & ~x7;
  assign n736 = x1 ? (~x5 | x6) : (x5 | ~x6);
  assign n737 = x6 & n665 & n738 & (~x4 | ~x5);
  assign n738 = x0 & ~x1;
  assign n739 = x1 ? (~x3 | ~x4) : (x3 | x4);
  assign z017 = ~n749 | n748 | n747 | n741 | n744;
  assign n741 = ~x0 & ((n742 & n686) | (x7 & ~n743));
  assign n742 = ~x3 & ~x1 & x2;
  assign n743 = (~x1 | ((x2 | x3 | x4 | ~x5 | ~x6) & (~x2 | ~x3 | ~x4 | x5 | x6))) & (x1 | ~x2 | x3 | x4 | x5 | x6);
  assign n744 = ~x1 & ((~x3 & n745 & ~x0 & x2) | (x3 & n746 & x0 & ~x2));
  assign n745 = ~x7 & ~x4 & x5;
  assign n746 = x4 & (x5 ^ ~x7);
  assign n747 = ~x7 & ((~x0 & ~x3 & (x1 ? (~x2 & ~x4) : (x2 & x4))) | (x0 & ~x1 & ~x2 & x3 & ~x4));
  assign n748 = ~x1 & (x0 ? (x2 ? x7 : (~x3 & ~x7)) : (x2 ? (x3 & ~x7) : x7));
  assign n749 = ~n751 & ~n752 & (~n750 | ~n753) & (~n698 | ~n754);
  assign n750 = x2 & ~x0 & x1;
  assign n751 = x1 & x7 & (x0 ? (~x2 & ~x3) : (x2 ^ x3));
  assign n752 = ~x0 & x1 & x7 & (x2 ? (x3 & ~x4) : (~x3 & x4));
  assign n753 = ~x7 & x5 & x3 & x4;
  assign n754 = x3 & ~x2 & x0 & x1;
  assign z018 = n756 | ~n760 | (~x2 & (~n765 | n766 | n771));
  assign n756 = n616 & ((n757 & n758) | (~x1 & ~n759));
  assign n757 = ~x6 & x4 & ~x5;
  assign n758 = x1 & x3;
  assign n759 = (x3 | x4 | x5 | x6) & (~x3 | ~x4 | ~x5 | ~x6);
  assign n760 = ~n761 & n763 & n764 & (~n588 | ~n762);
  assign n761 = ~x1 & ((x0 & x3 & (~x2 ^ x4)) | (~x3 & x4 & ~x0 & ~x2));
  assign n762 = ~x7 & x6 & x4 & ~x5;
  assign n763 = ~x1 | ((~x0 | x2 | x3) & (~x3 | x4 | x0 | ~x2));
  assign n764 = (x0 | (x1 ? (x3 | (~x2 & (x4 | x5))) : (x2 | ~x3))) & (x1 | x2 | ~x3 | ~x4 | x5);
  assign n765 = x0 ? ((x1 | x3 | ~x4 | ~x5 | ~x6) & (~x1 | ~x3 | x4 | x5 | x6)) : (x3 | x4 | ~x5 | (x1 ^ ~x6));
  assign n766 = x0 & ((n767 & n770) | (n768 & n769));
  assign n767 = ~x7 & ~x5 & x6;
  assign n768 = x7 & x5 & ~x6;
  assign n769 = x4 & ~x1 & ~x3;
  assign n770 = ~x4 & x1 & x3;
  assign n771 = n664 & n772;
  assign n772 = x5 & x6 & (x3 ? (x4 & x7) : (~x4 & ~x7));
  assign z019 = x0 ? (~n777 | (~x2 & ~n778)) : (~n774 | ~n776);
  assign n774 = x1 ? n775 : (~n563 | ~n698);
  assign n775 = (~x4 | ((~x2 | ((x6 | ~x7 | x3 | ~x5) & (~x3 | x5 | ~x6 | x7))) & (x2 | ~x3 | ~x5 | ~x6 | x7))) & (x2 | ~x3 | x4 | x5 | x6 | ~x7);
  assign n776 = (~x6 | ((~x1 | ((~x3 | x4) & (~x2 | x3 | ~x4 | ~x5))) & (x1 | x2 | x3 | x4 | x5))) & (x4 | ((~x2 | ~x3) & (x1 | x6 | (~x2 ^ x5)))) & (~x3 | (((x2 & x6) | (x5 ? x1 : ~x4)) & (x1 | ~x4 | x5) & (x2 | ~x5 | x6)));
  assign n777 = (x2 | ((~x1 | x3 | (~x4 & (~x5 | ~x6))) & (~x3 | x5 | (x1 & (x4 | x6))))) & (x1 | (x3 ? x4 : (~x4 | (~x6 & (~x2 | ~x5)))));
  assign n778 = (x1 | x3 | ~x4 | x6 | (~x5 ^ x7)) & (x5 | ~x6 | x7 | ~x1 | ~x3 | x4);
  assign z020 = ~n780 | n791 | (~x0 & (~x4 | ~n789) & (x4 | ~n790));
  assign n780 = n782 & ~n787 & (x6 ? (x3 | n788) : n781);
  assign n781 = (~x0 | ((~x1 | x2 | x4 | (~x3 ^ x5)) & (x3 | ~x4 | x5 | x1 | ~x2))) & (~x3 | ~x4 | ~x5 | x0 | x1 | ~x2);
  assign n782 = ~n784 & (n785 | (x3 ? n786 : (~n598 | n783)));
  assign n783 = ~x4 ^ ~x6;
  assign n784 = ~x1 & ((x5 & (x0 ? (~x4 & (x2 | ~x3)) : (x4 & (x2 ^ x3)))) | (x3 & ~x5 & (x0 ? (~x2 & x4) : (~x2 ^ x4))));
  assign n785 = x2 ^ ~x5;
  assign n786 = (~x4 | x6 | x0 | ~x1) & (x4 | ~x6 | ~x0 | x1);
  assign n787 = x1 & ((~x0 & (x2 ? (x3 ? (~x4 & x5) : (x4 & ~x5)) : (x4 & (x3 ^ x5)))) | (~x3 & ~x4 & ~x5 & x0 & ~x2));
  assign n788 = (x1 | x2 | x4 | x5) & (~x1 | ((x0 | (x2 ? (x4 | ~x5) : (~x4 | x5))) & (~x4 | ~x5 | ~x0 | x2)));
  assign n789 = ((x3 ? (x5 | ~x6) : (~x5 | x6)) | (x1 ? (~x2 | x7) : (x2 | ~x7))) & (~x1 | x2 | ~x3 | ~x5 | ~x6 | x7) & (x1 | ~x2 | x3 | x5 | x6 | ~x7);
  assign n790 = (~x7 | ((~x1 | x2 | x3 | ~x5 | x6) & (x1 | ((~x2 | ~x3 | ~x5 | ~x6) & (x2 | x3 | x5 | x6))))) & (~x1 | x2 | x7 | (x3 ? (x5 | x6) : (~x5 | ~x6)));
  assign n791 = x0 & ((x7 & n538 & ~n793) | (~x2 & ~n792));
  assign n792 = (x5 | ~x6 | x7 | ~x1 | ~x3 | x4) & (x6 | ((~x5 | ~x7 | x3 | ~x4) & (x1 | ((~x5 | ~x7 | ~x3 | x4) & (x3 | ~x4 | x5 | x7)))));
  assign n793 = (x5 | ~x6 | x3 | x4) & (~x3 | (x4 ? (~x5 | ~x6) : (x5 | x6)));
  assign z021 = n795 | ~n799 | n805 | n807 | (~x2 & ~n798);
  assign n795 = ~x1 & ((~x2 & ~n796) | (x0 & x2 & ~n797));
  assign n796 = x0 ? (~x3 | ((~x4 | ~x7 | (~x5 ^ ~x6)) & (x4 | ~x5 | x6 | x7))) : (x3 | ((~x6 | ~x7 | x4 | x5) & (x6 | x7 | ~x4 | ~x5)));
  assign n797 = (x5 | x6 | x7 | ~x3 | x4) & (x3 | ((x4 | x5 | ~x6 | x7) & (x6 | ~x7 | ~x4 | ~x5)));
  assign n798 = x4 ? ((x0 | (((x3 ^ x5) | (x1 ^ ~x6)) & (~x1 | x3 | ~x5 | ~x6))) & (~x0 | x1 | x3 | ~x5 | x6)) : (((x0 ? (x3 | x6) : (~x3 | ~x6)) | (x1 ^ x5)) & (~x0 | ((x1 | x3 | ~x5 | ~x6) & (x5 | x6 | ~x1 | ~x3))) & (x0 | x3 | (x1 ? (x5 | ~x6) : (~x5 | x6))));
  assign n799 = ~n802 & ~n803 & (n800 | n804) & (~x2 | n801);
  assign n800 = x5 ^ ~x7;
  assign n801 = (x0 | (((x1 ? (~x3 | ~x6) : (x3 | x6)) | (~x4 ^ ~x5)) & (~x1 | x3 | x4 | ~x5 | x6) & (~x4 | x5 | ~x6 | x1 | ~x3))) & (x4 | ~x5 | ~x6 | ~x0 | x1 | ~x3);
  assign n802 = x2 & ((x0 & ~x1 & ~x3 & ~x5 & ~x6) | ((x3 ^ x6) & ((~x1 & x5) | (~x0 & x1 & ~x5))));
  assign n803 = ~x2 & ~x5 & ((x0 & x6 & (x1 ^ x3)) | (x3 & ~x6 & ~x0 & ~x1));
  assign n804 = (((~x3 | ~x6 | x1 | ~x2) & (~x1 | x2 | x3 | x6)) | (x0 ^ x4)) & (x0 | ~x1 | ~x4 | (x2 ? (x3 | x6) : (~x3 | ~x6)));
  assign n805 = ~n806 & ((~x2 & ~x3 & ~x6 & x0 & ~x1) | (~x0 & ((x1 & x2 & x3 & x6) | (~x1 & (x2 ? (~x3 & ~x6) : (x3 & x6))))));
  assign n806 = x4 ? (x5 | x7) : (~x5 | ~x7);
  assign n807 = n808 & ((~x0 & ((x3 & ~x6 & (~x5 ^ x7)) | (~x3 & x5 & x6 & x7))) | (x0 & x3 & ~x5 & x6 & ~x7));
  assign n808 = ~x4 & x1 & ~x2;
  assign z022 = n810 | n813 | ~n818 | (~n662 & ~n817);
  assign n810 = x0 & ((~x1 & ~n812) | (n686 & n811));
  assign n811 = x3 & x1 & ~x2;
  assign n812 = (~x2 | (x3 ? (~x4 | (~x6 ^ x7)) : (x4 | ((x6 | ~x7) & (x5 | ~x6 | x7))))) & (~x4 | ~x5 | ((~x3 | ~x6 | x7) & (x6 | ~x7 | x2 | x3)));
  assign n813 = ~x0 & ((n814 & ~n816) | (~x4 & ~n815));
  assign n814 = x3 & x4;
  assign n815 = (x6 | ((x3 | (x1 ? ((~x5 | x7) & (~x2 | x5 | ~x7)) : (x5 | (x2 ^ ~x7)))) & (~x5 | ~x7 | ~x2 | ~x3))) & (~x3 | ~x6 | ((~x5 | x7) & (x1 | (x2 ? x7 : (x5 | ~x7)))));
  assign n816 = x6 ? (x7 | ((x2 | x5) & (~x1 | (x2 & x5)))) : (~x7 | ((~x1 | ~x2 | x5) & (~x5 | (x1 & x2))));
  assign n817 = (x0 | ((~x5 | ((x1 | ~x2 | (~x3 ^ ~x4)) & (x3 | ~x4 | (~x1 & x2)))) & (~x1 | x2 | x4 | (~x3 & x5)) & (~x4 | x5 | ~x2 | x3))) & (~x0 | ((x3 | ((x2 | (~x4 ^ x5)) & (~x4 | ~x5 | x1 | ~x2))) & (x1 | ((~x3 | x4 | x5) & (x2 | (x4 & x5)))))) & (x2 | x3 | ~x4 | (x1 ^ x5));
  assign n818 = ~n822 & (~x2 | n819) & (n820 | n821);
  assign n819 = (x1 | (x0 ? ((x3 | ~x4 | x5 | x6) & (~x5 | ~x6 | ~x3 | x4)) : (~x4 | (x3 ? (x5 | x6) : (~x5 | ~x6))))) & (x0 | ~x1 | ~x3 | (x4 ? (~x5 | x6) : (x5 | ~x6)));
  assign n820 = (x2 | (x0 ? (x4 ? (~x6 | x7) : (x6 | ~x7)) : (x4 ? (x6 | ~x7) : (~x6 | x7)))) & (x0 | ~x2 | x4 | x6 | ~x7);
  assign n821 = x1 ? (x3 | ~x5) : x5;
  assign n822 = ~x6 & n563 & ((x0 & x1 & ~x4 & ~x5) | (~x0 & (x1 ? (x4 & ~x5) : (~x4 & x5))));
  assign z023 = n825 | ~n832 | (~n800 & ~n830) | (~n824 & ~n831);
  assign n824 = ~x5 ^ ~x7;
  assign n825 = ~x2 & (~n827 | (~x0 & ~n826));
  assign n826 = (~x6 | ((x7 | ((x1 | x3 | ~x4 | ~x5) & (~x1 | (x3 ? (~x4 | ~x5) : (x4 | x5))))) & (x4 | x5 | ~x7 | x1 | ~x3))) & (x3 | x6 | ~x7 | (x1 ? ~x4 : (x4 | ~x5)));
  assign n827 = ~n829 & (~n738 | ~n828) & (~n586 | ~n587);
  assign n828 = x7 & x4 & ~x5;
  assign n829 = ~x4 & ((x0 & ((~x1 & x6 & ~x7) | (~x6 & x7 & x1 & ~x5))) | (~x0 & x1 & x5 & ~x6 & ~x7));
  assign n830 = x1 ? ((~x0 | x2 | x3 | x4 | ~x6) & (x0 | ((x2 | ~x4 | (~x3 ^ x6)) & (x4 | ~x6 | ~x2 | ~x3)))) : (x0 ? (x2 ? (x3 | ~x4) : (x4 | x6)) : ((~x2 | (x3 ? (~x4 | ~x6) : x4)) & (~x4 | x6 | x2 | x3)));
  assign n831 = (x6 | ((~x0 | x1 | x2 | ~x4) & (x3 | x4 | x0 | ~x1))) & (x1 | ((~x2 | (x0 ? (x4 | (~x3 & ~x6)) : (x3 | ~x4))) & (x0 | x2 | ~x6 | (~x3 ^ ~x4)))) & (x0 | ((~x4 | ~x6 | ~x2 | x3) & (~x1 | ~x3 | (x2 ^ x4)))) & (~x0 | ~x1 | x2 | x3 | ~x4);
  assign n832 = (n592 | n833) & (~x2 | (~n835 & (x1 | n834)));
  assign n833 = x0 ? ((~x1 | x2 | x3 | ~x5 | x6) & (~x3 | x5 | ~x6 | x1 | ~x2)) : ((x1 | x2 | (x3 ? x6 : (x5 | ~x6))) & (~x1 | ~x2 | x3 | ~x5 | ~x6));
  assign n834 = (x7 | (x0 ? (x3 ? (~x4 | ~x5) : (x4 | x6)) : (~x3 | x4 | (~x5 & ~x6)))) & (x0 | ~x4 | ~x7 | (x3 ? x6 : (x5 | ~x6)));
  assign n835 = n664 & (x3 ? (~x4 & n836) : (n837 | n838));
  assign n836 = x7 & ~x5 & ~x6;
  assign n837 = x7 & x6 & ~x4 & ~x5;
  assign n838 = ~x7 & x4 & ~x6;
  assign z024 = ~n845 | (x3 ? ~n840 : (x2 ? ~n844 : ~n843));
  assign n840 = x1 ? n842 : n841;
  assign n841 = (x7 | ((x4 | ((x0 | (x2 ? (x5 | x6) : (~x5 | ~x6))) & (x5 | ~x6 | ~x0 | ~x2))) & (~x0 | ~x4 | ((x5 | x6) & (x2 | ~x5 | ~x6))))) & (~x2 | ~x4 | ~x7 | (x0 ? (~x5 | x6) : (x5 | ~x6)));
  assign n842 = (x0 | (x4 ? ((~x2 | ~x7 | (~x5 ^ ~x6)) & (~x6 | x7 | x2 | x5)) : (x6 | ((~x5 | x7) & (x2 | x5 | ~x7))))) & (x5 | ~x6 | x7 | ~x0 | x2 | x4);
  assign n843 = x0 ? ((~x4 | ((~x5 | x6 | x7) & (x1 | ((~x5 | ~x6 | ~x7) & (x6 | x7))))) & (~x1 | x4 | x5 | ~x6 | ~x7)) : ((~x1 | ((x4 | ~x5 | x6 | x7) & (~x6 | ~x7 | ~x4 | x5))) & (x4 | ~x7 | (~x5 ^ ~x6)) & (x1 | ((~x6 | x7 | x4 | x5) & (x6 | ~x7 | ~x4 | ~x5))));
  assign n844 = (~x7 | ((x1 | ((x0 | x4 | ~x5 | ~x6) & (x5 | (x0 ? (~x4 ^ x6) : (x4 | x6))))) & (x0 | ~x1 | (x4 ? (x5 | ~x6) : (~x5 | x6))))) & (x0 | ~x4 | ~x6 | x7 | (x1 ^ x5));
  assign n845 = n849 & (n846 | n848) & (~x3 | n847);
  assign n846 = ~x5 ^ ~x6;
  assign n847 = (~x0 | ((~x1 | x2 | x4 | x5 | x6) & (~x4 | ~x5 | ~x6 | x1 | ~x2))) & (x1 | x2 | ~x4 | ~x5 | x6) & (x0 | (x1 ? (x5 | ~x6 | (~x2 & x4)) : (~x5 | (x4 ? x6 : ~x2))));
  assign n848 = (x1 | (x0 ? (x4 | (x2 & ~x3)) : (x3 | ~x4))) & (x0 | ~x1 | (x2 ? (x3 | x4) : (~x3 | ~x4)));
  assign n849 = (x3 | (x0 ? (n850 | (x1 ^ ~x2)) : n851)) & (x0 | x1 | x2 | ~x3 | n850);
  assign n850 = x4 ? (x5 | ~x6) : (~x5 | x6);
  assign n851 = (x1 | ~x2 | x4 | x5 | ~x6) & (~x1 | ((~x4 | ~x5 | x6) & (x2 | x4 | x5 | ~x6)));
  assign z025 = ~n859 | (x2 ? ~n855 : (x5 ? ~n854 : ~n853));
  assign n853 = x1 ? ((x3 | ~x4 | x6 | ~x7) & (~x0 | ~x3 | x4 | ~x6 | x7)) : (x0 ? ((~x6 | x7 | ~x3 | ~x4) & (x4 | x6 | ~x7)) : ((~x6 | ~x7 | ~x3 | x4) & (~x4 | x6 | (x3 & ~x7))));
  assign n854 = (x1 | ((~x0 | (x4 ? (~x6 | x7) : (x6 | ~x7))) & (~x4 | x6 | ~x7 | x0 | ~x3))) & (x0 | x7 | ((x4 | ~x6) & (~x1 | x3 | ~x4 | x6)));
  assign n855 = (x0 | n858) & (n856 | n857) & (~x0 | ~n605 | ~n587);
  assign n856 = (x6 | ~x7 | x4 | x5) & (~x6 | x7 | ~x4 | ~x5);
  assign n857 = x0 ^ ~x1;
  assign n858 = (x4 | ((x1 | ~x6 | (x3 ? ~x5 : x7)) & (~x1 | ~x3 | x5 | x6 | x7))) & (x1 | ~x4 | x5 | x6 | ~x7);
  assign n859 = (n630 | n860) & (n662 | n861);
  assign n860 = (~x1 | ((x0 | ~x4) & (x3 | x4 | ~x0 | x2))) & (x1 | (x0 ? (x2 ? x4 : (x3 | ~x4)) : (x2 | x4))) & (x0 | ~x2 | ~x4);
  assign n861 = x4 ? (x1 ? ((~x0 | x2 | x3) & (~x3 | x5 | x0 | ~x2)) : (x0 ^ (~x5 | (x2 & x3)))) : ((x1 | (x0 ? (~x5 | (x2 & x3)) : (~x2 | x5))) & (x0 | ((~x2 | x3 | x5) & (~x1 | (x2 & ~x5)))));
  assign z026 = ~n874 | ((~x0 | ~n863) & (n867 | n870 | x0 | n866));
  assign n863 = (n824 | n865) & (~x1 | ~n665 | ~n698) & (x1 | n864);
  assign n864 = (~x5 | x6 | ~x7 | x2 | x4) & (x5 | ((x2 | ~x4 | (x3 ? (~x6 | ~x7) : (x6 | x7))) & (~x2 | ~x3 | x4 | x6 | x7)));
  assign n865 = (x2 | ((~x4 | x6 | x1 | ~x3) & (x4 | ~x6 | ~x1 | x3))) & (x1 | ~x2 | (x6 ? (~x3 & ~x4) : x3));
  assign n866 = ~n824 & (x1 ? (~x2 & (x6 | (~x3 & x4))) : (x2 & (x6 ? x3 : (~x3 | ~x4))));
  assign n867 = ~n868 & ((~x1 & ~x2 & x3 & n543) | (x1 & x2 & n869));
  assign n868 = ~x4 ^ ~x5;
  assign n869 = ~x7 & ~x3 & x6;
  assign n870 = n873 & ((n563 & n872) | (n871 & n757));
  assign n871 = x2 & x3;
  assign n872 = x6 & ~x4 & x5;
  assign n873 = ~x1 & ~x7;
  assign n874 = (x0 | n877) & (n800 | n875) & (~x0 | n876);
  assign n875 = (x2 | ((~x0 | (x1 ? (x3 | x6) : (x4 | ~x6))) & (~x3 | ((x1 | x4 | ~x6) & (~x4 | x6 | x0 | ~x1))) & (x1 | ((x3 | ~x4 | ~x6) & (x0 | (x6 ? ~x4 : x3)))))) & (x0 | ~x2 | ((x3 | (x1 ? x6 : (x4 | ~x6))) & (~x1 | (x6 ? ~x3 : x4))));
  assign n876 = (~x4 | ~x5 | ~x6 | ~x1 | x2 | x3) & (x1 | ((x5 | x6 | x2 | x4) & (~x2 | ((x5 | ~x6 | x3 | x4) & (~x3 | ~x5 | x6)))));
  assign n877 = (x6 | (x1 ? ((x2 | x4 | ~x5) & (~x4 | x5 | ~x2 | ~x3)) : (~x3 | ~x4 | (x2 ^ x5)))) & (~x2 | x3 | ~x6 | (x1 ? (x4 | ~x5) : (~x4 | x5)));
  assign z027 = n879 | n882 | n884 | ~n888 | (~x0 & ~n881);
  assign n879 = ~n620 & ~n880;
  assign n880 = (~x5 | ((~x0 | x1 | x2 | ~x3 | ~x4) & (~x2 | x3 | x4 | x0 | ~x1))) & ((x0 ? (~x1 | x2) : (x1 | ~x2)) | (x3 ? (x4 | x5) : ~x4)) & (x3 | ((x0 | ((x1 | x2 | x4) & (~x2 | ~x4 | x5))) & (~x0 | x1 | ~x2 | x4)));
  assign n881 = (~x4 | ((~x6 | ((x1 | ~x2 | ~x3 | x5) & (~x1 | x3 | (x2 ^ x5)))) & (x1 | x2 | ~x3 | ~x5 | x6))) & (~x2 | x4 | ((~x5 | ~x6 | x1 | ~x3) & (x5 | x6 | ~x1 | x3)));
  assign n882 = ~n662 & ~n883;
  assign n883 = x0 ? (x1 | ((~x4 | ~x5 | x2 | x3) & (~x3 | (x2 ? (~x4 ^ x5) : (x4 | x5))))) : ((~x1 | (x2 ? (~x3 | ~x4) : x4)) & (~x3 | (x2 ? (~x4 | ~x5) : ((x4 | ~x5) & (x1 | ~x4 | x5)))));
  assign n884 = ~x2 & ((~x3 & ~n885 & ~n886) | (~x1 & x3 & ~n887));
  assign n885 = ~x1 ^ ~x4;
  assign n886 = (~x0 | x5 | x6 | x7) & (x0 | ~x5 | ~x6 | ~x7);
  assign n887 = (~x5 | x6 | x7 | ~x0 | ~x4) & (x0 | x4 | x5 | ~x6 | ~x7);
  assign n888 = ~n890 & ~n891 & (x3 ? (~n538 | n887) : n889);
  assign n889 = x0 ? ((x1 | ~x2 | ~x4 | ~x6) & (~x1 | x2 | x4 | x6)) : (x1 | (x2 ? (x4 | x6) : (~x4 | ~x6)));
  assign n890 = ~x0 & x1 & x3 & (x2 ? (~x4 & x6) : (x4 & ~x6));
  assign n891 = n738 & (n892 | (~x2 & ~x6 & ~n627));
  assign n892 = x6 & ~x5 & ~x4 & x2 & x3;
  assign z028 = n896 | n902 | n903 | (x1 ? ~n894 : ~n895);
  assign n894 = (x0 | (x4 ? (x2 ? (x3 | (x5 ^ x7)) : (~x7 | (~x3 & x5))) : (x7 | (x2 & (x3 | ~x5))))) & (x2 | x4 | x5 | ((~x3 | x7) & (~x0 | x3 | ~x7)));
  assign n895 = x4 ? ((~x7 | ((~x0 | (x2 ? x3 : x5)) & (x2 | x3 | x5) & (x0 | (x2 ? (~x3 | x5) : ~x5)))) & (x0 | x7 | (x2 ? (x3 | ~x5) : (~x3 | x5)))) : ((~x0 | ((x2 | (x5 ^ x7)) & (x7 | (x5 ? ~x2 : x3)))) & (~x5 | x7 | x0 | x2));
  assign n896 = ~x3 & (~n899 | (x6 & n897 & ~n898));
  assign n897 = ~x0 & ~x2;
  assign n898 = (~x5 | x7 | ~x1 | ~x4) & (x1 | x4 | (~x5 ^ ~x7));
  assign n899 = x4 ? (x7 | ((~x5 | n900) & (~x0 | x5 | n901))) : (~x7 | ((x5 | n900) & (x0 | ~x5 | n901)));
  assign n900 = (~x2 | x6 | x0 | ~x1) & (x2 | ~x6 | ~x0 | x1);
  assign n901 = x1 ? (x2 | ~x6) : (~x2 | x6);
  assign n902 = ~n592 & (x0 ? ((x3 & ~x5 & ~x1 & x2) | (x1 & ~x2 & ~x3 & x5)) : (x2 & ((~x1 & ~x3 & ~x5) | (x3 & (x1 | x5)))));
  assign n903 = ~n550 & n904 & (x2 ? (x6 ^ ~x7) : (~x6 ^ ~x7));
  assign n904 = ~x1 & x3;
  assign z029 = n907 | n908 | ~n909 | n915 | (~n906 & ~n914);
  assign n906 = x3 ^ ~x7;
  assign n907 = ~x0 & (x1 ? ((x3 & x4 & ~x5) | (~x4 & x5 & x2 & ~x3)) : (x4 & (~x3 ^ x5)));
  assign n908 = x0 & ~x4 & ((~x2 & (x1 ? (~x3 & ~x5) : x5)) | (~x1 & ((x3 & x5) | (x2 & ~x3 & ~x5))));
  assign n909 = n913 & ~n911 & (~n597 | n910 | x6 | ~n732);
  assign n910 = x1 ^ ~x2;
  assign n911 = ~n912 & ((x3 & ~x4 & ~x0 & ~x1) | (x4 & ~n910 & x0 & ~x3));
  assign n912 = x5 ^ ~x6;
  assign n913 = (x0 | ~x1 | ((~x5 | ~x6 | x3 | ~x4) & (x5 | x6 | ~x3 | x4))) & (~x4 | ~x5 | ~x6 | ~x0 | x1 | ~x3);
  assign n914 = (x0 | ((~x1 | ((~x4 | ~x5 | x6) & (x5 | ~x6 | ~x2 | x4))) & (~x5 | ~x6 | x1 | x4))) & (~x4 | x5 | x6 | ~x0 | x1 | ~x2);
  assign n915 = ~x2 & ((~n917 & ~n918) | (x7 & n916 & ~n919));
  assign n916 = ~x3 & ~x5;
  assign n917 = (~x4 | x6 | ~x0 | x1) & (x4 | ~x6 | x0 | ~x1);
  assign n918 = x3 ? (x5 | x7) : (~x5 | ~x7);
  assign n919 = (x0 | x1 | x4 | x6) & (~x0 | (x1 ? (~x4 | x6) : (x4 | ~x6)));
  assign z030 = n922 | n926 | n930 | n932 | (n677 & n921);
  assign n921 = x6 & ~x5 & ~x3 & ~x4;
  assign n922 = x6 & ((~n592 & ~n925) | (n923 & n691 & n924));
  assign n923 = ~x3 & x4;
  assign n924 = ~x2 & ~x0 & x1;
  assign n925 = (x2 | x3 | x5 | ~x0 | x1) & (x0 | (x1 ? (x5 | (~x2 & ~x3)) : ~x5));
  assign n926 = ~x6 & ((~n927 & ~n928) | (~x2 & ~n929));
  assign n927 = ~x4 ^ ~x7;
  assign n928 = (x2 | x3 | x5 | ~x0 | ~x1) & ((~x2 & ~x3) | (x0 ? (x1 | x5) : (~x1 | ~x5)));
  assign n929 = (x0 | ~x1 | x3 | ~x4 | ~x5 | ~x7) & (~x0 | x4 | x7 | (x1 ? (~x3 | x5) : (x3 | ~x5)));
  assign n930 = x4 & ~n931;
  assign n931 = (x1 | ((x0 | ~x5 | x6) & (x2 | x3 | ((x5 | x6) & (~x0 | ~x5 | ~x6))))) & (x0 | ~x1 | (x5 ? ~x6 : (x6 | (~x2 & ~x3))));
  assign n932 = ~n933 & (x0 ? (x4 ? x6 : (x5 & ~x6)) : (~x5 & (x4 ^ x6)));
  assign n933 = x1 ^ (~x2 & ~x3);
  assign z031 = n938 | (x2 ? ~n939 : (~n935 | ~n940));
  assign n935 = (x3 | n936) & (~n698 | ~n937);
  assign n936 = (~x5 | (x4 ^ x6) | (x0 ? (x1 | ~x7) : (~x1 | x7))) & (x0 | ~x1 | x5 | (x4 ? (x6 ^ x7) : (~x6 | x7)));
  assign n937 = x3 & x0 & x1;
  assign n938 = ~x2 & ((~x1 & ((x6 & ~x7 & (x0 ^ ~x5)) | (~x0 & x5 & (~x6 | x7)))) | (~x6 & x7 & ~x0 & x5));
  assign n939 = (x1 | ((~x0 | (x5 ? x7 : (x6 | ~x7))) & (~x5 | (~x6 ^ ~x7)) & (~x6 | x7 | x0 | x5))) & (x0 | ((~x5 | ((x6 | ~x7) & (~x1 | ~x6 | x7))) & (~x1 | x5 | (~x6 ^ ~x7))));
  assign n940 = ((x6 ^ x7) | ((~x3 | x5 | x0 | ~x1) & (~x0 | x1 | (~x3 ^ ~x5)))) & (~x3 | ((x0 | ~x1 | ~x5 | ~x6 | x7) & (~x0 | x1 | x5 | x6 | ~x7))) & (~x0 | ~x1 | x3 | (~x5 ^ (~x6 & x7)));
  assign z032 = ~n946 | n942 | (~n945 & n947 & x4 & ~x6);
  assign n942 = ~x2 & ((~x4 & ~n944) | (n586 & n943));
  assign n943 = ~x7 & x6 & x4 & x5;
  assign n944 = (~x1 | x5 | ((~x0 | ~x3 | (~x6 ^ x7)) & (~x6 | ~x7 | x0 | x3))) & (x0 | x1 | x3 | ~x5 | x6 | x7);
  assign n945 = ~x1 ^ ~x7;
  assign n946 = (x0 & (((x2 | x3) & (x1 | (~x6 & ~x7))) | (x6 & x7) | (x1 & ~x6 & ~x7))) | (~x0 & ((~x1 & ((~x6 & x7) | (~x2 & ~x3 & ~x7))) | (x6 & ~x7) | (~x6 & x7 & ~x2 & ~x3))) | (x6 & ((x1 & x7) | (~x1 & ~x2 & ~x3 & ~x7)));
  assign n947 = ~x3 & ~x0 & ~x2;
  assign z033 = n951 | ~n953 | (~x2 & ~n950) | (n949 & ~n952);
  assign n949 = x6 & ~x2 & ~x3;
  assign n950 = (x4 | ~x5 | x7 | x0 | x1 | x3) & (~x0 | x5 | ((x1 | x3 | ~x4 | ~x7) & (~x1 | ~x3 | x4 | x7)));
  assign n951 = ~x2 & ~x3 & ((~x0 & (x1 ? (~x4 ^ x7) : (x4 & ~x7))) | (~x4 & x7 & x0 & ~x1));
  assign n952 = (x0 | x4 | (x1 ? (~x5 | ~x7) : (x5 | x7))) & (~x0 | x1 | ~x4 | ~x5 | x7);
  assign n953 = (x2 | x3 | x7 | ~x0 | ~x1) & ((~x2 & ~x3) | ((x1 | x7) & (x0 | ~x1 | ~x7)));
  assign z035 = ~x2 & (n955 | ~n956 | ~n960);
  assign n955 = ~x0 & ~x4 & (x1 ? (x3 & ~x5) : (~x3 & x5));
  assign n956 = n959 & (~n957 | ~n586) & (~n698 | ~n958);
  assign n957 = x6 & x4 & x5;
  assign n958 = ~x3 & ~x0 & ~x1;
  assign n959 = x0 ? (x1 | ~x3 | (x4 & x5)) : (x3 | ~x4);
  assign n960 = ~n961 & (~x5 | n906 | n917);
  assign n961 = ~x0 & ~x4 & ((~x1 & ~x3 & ~x5 & x6) | (x5 & ~x6 & x1 & x3));
  assign z036 = ~n964 | ~n963 | (n723 & n665 & ~n917);
  assign n963 = x0 | (x2 ? (x3 | (~x1 & x4)) : (~x3 | (x1 & ~x4)));
  assign n964 = n966 & (~x3 | ((~n957 | ~n534) & (~n965 | ~n750)));
  assign n965 = ~x6 & ~x4 & ~x5;
  assign n966 = x1 | ~x2 | ((x3 | ~x4 | x5) & (~x0 | (x3 & x4)));
  assign z037 = n968 | n970 | n972 | ~n973 | (x3 & ~n971);
  assign n968 = ~x1 & ((x4 & ~n969) | (~x4 & ~x5 & ~n620 & n947));
  assign n969 = (x7 | ((~x3 | x5 | x6 | x0 | ~x2) & (~x0 | x3 | ~x6 | (~x2 ^ x5)))) & (~x5 | x6 | ~x7 | ~x0 | x2);
  assign n970 = ~x0 & ((~x1 & ~x2 & x3 & x4 & ~x5) | (x2 & ((x1 & ~x4 & (~x3 ^ x5)) | (x4 & x5 & ~x1 & ~x3))));
  assign n971 = (~x4 | ~x5 | ~x6 | ~x0 | x1 | x2) & (x0 | ((x1 | x2 | ~x4 | ~x5 | x6) & (~x1 | ~x2 | x4 | x5 | ~x6)));
  assign n972 = ~x1 & (x0 ? (x2 & (x3 ^ ~x4)) : (x3 & ~x4));
  assign n973 = n977 & (n974 | ~n975) & (x6 | ~n610 | n976);
  assign n974 = (x4 | ~x5 | ~x6 | ~x7) & (x5 | x6 | x7 | x3 | ~x4);
  assign n975 = ~x2 & ~x0 & x1;
  assign n976 = (~x4 | x5 | x1 | ~x2) & (x4 | ~x5 | ~x1 | x2);
  assign n977 = ~x1 | ((x0 | ~x3 | ~x4) & (x3 | x4 | x5 | ~x0 | x2));
  assign z038 = ~n982 | (x4 & (~n981 | (x2 ? ~n979 : ~n980)));
  assign n979 = (x1 | ((x0 | ~x3 | x5 | x6 | ~x7) & (~x0 | ~x6 | (x3 ? (~x5 | x7) : (x5 | ~x7))))) & (x0 | ~x1 | x5 | x7 | (~x3 ^ x6));
  assign n980 = (~x5 | x6 | ~x7 | ~x0 | x1 | ~x3) & (x3 | ((~x0 | ~x5 | (x1 ? (x6 | x7) : (~x6 | ~x7))) & (x0 | ~x1 | x5 | x6 | ~x7)));
  assign n981 = (x0 | ((~x3 | x5 | ~x6 | x1 | ~x2) & (~x1 | x6 | (x2 ? (x3 | x5) : (~x3 | ~x5))))) & (x1 | ~x3 | ~x5 | ((x2 | ~x6) & (~x0 | ~x2 | x6)));
  assign n982 = ~n984 & n987 & ~n988 & (~x3 | ~n670 | ~n983);
  assign n983 = ~x6 & ~x4 & x5;
  assign n984 = ~x4 & ((n537 & n985 & n924) | (~x1 & ~n986));
  assign n985 = x3 & x5;
  assign n986 = (x7 | ((~x3 | x5 | x6 | ~x0 | ~x2) & (x0 | ~x5 | (x2 ? (x3 | x6) : (~x3 | ~x6))))) & (x0 | x2 | x3 | x5 | ~x6 | ~x7);
  assign n987 = x1 ? ((x2 | ~x4 | (x0 ? (x3 | x5) : (~x3 ^ x5))) & (x4 | ~x5 | x0 | ~x2)) : (x5 ? ((~x2 | x3 | ~x4) & (x0 | (x2 ? ~x4 : (x3 | x4)))) : ((~x0 | ((x3 | x4) & (~x2 | ~x3 | ~x4))) & (x4 | (~x2 ^ x3))));
  assign n988 = ~n989 & ((x0 & ~x2 & ~x3 & ~x4 & x5) | (~x0 & ~x5 & (x2 ? (x3 & ~x4) : (~x3 & x4))));
  assign n989 = ~x1 ^ ~x6;
  assign z039 = n996 | (x2 ? (~n994 | ~n998) : (~n991 | ~n995));
  assign n991 = x0 ? (x1 | n993) : n992;
  assign n992 = (x1 | ~x3 | ~x6 | (x4 ? (x5 | x7) : (~x5 | ~x7))) & (x3 | ((x6 | x7 | ~x4 | ~x5) & (x5 | ((~x6 | ~x7 | x1 | x4) & (~x1 | (x4 ? (x6 | ~x7) : (~x6 | x7)))))));
  assign n993 = (x4 | x5 | ~x6 | x7) & (~x4 | ~x5 | ~x7 | (~x3 ^ x6));
  assign n994 = (x1 | ((~x0 | (x3 ? (~x4 | x5) : (~x5 | x6))) & (x3 | ~x4 | ~x5 | x6) & (~x3 | ((x5 | ~x6) & (~x5 | x6 | x0 | x4))))) & (x0 | (x3 ? (x5 | ~x6) : (~x5 | (x6 ? x4 : ~x1))));
  assign n995 = (x3 | ((x0 | ((~x4 | x5 | ~x6) & (~x5 | x6 | x1 | x4))) & (~x1 | ((x4 | x5 | x6) & (~x0 | ~x5 | ~x6))))) & (x1 | ((~x0 | ((x5 | x6) & (x4 | ~x5 | ~x6))) & (~x3 | ((~x4 | ~x5 | ~x6) & (x0 | x4 | x5))))) & (x0 | ~x3 | ((~x4 | ~x5 | ~x6) & (x5 | x6)));
  assign n996 = ~n824 & ~n997;
  assign n997 = (x3 | ~x4 | x6 | ~x0 | ~x1 | x2) & (x0 | x4 | ((~x3 | ~x6 | ~x1 | x2) & (x1 | ~x2 | x3 | x6)));
  assign n998 = (x7 | ((~n732 | n1000) & (~x5 | n999))) & n1001 & (x5 | ~x7 | n999);
  assign n999 = (~x3 | x4 | x6 | ~x0 | x1) & (x0 | ~x4 | (x1 ? (x3 | ~x6) : (~x3 | x6)));
  assign n1000 = (~x1 | x4 | x5 | x6) & (x1 | ~x4 | ~x5 | ~x6);
  assign n1001 = (~x0 | x1 | (x3 ? ~n587 : (~x6 | n1002))) & (x0 | ~x1 | ~x3 | x6 | n1002);
  assign n1002 = x4 ? (x5 | ~x7) : (~x5 | x7);
  assign z040 = ~n1006 | ~n1011 | (x0 ? ~n1004 : ~n1005);
  assign n1004 = (x1 | ((x6 | x7 | x2 | x4) & (~x3 | ((~x2 | x4 | (~x6 ^ x7)) & (x2 | ~x4 | ~x6 | x7))))) & (~x4 | x6 | ~x7 | ~x1 | x2 | x3);
  assign n1005 = (~x7 | ((~x2 | ((~x4 | ~x6 | ~x1 | x3) & (x1 | x6 | (~x3 ^ ~x4)))) & (~x1 | x2 | (x3 ? (x4 | ~x6) : (~x4 | x6))))) & (x3 | x7 | ((~x4 | x6 | ~x1 | ~x2) & (x1 | ~x6 | (~x2 ^ x4))));
  assign n1006 = (n1007 | n1009) & (x0 | n1008) & (~x0 | x4 | n1010);
  assign n1007 = x3 ? (x5 | x6) : (~x5 | ~x6);
  assign n1008 = x2 ? ((x6 | ((~x4 | x5 | x1 | x3) & (~x1 | ~x5 | (~x3 ^ ~x4)))) & (~x3 | x4 | ~x6 | (x1 & x5))) : (x1 ? (x5 | ((x4 | x6) & (~x3 | ~x4 | ~x6))) : (~x3 | ~x5 | (x4 ^ x6)));
  assign n1009 = (x0 | x1 | x2 | x4) & (~x0 | (x1 ? (x2 | x4) : (~x2 | ~x4)));
  assign n1010 = (~x1 | x2 | x3 | x5 | ~x6) & (x1 | (x2 ? (x3 | x6) : (~x5 | ~x6)));
  assign n1011 = x7 ? (~n1017 & ~n1018 & (x3 | n1016)) : n1012;
  assign n1012 = (~x2 | n1015) & (x2 | n1013) & (n783 | n1014);
  assign n1013 = (~x4 | x5 | ((x0 | (x1 ? (x3 | ~x6) : (~x3 | x6))) & (x3 | ~x6 | ~x0 | x1))) & (x4 | ~x5 | x6 | x0 | x3);
  assign n1014 = (x2 | x3 | x5 | ~x0 | ~x1) & (x0 | ~x3 | (x1 ? (x2 | ~x5) : (~x2 | x5)));
  assign n1015 = ((x3 ^ x5) | ((x4 | ~x6 | x0 | ~x1) & (~x4 | x6 | ~x0 | x1))) & (x0 | x1 | x3 | ~x4 | ~x5 | x6);
  assign n1016 = (x0 | ((x5 | ~x6 | x2 | x4) & (~x2 | ((~x5 | ~x6 | x1 | ~x4) & (x5 | x6 | ~x1 | x4))))) & (x1 | x2 | (x4 ? (~x5 | (~x0 & x6)) : (x5 | ~x6)));
  assign n1017 = ~n627 & ((~x0 & x3 & (x1 ? (x2 & ~x6) : (~x2 & x6))) | (x0 & ~x1 & x2 & ~x3 & x6));
  assign n1018 = n1021 & (n1020 | (~x2 & ~n1019));
  assign n1019 = x4 ? (~x5 | x6) : (x5 | ~x6);
  assign n1020 = x6 & x5 & x2 & x4;
  assign n1021 = x3 & x0 & ~x1;
  assign z041 = ~n1025 | (~x0 & (n1024 | (x3 & ~n1023)));
  assign n1023 = (~x5 | ((x7 | ((x6 | (x1 ? (x2 ^ ~x4) : (x2 | x4))) & (x1 | ~x2 | ~x4 | ~x6))) & (x2 | ~x6 | ~x7 | (x1 ^ x4)))) & (x2 | x5 | ((x6 | ~x7 | x1 | ~x4) & (~x1 | x4 | (x6 ^ x7))));
  assign n1024 = ~x5 & n563 & (x1 ? (~x4 & n537) : (x4 & ~n662));
  assign n1025 = n1029 & (~n738 | n1028) & (x2 ? n1027 : n1026);
  assign n1026 = x4 ? (x1 ? (x5 | ((x3 | ~x7) & (x0 | ~x3 | x7))) : (x0 ? ((x5 | x7) & (~x3 | ~x5 | ~x7)) : (~x5 | (~x3 ^ x7)))) : ((x5 | ((~x0 | (x1 ? (~x3 | x7) : ~x7)) & (x1 | x3 | ~x7) & (x0 | x7 | (x1 ^ ~x3)))) & (~x1 | ~x5 | (x0 ? (x3 | x7) : ~x7)));
  assign n1027 = x0 ? (x1 | (((~x3 ^ ~x7) | (~x4 ^ ~x5)) & (~x4 | x5 | (~x3 ^ x7)))) : (x3 ? (x1 ? (x4 ? (~x5 | x7) : (x5 ^ x7)) : (x4 ? (x5 | ~x7) : (~x5 | x7))) : ((~x1 | ((x5 | ~x7) & (x4 | ~x5 | x7))) & (x4 | x5 | ~x7) & (x1 | ~x4 | (x5 ^ x7))));
  assign n1028 = (~x4 | ((x2 | ~x6 | (x5 ? x3 : ~x7)) & (~x2 | ~x3 | ~x5 | x6 | x7))) & (~x2 | x3 | x4 | ~x5 | (x6 ^ x7));
  assign n1029 = x6 ? (x7 | (n1030 & (x2 | ~x5 | n1031))) : ((~x7 | n1030) & (~x2 | n1031 | (x5 ^ x7)));
  assign n1030 = ((x1 ^ x4) | ((~x3 | x5 | x0 | ~x2) & (x3 | ~x5 | ~x0 | x2))) & (x3 | x4 | x5 | ~x0 | ~x1 | x2);
  assign n1031 = (x0 | x3 | (x1 ^ x4)) & (~x3 | x4 | ~x0 | x1);
  assign z042 = ~n1040 | (x1 & ~n1039) | (x5 & ~n1033) | (~x5 & ~n1036);
  assign n1033 = (x0 | n1034) & (~n1035 | (x2 ? ~n544 : n662));
  assign n1034 = (~x2 | ((~x7 | (x1 ? (x3 ? (x4 | x6) : (~x4 | ~x6)) : (x3 ? (~x4 | x6) : (x4 | ~x6)))) & (x1 | x3 | ~x4 | ~x6 | x7))) & (x1 | x2 | x3 | x4 | x6 | ~x7);
  assign n1035 = x4 & ~x3 & x0 & ~x1;
  assign n1036 = x4 ? n1038 : n1037;
  assign n1037 = (x6 | (x0 ? (~x3 | (x1 ? (x2 | x7) : (~x2 | ~x7))) : (x3 | (x1 ? (~x2 | x7) : ~x7)))) & (x2 | ~x6 | ((x0 | (x1 ? (x3 | ~x7) : (~x3 | x7))) & (~x0 | x1 | x3 | x7)));
  assign n1038 = (~x0 | x1 | x2 | x3 | ~x6 | ~x7) & (x0 | ((~x1 | ~x2 | x3 | x6 | ~x7) & (x1 | ((~x6 | ~x7 | x2 | ~x3) & (x6 | x7 | ~x2 | x3)))));
  assign n1039 = (~x0 | x2 | x3 | x4 | x5 | ~x6) & (x0 | ((~x5 | x6 | x3 | x4) & (x5 | ((~x2 | ((~x4 | ~x6) & (~x3 | x4 | x6))) & (x4 | ~x6 | x2 | ~x3)))));
  assign n1040 = ~n1043 & ~n1044 & (n1041 | n1042) & (x1 | n1045);
  assign n1041 = x4 ^ ~x6;
  assign n1042 = (x1 | ((x3 | ~x5 | x7 | x0 | x2) & (~x0 | ~x2 | (x3 ? (~x5 | ~x7) : (x5 | x7))))) & (x0 | ~x1 | ~x5 | (x2 ? (~x3 | x7) : (x3 | ~x7)));
  assign n1043 = ~n850 & ((~x0 & ~x1 & x2 & x3 & ~x7) | (~x2 & ((x3 & ~x7 & ~x0 & x1) | (x0 & (x1 ? (~x3 & ~x7) : (x3 & x7))))));
  assign n1044 = ~n846 & ((~x2 & (x1 ? (x4 & (~x0 | ~x3)) : (x3 & ~x4))) | (~x1 & ((x2 & x3 & x4) | (x0 & ~x3 & ~x4))));
  assign n1045 = (x5 | ~x6 | ((~x2 | ~x3 | x4) & (x0 | (x2 ? x4 : (x3 | ~x4))))) & (~x4 | ~x5 | x6 | (x2 ^ ~x3));
  assign z043 = n1047 | n1050 | ~n1054 | (~n800 & ~n1053);
  assign n1047 = x6 & ((n664 & ~n1049) | (~x1 & ~n1048));
  assign n1048 = (~x2 | ((~x5 | ~x7 | x3 | ~x4) & (~x3 | (x0 ? (x4 ? (x5 | x7) : (~x5 | ~x7)) : (x5 | (x4 ^ x7)))))) & (x0 | x3 | x4 | ~x5 | ~x7) & (x2 | ((x0 | ((x5 | x7 | x3 | x4) & (~x5 | ~x7 | ~x3 | ~x4))) & (~x4 | ~x7 | ~x0 | x3)));
  assign n1049 = (x3 | ((x2 | (x4 ? (x5 | x7) : (~x5 | ~x7))) & (~x2 | ~x4 | ~x5 | ~x7))) & (~x2 | ~x3 | x4 | (~x5 ^ ~x7));
  assign n1050 = ~x6 & (x1 ? ~n1051 : ~n1052);
  assign n1051 = (x2 | ((x5 | ((x4 | (x0 ? (~x3 ^ ~x7) : (~x3 | x7))) & (~x4 | x7 | x0 | x3))) & (~x4 | ~x5 | ~x7 | x0 | x3))) & (x0 | ~x2 | ((x3 | ~x4 | ~x5 | x7) & (~x3 | ((~x5 | ~x7) & (~x4 | x5 | x7)))));
  assign n1052 = (~x4 & (x0 ? (x3 ? x2 : x7) : (~x3 & ~x7))) | (x7 & (~x5 | (x2 & ~x3) | (x3 & ((~x2 & x4) | (~x0 & (~x2 | x4)))))) | (x5 & ~x7) | (x2 & ~x3 & x4);
  assign n1053 = (x2 | ((~x6 | ((~x1 | x3 | (x0 ^ x4)) & (~x3 | ((x1 | ~x4) & (x0 | (x1 & ~x4)))))) & (x0 | x1 | ~x3 | ~x4))) & (x3 | ((x1 | ((~x2 | x4 | x6) & (~x0 | (~x4 ^ x6)))) & (x4 | x6 | x0 | ~x2)));
  assign n1054 = (x0 | n1057) & (n620 | n1056) & (~x0 | n1055);
  assign n1055 = (x2 | x5 | ((~x1 | x3 | (~x4 ^ x6)) & (x4 | ~x6 | x1 | ~x3))) & (x4 | ~x5 | x6 | x1 | ~x2 | ~x3);
  assign n1056 = (x4 | ((~x0 | ((x3 | ~x5 | ~x1 | x2) & (~x3 | x5 | x1 | ~x2))) & (x0 | ~x1 | x2 | ~x3 | ~x5))) & (x0 | ~x2 | ~x4 | ((x3 | x5) & (x1 | ~x3 | ~x5)));
  assign n1057 = (x3 | (x1 ? (x4 | (x2 ? (~x5 | ~x6) : (x5 | x6))) : (~x4 | (x2 ? (~x5 | x6) : (x5 | ~x6))))) & (~x1 | ~x3 | x5 | (x2 ? (~x4 | ~x6) : (~x4 ^ x6)));
  assign z044 = n1059 | ~n1061 | (x0 ? ~n1067 : ~n1066);
  assign n1059 = x4 & ((n537 & n916 & n924) | (~x6 & ~n1060));
  assign n1060 = (x3 | ~x5 | x7 | x0 | ~x1 | ~x2) & (x1 | ((x0 | ~x2 | ~x3 | ~x5 | x7) & (x5 | ((x3 | ~x7 | x0 | ~x2) & (x2 | (x0 ? (x3 ^ x7) : (~x3 | x7)))))));
  assign n1061 = ~n1064 & ((x4 & (~x6 | n1065)) | (~x4 & x6 & n1062) | (~x6 & n1063 & n1065));
  assign n1062 = (x2 | ((~x0 | ((~x1 | x5 | x7) & (~x5 | ~x7 | x1 | x3))) & (x0 | ~x5 | ((x3 | x7) & (x1 | ~x3 | ~x7))) & (x5 | x7 | ~x1 | ~x3))) & (x0 | ~x2 | ((~x5 | x7 | ~x1 | ~x3) & (x1 | x5 | (x3 ^ x7))));
  assign n1063 = (~x0 | x1 | x2 | x3 | x5 | ~x7) & (x0 | ~x2 | ((x1 | ~x5 | (x3 ^ x7)) & (x5 | x7 | ~x1 | ~x3)));
  assign n1064 = ~n662 & (x0 ? ((x3 & ~x4 & ~x1 & x2) | (x1 & ~x2 & ~x3 & x4)) : ((x1 & ~x2 & (x3 ^ ~x4)) | (~x3 & x4 & ~x1 & x2)));
  assign n1065 = (~x5 | ((x0 | ~x1 | ~x2 | x3 | ~x7) & (x2 | ((~x0 | (x1 ? (x3 | x7) : (~x3 | ~x7))) & (~x3 | x7 | x0 | ~x1))))) & (x1 | x5 | ((~x0 | ~x2 | (x3 ^ x7)) & (~x3 | ~x7 | x0 | x2)));
  assign n1066 = x2 ? (x4 ? ((~x3 | x6 | ~x7) & (~x1 | ((x6 | ~x7) & (~x3 | ~x6 | x7)))) : ((~x6 | (x1 ? (~x3 ^ ~x7) : (~x3 | x7))) & (x6 | ~x7 | x1 | x3))) : (x4 ? ((x3 | ~x6 | x7) & (x1 | ((~x6 | x7) & (x3 | x6 | ~x7)))) : ((x1 | (x3 ? (x6 | x7) : (~x6 | ~x7))) & (~x1 | ~x3 | x6 | ~x7)));
  assign n1067 = (x3 | ((~x1 | x2 | x4 | x6 | ~x7) & (x1 | (x2 ? (x4 ? (x6 | ~x7) : ~x6) : (x4 ? ~x6 : (x6 | x7)))))) & (x1 | ~x3 | x7 | (x2 ? (~x4 | ~x6) : (~x4 ^ x6)));
  assign z045 = ~n1071 | (~x0 & ((x5 & ~n1069) | (x4 & ~x5 & ~n1070)));
  assign n1069 = (x1 | ~x3 | ((x6 | ~x7 | x2 | ~x4) & (~x2 | x4 | ~x6 | x7))) & (x3 | ~x4 | ~x6 | x7) & (~x1 | ((~x2 | ~x4 | ((~x6 | x7) & (x3 | x6 | ~x7))) & (x2 | x3 | x4 | x6 | x7)));
  assign n1070 = (~x3 | ((~x6 | x7 | ~x1 | ~x2) & (x6 | ~x7 | x1 | x2))) & (x1 | ~x2 | x3 | (~x6 ^ x7));
  assign n1071 = ~n1073 & n1076 & ((x7 & (~x6 | n1072)) | (n1075 & (n1072 | (x6 & ~x7))));
  assign n1072 = (x3 | ((~x4 | ((~x0 | x2 | (x1 ^ x5)) & (x1 | ~x2 | ~x5) & (x0 | (x1 ? (~x2 | x5) : ~x5)))) & (~x0 | x4 | x5 | (x1 ^ ~x2)))) & (x0 | ~x3 | (x1 ? ((~x4 | ~x5) & (x2 | x4 | x5)) : (~x4 | x5)));
  assign n1073 = x0 & ((~x1 & ~n1074) | (n698 & n811));
  assign n1074 = (~x4 | ~x5 | ((~x3 | ~x6 | x7) & (~x2 | x6 | ~x7))) & (~x3 | x4 | x5 | ((x6 | ~x7) & (x2 | ~x6 | x7)));
  assign n1075 = (x4 | ((x1 | ((x3 | x5 | x0 | ~x2) & (~x5 | ((x2 | ~x3) & (~x0 | (x2 & ~x3)))))) & (x0 | ~x1 | (x2 ? (~x3 ^ x5) : (x3 | x5))))) & (x3 | ~x4 | x5 | ~x0 | x1 | ~x2);
  assign n1076 = (~n694 | ~n1079) & (~x7 | n1077) & (x0 | n1078);
  assign n1077 = x1 ? ((~x0 | x2 | x3 | x4 | ~x5) & (x0 | ((~x3 | x4 | ~x5) & (~x4 | x5 | x2 | x3)))) : (x5 ? ((x0 | ((x3 | x4) & (~x2 | ~x3 | ~x4))) & (x3 | ((~x2 | x4) & (~x0 | x2 | ~x4)))) : (x0 ? ((~x3 | ~x4) & (x2 | x3 | x4)) : (~x3 | x4)));
  assign n1078 = (x2 | ((x5 | ~x6 | x7 | x1 | x3) & (~x1 | ((~x6 | x7 | ~x3 | x5) & (x3 | ~x5 | x6 | ~x7))))) & (x5 | x6 | ~x7 | ~x1 | ~x2 | x3);
  assign n1079 = ~x7 & x6 & ~x3 & ~x5;
  assign z046 = n1081 | ~n1085 | ~n1089 | (~n620 & ~n1084);
  assign n1081 = x0 & ((~x1 & ~n1083) | (n1082 & n559));
  assign n1082 = ~x3 & x1 & ~x2;
  assign n1083 = x6 ? (~x7 | ((x4 | ((x3 | ~x5) & (x2 | (x3 & ~x5)))) & (~x2 | ~x4 | x5))) : (x7 | ((x2 | ~x3 | ~x4 | ~x5) & (~x2 | (x3 ? (x4 | x5) : (~x4 | ~x5)))));
  assign n1084 = (x4 | ((x5 | ((~x0 | ((x2 | x3) & (x1 | ~x2 | ~x3))) & (x2 | (x1 ^ x3)) & (x0 | (x2 ? ~x1 : ~x3)))) & (~x0 | x1 | ~x5 | (~x2 ^ x3)))) & (x0 | ~x4 | ~x5 | (x1 & (~x2 | ~x3)));
  assign n1085 = (n1041 | n1087) & (x4 | n1086) & (x2 | ~x4 | n1088);
  assign n1086 = (x1 | ((x0 | x2 | x3 | ~x5 | ~x6) & (~x0 | x5 | x6 | (~x2 ^ x3)))) & (x0 | ~x1 | ~x6 | (x2 ? (~x3 | ~x5) : (x3 | x5)));
  assign n1087 = (~x5 | (x0 ? (x1 ? (x2 | x3) : (~x2 | ~x3)) : (~x1 | (~x2 ^ x3)))) & (x0 | x1 | ~x2 | x5);
  assign n1088 = (x0 | ~x1 | x3 | ~x5 | x6) & (~x0 | x1 | x5 | (x3 ^ x6));
  assign n1089 = (n662 | n1090) & (x0 | (x2 ? n1092 : n1091));
  assign n1090 = (x2 | ((x0 | ~x1 | ~x3 | ~x4 | x5) & (x3 | ((~x0 | ~x4 | (x1 ^ ~x5)) & (x4 | ~x5 | x0 | ~x1))))) & (~x3 | x4 | ~x5 | x0 | x1 | ~x2);
  assign n1091 = (x5 | ((~x6 | ~x7 | x1 | x4) & (~x1 | ((~x6 | ~x7 | x3 | ~x4) & (~x3 | x4 | x6 | x7))))) & (x1 | ((~x4 | x6 | x7) & (~x3 | x4 | ~x6 | ~x7)));
  assign n1092 = (~x6 | ~x7 | ((~x1 | ~x3 | x4 | x5) & (x1 | ~x5 | (~x3 ^ ~x4)))) & (~x1 | ~x4 | x6 | x7 | (~x3 & x5));
  assign z047 = n1095 | ~n1096 | ~n1103 | (~x0 & ~n1094);
  assign n1094 = (x3 | ((~x4 | ((x1 | x7 | (x2 ^ x5)) & (~x5 | ~x7 | ~x1 | x2))) & (~x1 | x4 | ~x5 | (x2 ^ x7)))) & (~x1 | ~x3 | x5 | x7 | (~x2 ^ x4));
  assign n1095 = ~x1 & ((~x5 & x7 & ~x0 & x2) | (x3 & x5 & (x0 ? (x2 ^ ~x7) : (x2 & ~x7))));
  assign n1096 = n1098 & (n912 | n1097);
  assign n1097 = x2 ? ((~x3 & ~x4) | (x0 ? (x1 | x7) : (~x1 | ~x7))) : ((x0 | (x1 ? (x7 | (~x3 ^ x4)) : (~x7 | (x3 & x4)))) & (x4 | ~x7 | x1 | x3));
  assign n1098 = ~n1101 & (~n720 | ~n686) & (n1099 | n1100 | ~n1102);
  assign n1099 = x3 ^ ~x4;
  assign n1100 = x1 ^ ~x7;
  assign n1101 = x1 & ((~x0 & ((x5 & x7 & ~x2 & x3) | (~x5 & ~x7 & x2 & ~x3))) | (~x3 & x5 & x7 & x0 & ~x2));
  assign n1102 = ~x5 & x0 & ~x2;
  assign n1103 = (n846 | n1104) & (x1 | n1105);
  assign n1104 = x0 ? (x1 | (x2 ? (x3 | ~x7) : (x3 ? (~x4 | ~x7) : x7))) : (x1 ? ((x4 | ~x7 | x2 | x3) & (~x4 | x7 | ~x2 | ~x3)) : (x7 | (x2 ? (x3 | x4) : ~x3)));
  assign n1105 = (n1107 | n1108) & (~x0 | ~n665 | ~n565) & (x0 | n1106);
  assign n1106 = (x5 | ~x6 | x7 | x2 | x3 | x4) & (~x2 | ~x4 | ((x6 | x7 | x3 | x5) & (~x6 | ~x7 | ~x3 | ~x5)));
  assign n1107 = x3 ? (x5 | ~x7) : (~x5 | x7);
  assign n1108 = (~x0 | ~x2 | x4 | x6) & (x0 | x2 | ~x4 | ~x6);
  assign z048 = ~n1111 | n1124 | (x6 ? (x7 ? ~n1110 : ~n1125) : (x7 ? ~n1125 : ~n1110));
  assign n1110 = (x1 | ((~x4 | (x0 ? (x2 | ~x3) : (x2 ? (~x3 | ~x5) : (x3 | x5)))) & (~x0 | ((x2 | ~x3 | ~x5) & (x4 | x5 | ~x2 | x3))))) & (x0 | ((x4 | ~x5 | x2 | x3) & (~x1 | (x2 ? (~x3 ^ x4) : (x3 | x4)))));
  assign n1111 = ~n1113 & ~n1114 & ~n1118 & (~n534 | ~n1112);
  assign n1112 = ~x6 & ~x5 & x3 & ~x4;
  assign n1113 = ~x1 & ((~x0 & x2 & x3 & ~x4 & ~x6) | (x6 & ((x3 & ~x4 & ~x0 & ~x2) | (x0 & ~x3 & (~x2 ^ x4)))));
  assign n1114 = ~n1115 & ((x4 & n598 & ~n1116) | (x0 & ~x4 & ~n1117));
  assign n1115 = x3 ^ ~x5;
  assign n1116 = x2 ^ ~x6;
  assign n1117 = x1 ? (x2 | x6) : (~x2 | ~x6);
  assign n1118 = n670 & n1122 & ((n1119 & n1121) | (n1120 & n1123));
  assign n1119 = x0 & x4;
  assign n1120 = ~x5 & x6;
  assign n1121 = x5 & ~x6;
  assign n1122 = ~x3 & x7;
  assign n1123 = ~x0 & ~x4;
  assign n1124 = x1 & ((~x0 & ((~x2 & x3 & x4 & ~x6) | (x2 & (x3 ? (x4 & x6) : (~x4 & ~x6))))) | (~x3 & x4 & ~x6 & x0 & ~x2));
  assign n1125 = x1 ? (x2 | ((x0 | (~x3 ^ x4)) & (x4 | x5 | ~x0 | x3))) : ((~x4 | ((~x3 | ~x5 | x0 | x2) & (~x0 | (x2 ? ~x3 : (x3 | x5))))) & (~x2 | (x0 ? (~x3 | ~x5) : (x3 | (x4 & x5)))));
  assign z049 = ~n1128 | n1129 | n1131 | (~x2 & ~n1127);
  assign n1127 = x3 ? (x0 ? (x4 | ((x5 | x7) & (x1 | ~x5 | ~x7))) : (x1 | ~x4 | (x5 ^ x7))) : (x1 ? (x4 | ((x5 | ~x7) & (~x0 | ~x5 | x7))) : (~x4 | ((x5 | ~x7) & (x0 | ~x5 | x7))));
  assign n1128 = (((~x3 | ~x7) & (~x2 | x3 | x7)) | (x0 ? (x1 | ~x4) : (~x1 | x4))) & ((x1 ^ x4) | ((x0 | (~x3 ^ x7)) & (x3 | x7 | ~x0 | x2)));
  assign n1129 = n538 & ~n1130 & (x3 ? (x5 ^ ~x7) : (~x5 ^ ~x7));
  assign n1130 = x0 ^ ~x4;
  assign n1131 = n1132 & (x4 ? (n544 & n738) : (n664 & n543));
  assign n1132 = x5 & ~x2 & ~x3;
  assign z050 = (~n933 & (x0 ? (~x4 ^ ~x5) : (x4 ^ ~x5))) | ~n1135 | (x4 & ~n1134);
  assign n1134 = (x1 | x2 | x3 | (~x0 ^ x5)) & (x0 | ~x1 | (~x2 & ~x3 & x5));
  assign n1135 = (~n677 | ~n921) & (~n670 | ~n1136 | n1137);
  assign n1136 = ~x3 & ~x6;
  assign n1137 = (x5 | ~x7 | x0 | x4) & (~x5 | x7 | ~x0 | ~x4);
  assign z051 = (n1132 & (~n1140 | ~n1141)) | ~n1142 | (~x2 & ~n1139);
  assign n1139 = (~x0 | x1 | (~x3 ^ ~x5)) & (~x1 | (x0 ? (x3 | ~x5) : (~x3 | x5)));
  assign n1140 = (x0 | ~x1 | x4 | ~x6 | x7) & (~x0 | x1 | ~x4 | x6 | ~x7);
  assign n1141 = (~x0 | x1 | ~x4 | ~x6) & (x0 | ~x1 | x4 | x6);
  assign n1142 = (x1 | ~x2 | ~x5) & (x0 | (x1 ? (x5 | (~x2 & (x3 | ~x4))) : ~x5));
  assign z052 = ~x6 & (~n1145 | (n677 & n1144));
  assign n1144 = x7 & ~x5 & ~x3 & ~x4;
  assign n1145 = (x0 & x1 & (x2 | (x3 & (x4 | x5)))) | (~x0 & ~x1 & ~x2 & ~x3 & ~x4 & ~x5);
  assign z053 = ~x7 & (~n1145 | (n677 & n921));
  assign z054 = ~x0 & (~n933 | ~n1149 | (n730 & n1148 & ~n1150));
  assign n1148 = ~x2 & ~x4;
  assign n1149 = x1 | x2 | x3 | (~x4 & ~x5 & ~x6);
  assign n1150 = x1 ? (~x3 | x7) : (x3 | ~x7);
  assign z055 = n1157 | ~n1158 | (~x6 & (n1152 | n1155));
  assign n1152 = n605 & (x0 ? (~x2 & n1153) : (~x5 & ~n1154));
  assign n1153 = ~x7 & x4 & x5;
  assign n1154 = x2 ? (~x4 | x7) : (x4 | ~x7);
  assign n1155 = n924 & n1156 & n650;
  assign n1156 = ~x5 & x7;
  assign n1157 = ~x2 & ((~x0 & ~x4 & x5 & (~x1 ^ x3)) | (~x3 & x4 & ~x5 & x0 & ~x1));
  assign n1158 = (x0 | (x2 ? (~x1 & (x3 | x4)) : ((~x3 | ~x4) & (x1 | (~x3 & ~x4))))) & ~n1159 & (x2 | x3 | x4 | ~x0 | x1);
  assign n1159 = x6 & n597 & n897 & (x1 ^ ~x3);
  assign z056 = ~n1162 | ~n1164 | ~n1165 | (~x3 & ~n1161);
  assign n1161 = (x1 | ((~x4 | x5 | ~x6 | x0 | ~x2) & (~x0 | ~x5 | (x2 ? (x4 | x6) : (~x4 | ~x6))))) & (x0 | ~x1 | x2 | x4 | ~x5 | x6);
  assign n1162 = (x1 | (x0 ? (x2 | (~x3 & ~n1163)) : (~x2 | ~x3))) & (x0 | ((~x2 | ~x3 | x4) & (~x1 | (x2 ? x3 : (~x3 | ~x4)))));
  assign n1163 = x7 & ~x6 & x4 & x5;
  assign n1164 = ~n664 | ((~x3 | ~x5 | (x2 ? (~x4 | x6) : x4)) & (x2 | x4 | x5 | (x3 & ~x6)));
  assign n1165 = ~n1167 & (x0 | ((~n808 | n1168) & (~n742 | ~n1166)));
  assign n1166 = x7 & ~x6 & x4 & ~x5;
  assign n1167 = x2 & ((x0 & ~x1 & ~x3 & ~x4 & ~x5) | (~x0 & x4 & (x1 ? (x3 & ~x5) : (~x3 & x5))));
  assign n1168 = (~x6 | x7 | x3 | ~x5) & (x6 | ~x7 | ~x3 | x5);
  assign z057 = n1174 | ~n1175 | (~x0 & (~n1170 | n1171 | n1173));
  assign n1170 = x2 ? ((~x4 | x5 | ~x6 | x1 | x3) & (~x5 | ((~x1 | (x3 ? (~x4 | ~x6) : (x4 | x6))) & (~x4 | x6 | x1 | ~x3)))) : (x4 | x5 | (x1 ? (~x3 | ~x6) : (~x3 ^ x6)));
  assign n1171 = ~x4 & ((x1 & (x2 ? (~x3 & n1172) : (x3 & n836))) | (~x3 & n836 & ~x1 & ~x2));
  assign n1172 = ~x7 & x5 & x6;
  assign n1173 = x4 & n538 & ((x3 & x5 & x6 & ~x7) | (~x6 & x7 & ~x3 & ~x5));
  assign n1174 = ~x0 & ((~x4 & ((x1 & (x2 ? (~x3 & ~x5) : (x3 & x5))) | (~x1 & ~x2 & ~x3 & x5))) | (~x1 & x2 & x4 & (x3 ^ x5)));
  assign n1175 = ~n1177 & n1178 & (~n1176 | ~n1179) & (~n568 | ~n1180);
  assign n1176 = x2 & x0 & ~x1;
  assign n1177 = ~x1 & ((x2 & x3 & ~x4) | (~x3 & ((~x2 & x4) | (x0 & (~x2 | x4)))));
  assign n1178 = ~x3 | ~x4 | ((x0 | ~x1 | x2) & (~x0 | x1 | ~x2 | x5));
  assign n1179 = x6 & x5 & ~x3 & ~x4;
  assign n1180 = x3 & x2 & x0 & ~x1;
  assign z058 = ~n1187 | (~x1 & (n1183 | ~n1186 | (~x0 & ~n1182)));
  assign n1182 = (~x4 | ((x2 | ~x3 | ~x5 | x6 | x7) & (~x2 | ~x7 | (x3 ? (~x5 | ~x6) : (x5 | x6))))) & (x2 | x3 | x4 | (x5 ? (~x6 | x7) : (x6 | ~x7)));
  assign n1183 = n1119 & ((n871 & n768) | (~x7 & n1184 & ~n1185));
  assign n1184 = ~x2 & ~x5;
  assign n1185 = ~x3 ^ ~x6;
  assign n1186 = x4 ? ((~x0 | ~x3 | (x2 ? (~x5 | ~x6) : (x5 | x6))) & (x0 | ~x2 | x3 | x5 | ~x6)) : (x0 ? (~x2 | (x3 ? (x5 | x6) : (~x5 | ~x6))) : (x2 | ((x5 | ~x6) & (x3 | ~x5 | x6))));
  assign n1187 = n1188 & (~n664 | (n1189 & (x4 | n1190)));
  assign n1188 = (x3 | ((~x0 | ((x2 | x4) & (x1 | ~x2 | ~x4))) & (~x4 | ~x5 | x1 | ~x2) & (~x1 | ((x2 | x4 | x5) & (x0 | ~x2 | ~x4))))) & (x0 | x2 | ~x3 | ~x4 | x5) & (x4 | (x0 ? (x1 | x2) : (~x3 | ((x2 | ~x5) & (x1 | ~x2 | x5)))));
  assign n1189 = (x2 | x3 | x4 | ~x5 | x6) & (~x3 | ((~x2 | (x4 ? (~x5 | ~x6) : (x5 | x6))) & (x5 | ~x6 | x2 | x4)));
  assign n1190 = (x2 | ~x3 | x5 | x6 | ~x7) & (~x6 | ((x2 | x3 | ~x5 | x7) & (~x2 | (x3 ? (x5 | x7) : (~x5 | ~x7)))));
  assign z059 = ~n1196 | (x1 ? ~n1192 : (x5 ? ~n1194 : ~n1195));
  assign n1192 = x0 ? (~n563 | ~n686) : n1193;
  assign n1193 = (~x2 | ((~x3 | x4 | x5 | ~x6 | ~x7) & (x3 | ~x4 | ~x5 | x6 | x7))) & (x2 | ~x3 | x4 | x5 | x6 | ~x7) & (x3 | ((~x6 | ~x7 | x4 | ~x5) & (x2 | x7 | (x4 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n1194 = x2 ? (~x3 | ((~x6 | ~x7 | x0 | ~x4) & (~x0 | (x4 ? (x6 | ~x7) : (~x6 | x7))))) : ((x0 | x3 | x4 | ~x6 | ~x7) & (x6 | ((~x0 | x7 | (~x3 ^ x4)) & (~x4 | ~x7 | x0 | ~x3))));
  assign n1195 = (~x4 | ~x6 | ~x7 | ~x0 | x2 | ~x3) & (x3 | ((x6 | ((~x0 | (x2 ? (x4 | x7) : (~x4 | ~x7))) & (~x4 | ~x7 | x0 | ~x2))) & (x4 | ~x6 | x7 | x0 | ~x2)));
  assign n1196 = ~n1197 & ~n1199 & ~n1200 & (x2 ? n1201 : n1198);
  assign n1197 = x0 & ((x4 & ((x1 & ~x2 & ~x3 & ~x5) | (~x1 & (x2 ? (~x3 & ~x5) : (x3 & x5))))) | (~x1 & ~x2 & ~x4 & ~x5));
  assign n1198 = (~x4 | x5 | ~x6 | ~x0 | x1 | x3) & (x0 | ~x1 | ((x3 | ~x4 | x5 | x6) & (~x3 | x4 | (~x5 ^ x6))));
  assign n1199 = ~n868 & (x0 ? ((~x1 & x2 & x3 & x6) | (x1 & ~x2 & ~x3 & ~x6)) : (~x1 & (x2 ? (~x3 & ~x6) : (x3 & x6))));
  assign n1200 = ~x0 & ((~x1 & ((x3 & ~x4 & x5) | (x4 & ~x5 & ~x2 & ~x3))) | (x2 & ((x1 & ~x3 & x4 & ~x5) | (x3 & ~x4 & x5))) | (x1 & ~x2 & (x3 ? (x4 & x5) : (~x4 & ~x5))));
  assign n1201 = (x1 | (~x3 ^ x6) | (x0 ? (x4 | ~x5) : (~x4 | x5))) & (x0 | ~x1 | ((x5 | x6 | x3 | x4) & (~x5 | ~x6 | ~x3 | ~x4)));
  assign z060 = ~n1211 | (x5 ? ~n1203 : (x1 ? ~n1210 : ~n1209));
  assign n1203 = (n1204 | n1207) & (~x7 | n1206) & (x7 | ~n1205 | n1208);
  assign n1204 = ~x2 ^ ~x4;
  assign n1205 = ~x0 & x6;
  assign n1206 = (x0 | ((x3 | (x1 ? (x2 ? (x4 | ~x6) : (~x4 | x6)) : (x4 | (~x2 ^ x6)))) & (~x2 | ~x3 | (x1 ? (x4 | x6) : (~x4 | ~x6))))) & (x1 | ~x3 | ((x2 | ~x4 | x6) & (~x0 | ~x2 | x4 | ~x6)));
  assign n1207 = (x0 | ~x1 | x3 | x6 | ~x7) & (~x0 | x1 | (x3 ? (x6 | ~x7) : (~x6 | x7)));
  assign n1208 = (~x1 | x2 | ~x3 | ~x4) & (x1 | (x2 ? (~x3 | x4) : (x3 | ~x4)));
  assign n1209 = (x7 | (x0 ? (x3 | (x2 ? (~x4 ^ x6) : (x4 | x6))) : (x2 ? (x3 ? (x4 | x6) : (~x4 | ~x6)) : (x3 ? (x4 | ~x6) : (~x4 | x6))))) & (x3 | x6 | ~x7 | (x0 ? (~x2 ^ x4) : (x2 ^ x4)));
  assign n1210 = (x7 | ((x2 | ((~x4 | x6 | x0 | ~x3) & (~x0 | (x3 ? (x4 | x6) : (~x4 | ~x6))))) & (x0 | ~x2 | ~x6 | (~x3 ^ ~x4)))) & (x4 | x6 | ~x7 | x0 | x2 | ~x3);
  assign n1211 = ~n1214 & ~n1216 & (x0 ? (x1 | n1212) : n1213);
  assign n1212 = (~x2 | ~x3 | x4 | x5 | ~x6) & (x3 | ((x5 | ~x6 | x2 | ~x4) & (~x5 | (x2 ? (~x4 ^ x6) : (x4 | x6)))));
  assign n1213 = (x2 | (x1 ? (~x3 | (x4 ? (~x5 | x6) : ~x6)) : (x3 | (x4 ? (~x5 | x6) : (x5 | ~x6))))) & (x1 | ~x2 | ((~x5 | ~x6 | x3 | ~x4) & (~x3 | (x4 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n1214 = ~n1215 & ((~x2 & (x0 ? (x1 ? (~x3 & ~x4) : (x3 & x4)) : (x1 ? (~x3 & x4) : (x3 & ~x4)))) | (~x0 & x2 & ~x4 & (x1 | ~x3)));
  assign n1215 = x5 ? (x6 | x7) : (~x6 | ~x7);
  assign n1216 = ~n846 & ((x4 & (x0 ? (x1 ? (~x2 & ~x3) : (x2 & x3)) : (x1 ? x2 : (~x2 & x3)))) | (~x2 & ~x4 & (x0 ? (~x1 & x3) : (x1 & ~x3))));
  assign z061 = n1218 | ~n1223 | (~n620 & ~n1222) | (~n662 & ~n1221);
  assign n1218 = ~x2 & ((n544 & ~n1220) | (~x6 & ~n1219));
  assign n1219 = (~x0 | ((x1 | x3 | ~x4 | ~x5) & (~x1 | ~x3 | x4 | x5 | ~x7))) & (x1 | ((~x5 | ~x7 | x3 | ~x4) & (x4 | ((x3 | x5 | ~x7) & (x0 | ~x3 | (x5 ^ x7)))))) & (x0 | ~x1 | ~x5 | (x3 ? (~x4 | ~x7) : (~x4 ^ x7)));
  assign n1220 = (x5 | ((x1 | ~x3 | x4) & (x0 | (x1 ? (x3 | x4) : ~x3)))) & (~x3 | ~x4 | ~x5 | ~x0 | x1);
  assign n1221 = x1 ? ((x2 | ((x3 | x5) & (x0 | ~x3 | ~x5))) & (x0 | x5 | (x3 ? ~x2 : ~x4))) : ((~x0 | ((x3 | x4 | ~x5) & (x2 | ~x3 | x5))) & (x2 | (x3 ? (~x4 | x5) : (x4 | ~x5))) & (~x4 | ~x5 | x0 | x3) & (~x2 | ((x0 | ((~x4 | ~x5) & (x3 | x4 | x5))) & (~x5 | (~x3 ^ x4)))));
  assign n1222 = (x2 | ((~x5 | ((x0 | x1 | ~x3 | ~x4) & (~x0 | x4 | (~x1 ^ x3)))) & (~x4 | x5 | ((x1 | x3) & (x0 | ~x1 | ~x3))))) & (~x3 | x4 | x5 | x0 | x1 | ~x2);
  assign n1223 = ~n1225 & (~x2 | (~n1227 & (n630 | n1224) & n1228));
  assign n1224 = (x1 | ~x3 | ~x4) & (x0 | ~x1 | x3 | x4);
  assign n1225 = ~n1226 & ((x2 & ((~x1 & ~x3 & ~x4) | (~x0 & (x1 ? (x3 & x4) : ~x3)))) | (x1 & ~x2 & ((~x3 & x4) | (~x0 & x3 & ~x4))));
  assign n1226 = x5 ? (~x6 | x7) : (x6 | ~x7);
  assign n1227 = ~n1100 & n732 & x4 & n1120;
  assign n1228 = (~n1229 | ~n1231) & (n906 | n1041 | n1230);
  assign n1229 = x3 & x0 & ~x1;
  assign n1230 = x0 ? (x1 | x5) : (~x1 | ~x5);
  assign n1231 = x7 & ~x6 & ~x4 & x5;
  assign z062 = ~n1238 | (x2 ? (x4 ? ~n1236 : ~n1237) : ~n1233);
  assign n1233 = x4 ? n1235 : n1234;
  assign n1234 = (~x0 & (x1 ? (~x5 & x7) : (x3 ^ x5))) | (x3 & ((x0 & x5) | (x1 & ~x5 & x7))) | (x0 & x1 & (x5 | (~x3 & ~x7))) | (x6 & x7) | (~x7 & (~x6 | (~x3 & x5)));
  assign n1235 = (~x5 | ((x0 | ~x1 | ~x3 | (x6 ^ x7)) & (x7 | ((x1 | x3 | x6) & (~x0 | ((x3 | x6) & (x1 | (x3 & x6)))))))) & (x1 | ~x6 | ~x7 | (x0 ^ x3)) & (x5 | ((x0 | x1 | ~x3 | (~x6 ^ x7)) & (x3 | ((~x6 | ~x7) & (~x1 | x6 | x7)))));
  assign n1236 = ((~x6 ^ x7) | (x0 ? (x1 | (~x3 ^ ~x5)) : (x3 | (~x1 & ~x5)))) & (x0 | ~x3 | ((x5 | x6 | x7) & (x1 | ((x6 | x7) & (x5 | ~x6 | ~x7)))));
  assign n1237 = ((x6 ^ x7) | (x0 ? (x1 | ~x3) : ((x3 | x5) & (~x1 | ~x3 | ~x5)))) & (x1 | ((x0 | x6 | (x3 ? (x5 | ~x7) : x7)) & (~x0 | x3 | ~x5 | ~x6 | x7)));
  assign n1238 = ~n1240 & ~n1242 & ~n1245 & (x2 | n1239);
  assign n1239 = (x1 | ((x0 | ~x3 | x4 | x5 | ~x6) & (x6 | ((x3 | ~x4 | x5) & (~x0 | ((~x4 | x5) & (~x3 | x4 | ~x5))))))) & (x0 | ~x1 | ((x3 | ~x5 | ~x6) & (x5 | x6 | ~x3 | ~x4)));
  assign n1240 = ~n1241 & ((~x0 & x5 & (x1 ? (x2 & x6) : (~x2 & ~x6))) | (x0 & ~x1 & x2 & ~x5 & x6));
  assign n1241 = ~x3 ^ ~x4;
  assign n1242 = ~n783 & (n1244 | (x3 & n616 & ~n1243));
  assign n1243 = x1 ^ ~x5;
  assign n1244 = x5 & ~x3 & ~x2 & x0 & x1;
  assign n1245 = ~x3 & n538 & ((x0 & x4 & x5 & ~x6) | (~x0 & x6 & (x4 ^ x5)));
  assign z063 = ~n1250 | (~x7 & (n1248 | (x6 & ~n1247)));
  assign n1247 = (x0 | ((x3 | ((x1 | (x4 ? x2 : x5)) & (~x2 | (x4 ? ~x1 : x5)))) & (x2 | ~x3 | (x1 ? (x4 ^ x5) : (x4 | ~x5))))) & (x1 | ((~x4 | x5 | ((x2 | ~x3) & (~x0 | ~x2 | x3))) & (~x0 | ~x2 | ((x4 | ~x5) & (~x3 | (x4 & ~x5))))));
  assign n1248 = n534 & n1249;
  assign n1249 = ~x6 & x5 & ~x3 & x4;
  assign n1250 = ~n1253 & n1254 & (n662 | n1251) & (n806 | n1252);
  assign n1251 = ((x4 ^ x5) | ((~x0 | ~x1 | x2 | x3) & (x0 | ~x2 | (~x1 ^ x3)))) & (x1 | (x3 ? ((~x0 | ~x2 | x4 | ~x5) & (~x4 | x5 | x0 | x2)) : (x0 ? (x2 ? (~x4 | x5) : (x4 | ~x5)) : (~x5 | (~x2 ^ x4))))) & (x0 | ~x1 | ~x2 | ~x3 | ~x4 | x5);
  assign n1252 = (~x0 | ~x1 | x2 | x3) & (x0 | x1 | ~x2 | ~x3);
  assign n1253 = ~n868 & ((x2 & x3 & x7 & ~x0 & x1) | (~x1 & ((~x0 & ~x2 & x3 & x7) | (x0 & (x2 ? (~x3 & x7) : (x3 & ~x7))))));
  assign n1254 = (~x2 | n1257) & (~n543 | n1255) & (x2 | n1256);
  assign n1255 = (x0 | ((~x3 | ~x4 | ~x5 | x1 | ~x2) & (~x1 | x2 | x4 | x5))) & (x4 | ((~x0 | x1 | ~x2 | x3 | ~x5) & (~x3 | x5 | ~x1 | x2))) & (x1 | x2 | ~x4 | ((x3 | x5) & (~x0 | (x3 & x5))));
  assign n1256 = (x4 | ((~x5 | x7 | x0 | ~x1) & (x1 | ((~x0 | (x3 ? (~x5 | ~x7) : (x5 | x7))) & (~x5 | ~x7 | x0 | x3))))) & (x0 | ~x1 | ~x4 | (x3 ? (x5 | ~x7) : (x5 ^ x7)));
  assign n1257 = (~x4 | x5 | ~x7 | ~x0 | x1 | ~x3) & (x0 | ((~x5 | ((x1 | x3 | ~x4 | x7) & (~x1 | x4 | (~x3 ^ x7)))) & (x1 | x3 | ~x4 | x5 | ~x7)));
  assign z064 = n1259 | ~n1265 | (n664 & ~n1270) | (~x2 & ~n1269);
  assign n1259 = ~x1 & (n1261 | ~n1262 | (x0 & ~n1260));
  assign n1260 = (~x2 | ((x3 | x4 | x5 | ~x6 | ~x7) & (~x3 | ~x4 | ~x5 | x6 | x7))) & (~x3 | ~x5 | ~x6 | ~x7 | (x2 & ~x4));
  assign n1261 = ~n912 & ((~x7 & n616 & x3 & x4) | (~x3 & ~x4 & x7 & n651));
  assign n1262 = n1264 & (~n559 | ~n1263);
  assign n1263 = ~x3 & ~x0 & x2;
  assign n1264 = (x0 | x3 | ~x6 | ~x7 | (x2 ^ x4)) & (~x0 | ~x2 | ~x3 | x4 | x6 | x7);
  assign n1265 = (~x2 | n1268) & (n620 | n1266) & (n627 | n1267);
  assign n1266 = (x2 | ((~x1 | ((x4 | (x0 ? (~x3 ^ x5) : (~x3 | ~x5))) & (x0 | x3 | x5))) & (x0 | x5 | ((x3 | x4) & (x1 | ~x3 | ~x4))) & (x1 | ~x4 | ~x5 | (~x0 & x3)))) & (x3 | ~x4 | x5 | ~x0 | x1) & (~x2 | ((x1 | (x3 ? (x4 | ~x5) : (~x4 | x5))) & (x0 | ~x1 | (x4 ^ x5))));
  assign n1267 = (~x3 | ~x6 | ~x7 | x0 | x1 | ~x2) & (x2 | (x1 ? (~x6 | ~x7) : (x6 | x7)) | (~x0 ^ x3));
  assign n1268 = (x1 | ((~x0 | ~x4 | ~x6 | (~x3 ^ x5)) & (x4 | x6 | ((x3 | ~x5) & (x0 | ~x3 | x5))))) & (x0 | ~x1 | ((~x5 | ~x6 | x3 | x4) & (x5 | x6 | ~x3 | ~x4)));
  assign n1269 = x4 ? ((x0 | x1 | ~x3 | ~x5 | ~x6) & (x6 | ((x0 | x1 | x3 | x5) & (~x0 | (x1 ? (x3 | ~x5) : (~x3 | x5)))))) : (x5 | (x1 ? (x6 | (~x0 ^ x3)) : (~x3 | ~x6)));
  assign n1270 = x6 ? ((~x7 | (x2 ? (~x3 | (x4 & ~x5)) : (x3 | ~x4))) & (x2 | x3 | x4 | ~x5 | x7)) : (x7 | ((x2 | ~x3 | ~x4 | ~x5) & (x3 | (x4 ? ~x2 : x5))));
  assign z065 = n1272 | ~n1276 | (~n800 & ~n1275);
  assign n1272 = ~x0 & ((x1 & ~n1273) | (n538 & ~n1274));
  assign n1273 = x6 ? ((~x5 | ~x7 | ~x3 | ~x4) & (x3 | x4 | x5 | x7)) : ((x2 | x3 | x4 | ~x5 | x7) & (~x2 | ((~x5 | ~x7 | x3 | ~x4) & (~x3 | x5 | (~x4 ^ ~x7)))));
  assign n1274 = (x3 | x4 | x5 | ~x6 | ~x7) & (~x3 | ((~x5 | ~x6 | ~x7) & (x4 | x5 | x6 | x7)));
  assign n1275 = (x1 | ((x4 | ((~x0 | ((x3 | x6) & (~x2 | ~x3 | ~x6))) & (x3 | ~x6 | x0 | x2))) & (~x3 | x6 | ((x2 | ~x4) & (x0 | (x2 & ~x4)))))) & (x0 | ((x2 | ~x3 | ~x4 | x6) & (~x6 | ((~x2 | x3 | ~x4) & (~x1 | ((x3 | ~x4) & (~x2 | ~x3 | x4))))))) & (~x0 | ~x1 | x2 | x3 | x6);
  assign n1276 = ~n1280 & (~n738 | n1278) & (x2 ? n1277 : n1279);
  assign n1277 = ((x0 ^ ~x1) | ((~x5 | x7 | ~x3 | ~x4) & (x3 | (x4 ? (x5 | x7) : (~x5 | ~x7))))) & (x1 | ((~x3 | ((x0 | x4 | (~x5 ^ x7)) & (x5 | ~x7 | ~x0 | ~x4))) & (x0 | x3 | x4 | x5 | x7)));
  assign n1278 = (x7 | ((~x3 | x4 | x5 | x6) & (~x6 | ((x3 | x4 | x5) & (x2 | (x3 ? (x4 | ~x5) : ~x4)))))) & (~x4 | ~x5 | ~x7 | ((x3 | x6) & (x2 | ~x3 | ~x6)));
  assign n1279 = x0 ? (x1 ? ((~x5 | ~x7 | x3 | ~x4) & (x5 | x7 | ~x3 | x4)) : (x4 | ~x7 | (~x3 ^ x5))) : ((~x4 | ~x5 | ~x7 | x1 | ~x3) & ((~x5 ^ x7) | (x1 ? (~x3 | x4) : (x3 | ~x4))));
  assign n1280 = ~n806 & (x0 ? ~n1281 : (n1282 | (n538 & n1136)));
  assign n1281 = (~x3 | x6 | x1 | ~x2) & (x3 | ~x6 | ~x1 | x2);
  assign n1282 = ~x2 & (x3 ^ ~x6);
  assign z066 = ~n1286 | ~n1292 | (~x3 & (n1285 | (~x1 & ~n1284)));
  assign n1284 = (~x4 | ((~x0 | x2 | x5 | x6 | ~x7) & (~x5 | ((~x0 | (x2 ? (~x6 | ~x7) : (x6 | x7))) & (~x6 | x7 | x0 | ~x2))))) & (x0 | x4 | ~x5 | (x2 ? (x6 ^ x7) : (~x6 | x7)));
  assign n1285 = n664 & ((x7 & (x2 ? (~x5 & (~x4 ^ x6)) : (x5 & (x4 ^ x6)))) | (~x5 & ~x7 & (x2 ? (x4 & ~x6) : (~x4 & x6))));
  assign n1286 = (n620 | n1291) & (~x3 | n1287) & (x2 | n1290);
  assign n1287 = (n976 | ~n1289) & (~n534 | ~n678) & (n846 | n1288);
  assign n1288 = (~x2 | x4 | x7 | ~x0 | x1) & (x0 | ((~x1 | x2 | ~x4 | x7) & (x4 | ~x7 | x1 | ~x2)));
  assign n1289 = ~x0 & (x6 ^ ~x7);
  assign n1290 = x4 ? (~x6 | x7 | ((~x1 | x3) & (x0 | x1 | ~x3))) : (x6 | (x0 ? (x1 ? (x3 | x7) : (~x3 | ~x7)) : (x1 ? (x3 | ~x7) : (~x3 | x7))));
  assign n1291 = (x1 | ((~x0 | ((~x4 | x5 | ~x2 | ~x3) & (x3 | x4 | ~x5))) & (x3 | ~x4 | x5 | x0 | x2))) & (~x3 | x4 | ~x5 | x0 | ~x1 | ~x2);
  assign n1292 = ~n1295 & n1296 & (x0 ? (x1 | n1294) : n1293);
  assign n1293 = ((x4 ^ x6) | ((~x1 | x2 | ~x3 | x5) & (x1 | ~x2 | (x3 ^ x5)))) & (x4 | ~x5 | x6 | ~x1 | ~x2 | x3) & (x1 | x2 | ((~x5 | ~x6 | ~x3 | x4) & (x3 | (x4 ? (~x5 | x6) : (x5 | ~x6)))));
  assign n1294 = (~x6 | ((~x2 | ~x3 | x4 | x5) & (x2 | (x3 ? (~x4 | ~x5) : (x4 | x5))))) & (~x2 | ~x4 | x6 | (x3 ^ x5));
  assign n1295 = ~n1019 & (x1 ? ((~x0 & x2 & ~x7) | (~x3 & x7 & x0 & ~x2)) : ((x0 ^ x7) & (x2 ^ x3)));
  assign n1296 = (n1007 | n1297) & (~n537 | ~n814 | ~n750);
  assign n1297 = (x0 | ~x1 | ~x2 | ~x4) & (~x0 | x2 | (~x1 ^ x4));
  assign z067 = ~n1309 | (x5 ? (n1305 | (~x1 & ~n1304)) : ~n1299);
  assign n1299 = ~n1300 & ~n1302 & ~n1303 & (~n814 | ~n534 | ~n540);
  assign n1300 = x7 & ~n1301;
  assign n1301 = (~x6 | (x0 ? (x1 | (x2 ? (x3 | x4) : (~x3 | ~x4))) : (~x1 | ~x4 | (~x2 ^ ~x3)))) & (x1 | x4 | x6 | (x0 ? (~x2 | ~x3) : (x2 | x3)));
  assign n1302 = ~n599 & ((x0 & ~x2 & ~x3 & x4 & ~x7) | (~x0 & ((~x2 & x3 & x4 & x7) | (x2 & ~x4 & (x3 ^ x7)))));
  assign n1303 = ~n989 & ((x0 & ~x2 & ~x3 & x4 & x7) | (~x0 & x3 & (x2 ? (~x4 & x7) : (x4 & ~x7))));
  assign n1304 = x2 ? ((x3 | ~x4 | x6 | x7) & (~x6 | ~x7 | ~x3 | x4)) : ((~x0 | x7 | (x3 ? (~x4 | ~x6) : (x4 | x6))) & (x0 | x3 | x4 | ~x6 | ~x7));
  assign n1305 = n664 & (x2 ? ~n1306 : (n1308 | (x3 & ~n1307)));
  assign n1306 = (~x6 | x7 | x3 | ~x4) & (x6 | ~x7 | ~x3 | x4);
  assign n1307 = x4 ? (~x6 | ~x7) : (x6 | x7);
  assign n1308 = ~x7 & x6 & ~x3 & ~x4;
  assign n1309 = ~n1310 & ~n1313 & (x0 ? (x1 | n1312) : n1314);
  assign n1310 = ~n1311 & ((x0 & ((x3 & ~x5 & ~x1 & x2) | (x1 & ~x2 & ~x3 & x5))) | (~x1 & ~x2 & ((x3 & x5) | (~x0 & ~x3 & ~x5))));
  assign n1311 = x4 ? (x6 | ~x7) : (~x6 | x7);
  assign n1312 = (x2 | ~x3 | x4 | x5 | ~x7) & (x3 | ((x2 | ~x5 | (~x4 ^ x7)) & (x5 | x7 | (~x2 & x4))));
  assign n1313 = ~n906 & (x1 ? ((~x2 & ~x4 & ~x5) | (~x0 & x4 & (x2 ^ x5))) : (x2 & x5));
  assign n1314 = x1 ? ((~x5 | ((x4 | ~x7 | x2 | ~x3) & (~x2 | (x3 ? (~x4 | ~x7) : (x4 | x7))))) & (x2 | x3 | ~x4 | x5 | x7)) : ((x5 | ((x4 | ~x7 | x2 | ~x3) & (~x2 | (x3 ? (~x4 | ~x7) : x7)))) & (x2 | x3 | ~x5 | x7));
  assign z068 = n1316 | ~n1322 | (x5 & ~n1321) | (~n857 & ~n1320);
  assign n1316 = ~x2 & ((x6 & n1317 & ~n1319) | (~x3 & ~n1318));
  assign n1317 = ~x0 & x3;
  assign n1318 = (~x4 | ((~x7 | (x0 ? (~x5 | (x1 ^ x6)) : (x5 | ~x6))) & (x6 | x7 | x0 | x5))) & (~x0 | ~x1 | x4 | ~x5 | (~x6 ^ x7));
  assign n1319 = (~x4 | ~x5 | ~x7) & (x1 | x4 | x7);
  assign n1320 = (x4 | (x6 ? ((x3 ^ x5) | (x2 ^ x7)) : ((~x2 | x3 | x5 | x7) & (x2 | ~x5 | ~x7)))) & (~x2 | ~x4 | ((x3 | ~x5 | (~x6 ^ x7)) & (~x6 | ~x7 | ~x3 | x5)));
  assign n1321 = x3 ? (~x4 | ((x0 | ~x2 | x6) & (x1 | ((~x2 | x6) & (~x0 | x2 | ~x6))))) : ((~x4 | x6 | x0 | x2) & (x4 | (x0 ^ ~x1) | (~x2 ^ x6)));
  assign n1322 = ~n1324 & ~n1327 & (n1323 | n1326) & (x5 | n1328);
  assign n1323 = x3 ^ ~x6;
  assign n1324 = ~n1325 & x2 & n598;
  assign n1325 = (x3 | x4 | x5 | x6 | x7) & (~x7 | ((~x3 | x4 | ~x5 | ~x6) & (x3 | (x4 ? (~x5 | x6) : (x5 | ~x6)))));
  assign n1326 = (x0 | ((x1 | x2 | x4 | ~x5 | ~x7) & (x5 | x7 | ~x2 | ~x4))) & (x5 | x7 | ((x1 | ~x2 | ~x4) & (~x0 | ~x1 | x2 | x4)));
  assign n1327 = ~n783 & ((~x0 & ((~x2 & x3 & ~x5) | (~x3 & x5 & ~x1 & x2))) | (~x2 & ~x5 & (x3 ? ~x1 : x0)));
  assign n1328 = (x0 | (x2 ? (x3 ? (x4 | ~x6) : (~x4 | x6)) : (x3 | x4 | (x1 ^ ~x6)))) & (x1 | ~x2 | (x3 ? (x4 | ~x6) : (~x4 | x6)));
  assign z069 = ~n1333 | (~x2 & (~n1330 | (x0 ? ~n1331 : ~n1332)));
  assign n1330 = (~x5 | ((x1 | (x3 ? (x4 | ~x7) : (~x4 | x7))) & (x4 | ~x7 | (x3 ? x0 : ~x1)))) & (~x4 | x5 | (x0 ? (x3 | x7) : (~x3 ^ x7)));
  assign n1331 = (x4 | x6 | ~x7 | (x1 ? (~x3 | x5) : x3)) & (x1 | ~x3 | ~x6 | x7 | (~x4 & x5));
  assign n1332 = (x5 | ~x6 | x7 | x1 | x3 | x4) & (~x1 | ((~x3 | x4 | x5 | ~x6 | x7) & (x3 | ((x6 | ~x7 | x4 | x5) & (~x6 | x7 | ~x4 | ~x5)))));
  assign n1333 = (n662 | n1335) & (~x2 | (n1334 & (x1 | n1336)));
  assign n1334 = (x0 & (x1 | (~x4 & x5))) | (x3 & ((x5 & x7) | (~x4 & (x5 | x7)))) | (x7 & ((~x4 & x5) | (~x0 & ~x1 & x4))) | (x4 & ~x5 & ~x7) | (~x3 & ((~x5 & ~x7) | (x4 & (~x5 | ~x7))));
  assign n1335 = x2 ? ((x0 & x1) | (x3 ? (x4 | ~x5) : (~x4 | x5))) : (x3 ? ((x0 & x1) | (x4 ^ x5)) : ((~x0 | ((x4 | x5) & (~x1 | ~x4 | ~x5))) & (x4 | ((~x1 | x5) & (x0 | x1 | ~x5)))));
  assign n1336 = (x0 | x6 | ~x7 | (x3 ? (~x4 ^ x5) : (~x4 | ~x5))) & (~x0 | x3 | x4 | ~x5 | ~x6 | x7);
  assign z070 = ~n1340 | ~n1345 | (~n620 & ~n1339) | (n605 & ~n1338);
  assign n1338 = (x0 | ((~x5 | ~x6 | ~x7 | x2 | ~x4) & (~x2 | ((x4 | ~x6 | ~x7) & (x6 | x7 | ~x4 | ~x5))))) & (~x0 | ~x2 | ~x4 | x5 | x6 | ~x7);
  assign n1339 = ((~x3 ^ x5) | (x2 ? (~x4 | (x0 & x1)) : (x4 | (~x0 & ~x1)))) & (x2 | ((x0 | ((~x3 | x4 | ~x5) & (~x4 | x5 | x1 | x3))) & (~x3 | ~x4 | ~x5 | ~x0 | x1))) & (x0 | ~x2 | x3 | x4 | x5);
  assign n1340 = n1342 & ((x4 & ~x5 & (~x3 | n1344)) | (n1341 & n1344) | (~x4 & x5 & (x3 | n1344)));
  assign n1341 = (x2 | x3 | x6 | ~x0 | ~x1) & (x0 | x1 | ~x3 | (x2 ^ x6));
  assign n1342 = (~n559 | ~n924) & (~n1176 | (~n587 & (~n537 | ~n1343)));
  assign n1343 = x3 & ~x5;
  assign n1344 = (x2 | x6 | x7 | ~x0 | x1) & (~x2 | ~x6 | ~x7 | x0 | ~x1);
  assign n1345 = n1347 & n1349 & (n627 | n1346);
  assign n1346 = x0 ? (x3 | ((~x1 | x2 | ~x6 | ~x7) & (x6 | x7 | x1 | ~x2))) : (~x3 | ((x2 | ~x6 | ~x7) & (x6 | x7 | x1 | ~x2)));
  assign n1347 = x3 ? (~x5 | ((x6 | n1348) & (x4 | n900))) : (x5 | ((~x6 | n1348) & (~x4 | n900)));
  assign n1348 = (~x2 | x4 | ~x0 | x1) & (x2 | ~x4 | x0 | ~x1);
  assign n1349 = (~n947 | n1351) & (n1350 | ~n598 | ~n1136);
  assign n1350 = x2 ? (~x4 | x5) : (x4 | ~x5);
  assign n1351 = (~x1 | ~x5 | x6 | x7) & (x1 | x5 | ~x6 | ~x7);
  assign z071 = x3 ? (~n1357 | ~n1366) : (~n1353 | ~n1367);
  assign n1353 = (x2 | n1356) & (n927 | n1355) & (~x2 | n1354);
  assign n1354 = (x1 | ((x0 | ~x4 | x5 | x6 | x7) & (~x5 | (x0 ? ((~x6 | ~x7) & (~x4 | x6 | x7)) : ((~x6 | x7) & (x4 | x6 | ~x7)))))) & (x0 | x4 | x5 | ((~x6 | ~x7) & (~x1 | x6 | x7)));
  assign n1355 = (~x6 | ((x2 | ~x5 | ~x0 | x1) & (x0 | (x1 ? ~x5 : (x2 | x5))))) & (~x0 | x5 | x6 | (x1 & x2));
  assign n1356 = x6 ? (x0 ? ((~x1 | (x4 ? (x5 | x7) : (~x5 | ~x7))) & (x1 | x4 | x5 | ~x7)) : ((x5 | ~x7 | ~x1 | x4) & (~x5 | x7 | x1 | ~x4))) : ((x0 | (x4 ? (x5 | x7) : (~x5 | ~x7))) & (~x5 | x7 | ~x0 | ~x4));
  assign n1357 = ~n1360 & ~n1363 & n1364 & (x1 | (n1358 & n1359));
  assign n1358 = (x5 | x6 | ~x7 | x0 | x2 | ~x4) & (~x2 | ((~x0 | ~x4 | x5 | (x6 ^ x7)) & (x0 | x4 | ~x5 | x6 | x7)));
  assign n1359 = (~x0 | ~x4 | ~x5 | ~x6 | x7) & (x0 | x4 | ~x7 | (~x5 ^ ~x6));
  assign n1360 = ~n912 & ((~x7 & n897 & ~n1361) | (~n927 & ~n1362));
  assign n1361 = x1 ^ ~x4;
  assign n1362 = x0 ? (x1 | x2) : (~x1 | ~x2);
  assign n1363 = ~n630 & ((x2 & ~x4 & x0 & ~x1) | (~x0 & x4 & (~x1 ^ ~x2)));
  assign n1364 = x0 | ~x1 | ((~n1365 | n1154) & (x4 | ~n836));
  assign n1365 = x5 & x6;
  assign n1366 = ((x0 ? (x1 | x2) : (~x1 | ~x2)) | (x4 ? (x5 | x7) : (~x5 | ~x7))) & (x2 | ((~x0 | ~x1 | x4 | x5 | x7) & (x0 | x1 | ~x5 | (x4 ^ x7))));
  assign n1367 = ((~x5 ^ x7) | (x0 ? (x4 | (x1 ^ ~x2)) : (~x1 | ~x4))) & (~x1 | x2 | ((~x5 | ~x7 | ~x0 | ~x4) & (x5 | x7 | x0 | x4))) & (x0 | ~x2 | x5 | ((~x4 | ~x7) & (x1 | x4 | x7)));
  assign z072 = n1369 | n1374 | ~n1375 | (~x5 & ~n1373);
  assign n1369 = ~x1 & (n1371 | n1372 | (~x0 & ~n1370));
  assign n1370 = x2 ? (~x5 | ((~x6 | ~x7 | ~x3 | ~x4) & (x3 | x4 | x6 | x7))) : (x5 | ((x3 | x4 | x6 | ~x7) & (~x6 | x7 | ~x3 | ~x4)));
  assign n1371 = ~n1019 & ((x0 & ~x2 & ~x3 & ~x7) | (~x0 & x7 & (~x2 ^ ~x3)));
  assign n1372 = n723 & n541 & (x2 ? (x3 & x6) : ~x6);
  assign n1373 = x2 ? ((~x3 | ~x4 | ~x6 | ~x0 | x1) & (x0 | ((x4 | x6 | x1 | x3) & (~x1 | ((~x4 | x6) & (x3 | x4 | ~x6)))))) : (((x3 ? (x4 | x6) : (~x4 | ~x6)) | (~x0 ^ ~x1)) & (~x3 | x4 | ~x6 | x0 | ~x1));
  assign n1374 = ~n1007 & (x2 ? (n738 & ~n592) : (n664 & ~n927));
  assign n1375 = n1376 & ~n1380 & (n662 | n1379);
  assign n1376 = (n620 | n1378) & (~x5 | n1377);
  assign n1377 = (x1 | (x0 ? (x2 ? (x4 | x6) : (~x4 | ~x6)) : (~x2 | ((x4 | ~x6) & (~x3 | ~x4 | x6))))) & (x0 | ~x1 | ~x4 | (x2 ? (~x3 | ~x6) : (x3 | x6)));
  assign n1378 = x1 ? ((x3 | ~x4 | ~x5 | ~x0 | x2) & (x0 | ((~x4 | x5 | x2 | x3) & (~x2 | x4 | ~x5)))) : ((~x0 | x4 | x5 | (~x2 ^ x3)) & (~x4 | ((~x0 | ~x2 | ~x3 | ~x5) & (x0 | (x2 ? x5 : (x3 | ~x5))))));
  assign n1379 = x0 ? ((x1 | ~x4 | x5 | (x2 & x3)) & (~x1 | x2 | x3 | x4 | ~x5)) : ((x4 | ((~x1 | x2 | x3 | x5) & (x1 | (x2 ? (~x3 | x5) : ~x5)))) & (~x1 | ~x4 | ~x5 | (~x2 ^ x3)));
  assign n1380 = x1 & ((~x4 & ~n1381) | (x3 & n616 & n1382));
  assign n1381 = (~x0 | x2 | x3 | x5 | x6 | ~x7) & (x0 | x7 | ((~x2 | x5 | (x3 ^ x6)) & (x2 | ~x3 | ~x5 | ~x6)));
  assign n1382 = x4 & (x5 ? (~x6 & ~x7) : (x6 & x7));
  assign z073 = ~n1388 | (~x0 & (~n1385 | (x5 & ~n1384)));
  assign n1384 = (x4 | ~x6 | ~x7 | ~x1 | x2 | ~x3) & (~x4 | ((x1 | x2 | ~x3 | ~x6 | x7) & ((x2 ? (~x3 | ~x6) : (x3 | x6)) | (x1 ^ ~x7))));
  assign n1385 = (~n1386 | ~n686) & (n1387 | (~n1112 & (x3 | n846)));
  assign n1386 = ~x3 & ~x1 & ~x2;
  assign n1387 = x1 ? (x2 | ~x7) : (~x2 | x7);
  assign n1388 = n1390 & (n912 | n1389) & (x3 ? n1395 : n1394);
  assign n1389 = x1 ? ((x3 | x4 | x7 | ~x0 | x2) & (x0 | (x2 ? (x3 ? ~x7 : (x4 | x7)) : (~x3 | x7)))) : (x0 ? ((~x2 | ~x3 | x7) & (x4 | ~x7 | x2 | x3)) : (~x7 | (x2 ? (x3 | x4) : ~x3)));
  assign n1390 = ~n1391 & ~n1392 & (~n738 | n1393);
  assign n1391 = x1 & ((~x3 & x5 & x7 & x0 & ~x2) | (~x0 & x2 & (x3 ? (~x5 & ~x7) : (x5 & x7))));
  assign n1392 = ~x1 & (x0 ? ((x5 & ~x7 & x2 & ~x3) | (~x2 & x3 & ~x5 & x7)) : (x3 & (x2 ? (x5 ^ x7) : (~x5 & ~x7))));
  assign n1393 = (x3 & x4 & (x6 | ~x7)) | (~x5 & x6) | (x2 & ~x7) | (x5 & ~x6) | (~x2 & x7);
  assign n1394 = (x0 | x1 | x2 | ~x4 | x5 | x7) & ((x1 ^ ~x7) | ((x0 | (x2 ? (~x4 | x5) : (x4 | ~x5))) & (~x4 | x5 | ~x0 | x2)));
  assign n1395 = (~x4 | ~x5 | ~x7 | ~x0 | x1 | ~x2) & (x2 | ((~x0 | x7 | (x1 ? (x4 | x5) : (~x4 | ~x5))) & (~x4 | ~x5 | ~x7 | x0 | ~x1)));
  assign z074 = n1398 | ~n1399 | ~n1406 | (~n620 & ~n1397);
  assign n1397 = x0 ? ((~x1 | x2 | x3 | x4) & (x1 | ((~x4 | ~x5 | ~x2 | ~x3) & (x2 | (~x3 ^ x4))))) : (x1 ? ((x2 | ~x3 | ~x4) & (x4 | x5 | ~x2 | x3)) : ((x4 | x5 | x2 | x3) & (~x2 | (x3 ? (x4 | x5) : ~x4))));
  assign n1398 = x0 & ((x1 & ~x2 & ~x3 & x4 & ~x6) | (~x1 & ((~x4 & x6 & x2 & x3) | (~x2 & (x3 ? (x4 & ~x6) : (~x4 & x6))))));
  assign n1399 = ~n1404 & ~n1405 & (~n1400 | ~n1401) & (~x2 | n1402);
  assign n1400 = x4 & ~x3 & ~x0 & ~x2;
  assign n1401 = x5 & (x1 ? (~x6 & ~x7) : (x6 & x7));
  assign n1402 = (x0 | ((x1 | ~n772) & (~x1 | ~x5 | x6 | n1403))) & (~x0 | x1 | x5 | ~x6 | n1403);
  assign n1403 = x3 ? (~x4 | x7) : (x4 | ~x7);
  assign n1404 = ~x0 & (x1 ? ((x4 & ~x6 & x2 & ~x3) | (~x2 & x3 & ~x4 & x6)) : (x4 & ~x6 & (x2 ^ ~x3)));
  assign n1405 = n1365 & n545 & (x1 ? (x2 ^ ~x3) : (~x2 & x3));
  assign n1406 = (x4 | n1407) & (n662 | n1408);
  assign n1407 = (x3 | x5 | ~x6 | x0 | x1 | ~x2) & (x6 | (x0 ? (x5 | (x1 ? (x2 | ~x3) : (~x2 | x3))) : (x1 | ~x5 | (~x2 ^ ~x3))));
  assign n1408 = (x1 | (x0 ? (~x2 | x3 | (~x4 & ~x5)) : (x2 | ~x3 | (x4 & x5)))) & (x0 | ~x1 | (x4 & x5) | (~x2 ^ ~x3));
  assign z075 = ~n1412 | (~x1 & (x6 ? (x7 & ~n1411) : ~n1410));
  assign n1410 = (~x7 | (x0 ? (~x5 | (x2 ? (x3 | ~x4) : (~x3 | x4))) : (x5 | (x2 ? (~x3 | x4) : (~x3 ^ ~x4))))) & (~x0 | x2 | x3 | ~x4 | x5 | x7);
  assign n1411 = (x0 | x2 | x3 | ~x4 | ~x5) & (~x2 | (~x3 ^ ~x4) | (~x0 ^ x5));
  assign n1412 = ~n1414 & n1418 & ~n1419 & ~n1420 & (x5 | n1413);
  assign n1413 = x2 ? (((~x3 ^ ~x4) | (x0 ? (x1 | x7) : (~x1 | ~x7))) & (~x0 | x1 | x3 | ~x4 | ~x7)) : ((~x0 | x4 | (x1 ? (~x3 ^ x7) : (~x3 | ~x7))) & (x0 | ~x1 | x3 | ~x4 | ~x7));
  assign n1414 = x1 & ((n1416 & ~n1417) | (n1415 & n1231));
  assign n1415 = ~x3 & x0 & ~x2;
  assign n1416 = ~x0 & ~x7;
  assign n1417 = ((x3 ? (x5 | x6) : (~x5 | ~x6)) | (~x2 ^ x4)) & (~x4 | ~x5 | ~x6 | ~x2 | ~x3);
  assign n1418 = ((~x2 ^ x4) | ((~x3 | x7 | ~x0 | x1) & (x0 | (x1 ? (~x3 | ~x7) : (x3 | x7))))) & (x0 | ~x2 | ~x4 | (x1 ? (x3 | x7) : (~x3 ^ x7)));
  assign n1419 = ~x2 & (((~x1 ^ ~x7) & (x0 ? (~x3 & x4) : (x3 & ~x4))) | (~x3 & ~x4 & (x0 ? (~x1 & ~x7) : (x1 & x7))));
  assign n1420 = n1421 & ((x3 & ~x4 & ~x7 & ~x0 & x2) | ((x3 ^ ~x4) & (x0 ? (x2 & x7) : (~x2 & ~x7))));
  assign n1421 = ~x1 & x5;
  assign z076 = ~n1427 | (x1 ? ~n1423 : (x3 ? ~n1425 : ~n1426));
  assign n1423 = x0 ? (~n563 | ~n568) : n1424;
  assign n1424 = x2 ? (x3 ? ((x6 | ~x7 | ~x4 | ~x5) & (x4 | (x5 ? (~x6 | x7) : (x6 | ~x7)))) : ((~x6 | x7 | ~x4 | x5) & (x4 | ~x5 | x6 | ~x7))) : ((~x5 | ((~x6 | x7 | ~x3 | ~x4) & (x3 | x6 | (~x4 ^ ~x7)))) & (~x3 | x5 | (x4 ? (x6 | ~x7) : (~x6 | x7))));
  assign n1425 = ((~x0 ^ ~x2) | ((x4 | ~x5 | x6 | x7) & (~x6 | ~x7 | ~x4 | x5))) & (~x5 | x6 | x7 | ~x0 | x2 | ~x4) & (x0 | ~x2 | x4 | x5 | ~x6 | ~x7);
  assign n1426 = x0 ? (x5 | ((~x2 | x4 | ~x6 | ~x7) & (x2 | (x4 ? (x6 | ~x7) : (~x6 | x7))))) : ((x2 | x4 | x5 | ~x6 | ~x7) & (~x2 | ~x4 | ~x5 | x6 | x7));
  assign n1427 = ~n1433 & ~n1432 & ~n1431 & ~n1428 & ~n1430;
  assign n1428 = ~n1429 & ((~x2 & ~x3 & ~x4 & x0 & x1) | (~x1 & (x0 ? (x2 ? (~x3 & x4) : (x3 & ~x4)) : (x2 ? (x3 ^ ~x4) : (~x3 & x4)))));
  assign n1429 = x5 ? (~x6 | ~x7) : (x6 | x7);
  assign n1430 = n664 & ((x2 & ~x4 & x6 & (x3 ^ x5)) | (x4 & ((~x2 & x5 & (x3 ^ x6)) | (~x5 & ~x6 & x2 & ~x3))));
  assign n1431 = ~x1 & ((x3 & x4 & x5 & ~x0 & ~x2) | (x2 & ((x4 & ~x5 & ~x0 & ~x3) | (x0 & ~x4 & (x3 ^ x5)))));
  assign n1432 = (~x0 ^ x4) & ((x1 & ~x2 & ~x3 & ~x5) | (~x1 & (x2 ? (x3 & x5) : (x3 ^ x5))));
  assign n1433 = ~n783 & ((~x2 & ~x3 & ~x5 & x0 & ~x1) | (~x0 & x1 & x3 & (~x2 ^ x5)));
  assign z077 = ~n1437 | (x7 & (x0 ? ~n1436 : ~n1435));
  assign n1435 = ((x3 ? (~x5 | x6) : (x5 | ~x6)) | (x1 ? (~x2 | ~x4) : (x2 | x4))) & (x1 | ((~x4 | x5 | ~x6 | x2 | ~x3) & (~x2 | ((x3 | ~x4 | ~x5 | x6) & (x5 | ~x6 | ~x3 | x4))))) & (~x1 | ((~x5 | x6 | x3 | x4) & (x2 | ((x3 | ~x5 | x6) & (x5 | ~x6 | ~x3 | x4)))));
  assign n1436 = (x2 | x3 | ~x4 | ~x5 | x6) & (x1 | ((~x2 | ~x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (x5 | ~x6 | x3 | x4) & (x2 | ~x4 | x6 | (x3 & ~x5))));
  assign n1437 = (~x0 | n1440) & (n846 | n1438) & (x0 | n1439);
  assign n1438 = ((~x2 ^ x4) | (x0 ? (x1 | ~x3) : (x3 | ~x7))) & (x1 | (x2 ? (x3 | ~x4) : (~x3 | x4)) | (x0 & ~x7)) & (~x1 | ((x0 | ((~x3 | ~x4 | ~x7) & (x3 | x4) & (~x2 | (x4 ? ~x3 : ~x7)))) & (x2 | x3 | (~x4 & ~x7)))) & (~x3 | ~x4 | ~x7 | x0 | ~x2);
  assign n1439 = x2 ? (x1 ? ((x3 | ~x4 | ~x5 | x6) & (x5 | ~x6 | ~x3 | x4)) : ((x5 | ~x6 | x3 | x4) & (~x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))))) : ((x1 | ~x3 | ~x4 | ~x5 | x6) & ((x4 ? (x5 | ~x6) : (~x5 | x6)) | (x1 ^ x3)));
  assign n1440 = (x4 | ((x1 | ((x3 | ~x5 | x6) & (x5 | ~x6 | x2 | ~x3))) & (~x1 | x2 | x3 | x5 | ~x6))) & (x1 | ~x4 | ((x3 | x5 | ~x6) & (~x5 | x6 | ~x2 | ~x3)));
  assign z078 = ~n1444 | (~x1 & (x2 ? ~n1442 : ~n1443));
  assign n1442 = (x0 | (((~x4 ^ x6) | (x3 ? (~x5 ^ x7) : (~x5 | ~x7))) & (~x4 | ~x6 | (x3 ? (~x5 | ~x7) : (x5 | x7))) & (x3 | x4 | x6 | (~x5 ^ x7)))) & (~x3 | x4 | x5 | x6 | x7) & (~x5 | ~x6 | ~x7 | ~x0 | x3 | ~x4);
  assign n1443 = (x3 | ~x4 | ~x5 | x6 | x7) & (x0 | (x3 ? (x4 ? (x5 ? (~x6 | x7) : (x6 ^ x7)) : (x5 ? (x6 | ~x7) : (~x6 | x7))) : ((x4 | ~x5 | ~x6 | x7) & (~x7 | (x4 ? (~x5 ^ ~x6) : (x5 | ~x6))))));
  assign n1444 = n1453 & ~n1452 & ~n1450 & ~n1448 & ~n1445 & ~n1447;
  assign n1445 = ~n1446 & ((x6 & ((~x0 & x1 & ~x3 & ~x5) | (x0 & ~x1 & (x3 ^ x5)))) | (~x0 & x1 & x3 & x5 & ~x6));
  assign n1446 = x2 ^ ~x4;
  assign n1447 = ~n846 & (x0 ? (~x1 & (x2 ? (x3 & x4) : (~x3 & ~x4))) : (x1 & (x2 ? (~x3 & x4) : (x3 & ~x4))));
  assign n1448 = ~x6 & n738 & (x2 ? (~x3 & ~n868) : (x3 & n1449));
  assign n1449 = ~x4 & x5;
  assign n1450 = ~n1451 & ((~x2 & x3 & x0 & ~x1) | (x1 & ((~x2 & ~x3) | (~x0 & x2 & x3))));
  assign n1451 = (~x4 | x5 | x6 | x7) & (x4 | ~x5 | ~x6 | ~x7);
  assign n1452 = ~n1215 & (x0 ? (~x1 & ((~x3 & ~x4) | (x2 & x3 & x4))) : (x1 & (x2 ? (~x3 & x4) : (x3 & ~x4))));
  assign n1453 = (n620 | n1456) & (~x1 | (n1455 & (x0 | n1454)));
  assign n1454 = (~x2 | x3 | x4 | x5 | x6 | x7) & (x2 | ((x3 | x4 | (x5 ? (x6 | ~x7) : (~x6 | x7))) & (~x5 | ~x6 | ~x7 | ~x3 | ~x4)));
  assign n1455 = (x4 | ~x5 | x6 | ~x0 | x2 | x3) & (x5 | ((~x0 | x2 | (x3 ? (x4 | x6) : (~x4 | ~x6))) & (x0 | ~x2 | ~x3 | ~x4 | ~x6)));
  assign n1456 = x3 ? (((x0 ? (x1 | x2) : (~x1 | ~x2)) | (x4 ^ x5)) & (x0 | ~x1 | x2 | ~x4 | x5) & (~x0 | x1 | ~x2 | x4 | ~x5)) : ((~x0 | x5 | (x1 ? (x2 | x4) : ~x4)) & (~x1 | ~x5 | ((x2 | ~x4) & (x0 | ~x2 | x4))));
  assign z079 = n1458 | n1462 | n1463 | ~n1464 | (~n662 & ~n1461);
  assign n1458 = ~x1 & (x2 ? ~n1459 : ~n1460);
  assign n1459 = (x0 | x3 | x4 | x5 | x6 | ~x7) & (~x0 | ~x3 | ~x4 | ~x5 | ~x6 | x7);
  assign n1460 = (~x0 | x3 | ~x4 | ~x5 | x6) & (x0 | ((x3 | x4 | x5 | ~x7) & (~x3 | ~x4 | ~x5 | ~x6 | x7)));
  assign n1461 = (~x3 & (x5 ? (x0 ? (x2 ? ~x4 : ~x1) : (x1 | (x2 & x4))) : ((~x2 & x4) | (~x0 & ~x1 & ~x4)))) | (x3 & ((~x0 & (x2 ? (x4 & ~x5) : (~x4 & x5))) | (x1 & (x0 | (x4 & ~x5))) | (x0 & x2 & (~x4 ^ x5)))) | (~x4 & ~x5 & x1 & x2) | (x4 & ((x1 & x2 & x5) | (x0 & ~x5 & (x1 | ~x2))));
  assign n1462 = ~n630 & ((~x1 & ((x0 & (x4 ? x3 : x2)) | (x2 & ~x3 & ~x4) | (~x0 & ((~x3 & x4) | (~x2 & x3 & ~x4))))) | (x1 & ~x2 & ~x3 & x4) | (~x0 & ((x2 & x3 & x4) | (x1 & ~x3 & ~x4))));
  assign n1463 = n808 & ((~x0 & ~x3 & x5 & x6) | (x0 & ~x5 & (x3 ? ~x7 : (~x6 & x7))));
  assign n1464 = (n1465 | ((x1 | x2) & ((x1 & x2) | (~x0 ^ x3)))) & (n1466 | (x0 ? x1 : ~x2));
  assign n1465 = (~x6 | x7 | x4 | ~x5) & (x6 | ~x7 | ~x4 | x5);
  assign n1466 = (~x3 | x4 | x5 | x6 | ~x7) & (x3 | ~x4 | ~x5 | ~x6 | x7);
  assign z080 = ~n1470 | ~n1479 | (~x0 & (x7 | ~n1469) & (~x7 | ~n1468));
  assign n1468 = ((~x4 ^ x6) | ((x1 | (x2 ? (~x3 | ~x5) : (~x3 ^ x5))) & (~x1 | x2 | x3 | x5))) & (x1 | (x2 ? ((x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (x5 | x6 | ~x3 | x4)) : ((x5 | x6 | x3 | x4) & (~x5 | ~x6 | ~x3 | ~x4)))) & (~x4 | ~x5 | ~x6 | ~x1 | ~x2 | ~x3);
  assign n1469 = ((x5 ^ x6) | ((~x1 | x2 | x3 | x4) & (x1 | (x2 ? (x3 | ~x4) : (~x3 | x4))))) & (x1 | (((~x2 ^ ~x3) | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (~x2 | x3 | x4 | x5 | ~x6) & (x2 | ~x3 | ~x4 | ~x5 | x6)));
  assign n1470 = n1474 & (n1471 | ~n1472) & (n1473 | (n1215 & n846));
  assign n1471 = x1 ? (~x3 | x6) : (x3 | ~x6);
  assign n1472 = ~x5 & ~x4 & x0 & ~x2;
  assign n1473 = ((~x2 ^ x4) | (x0 ? (x1 | x3) : (~x1 | ~x3))) & (~x2 | ~x3 | ~x4 | ~x0 | x1);
  assign n1474 = (~n750 | ~n1478) & (n1475 | n1477) & (~n559 | ~n1476);
  assign n1475 = x0 ? (x1 | ~x2) : (~x1 | x2);
  assign n1476 = ~x3 & ~x2 & x0 & ~x1;
  assign n1477 = (~x5 | x6 | x3 | ~x4) & (x5 | ~x6 | ~x3 | x4);
  assign n1478 = ~x6 & x5 & x3 & x4;
  assign n1479 = n1481 & (n633 | n1475) & (n620 | n1480);
  assign n1480 = ((x0 ? (x1 | x3) : (~x1 | ~x3)) | (x2 ? (~x4 | x5) : (x4 | ~x5))) & (~x3 | x4 | ~x5 | ~x0 | x1 | ~x2) & ((x4 ^ x5) | ((~x2 | x3 | x0 | ~x1) & (~x0 | x2 | (~x1 ^ x3))));
  assign n1481 = (x2 & (x0 | x3)) | (~x0 & ~x2) | (x1 & x3) | (n850 & n1451) | (~x1 & ~x3);
  assign z081 = n1483 | n1487 | ~n1488 | (~n662 & ~n1486);
  assign n1483 = ~x2 & (x0 ? ~n1484 : ~n1485);
  assign n1484 = (x4 | x5 | ((x6 | ~x7 | x1 | ~x3) & (~x1 | (x3 ? x7 : (x6 | ~x7))))) & (x1 | x3 | ~x4 | ~x5 | (~x6 ^ x7));
  assign n1485 = x1 ? ((~x3 | ~x4 | ~x5 | ~x6 | x7) & (x3 | x5 | (x4 ? (~x6 | x7) : (x6 | ~x7)))) : ((~x3 | x4 | x5 | x6 | ~x7) & (x3 | ~x4 | ~x5 | ~x6 | x7));
  assign n1486 = (x2 | ((x0 | ~x1 | ~x3 | ~x4 | x5) & ((x4 & ~x5) | ((~x1 | x3) & (~x0 | x1 | ~x3))))) & (~x2 | ((x0 | ~x1 | ~x3 | (x4 ^ x5)) & (x1 | ((~x4 | x5) & (x3 | (~x4 & x5)))))) & (x0 | ~x1 | x3 | x4 | ~x5) & (x1 | (x3 ? (x4 | ~x5) : (~x4 | x5)));
  assign n1487 = ~n630 & (x3 ? ((~x2 & ~x4) ? (~x0 & x1) : ~x1) : ((x0 & (x1 ? (~x2 & x4) : ~x4)) | (~x1 & ~x2 & ~x4) | (~x0 & x1 & x2 & x4)));
  assign n1488 = (n1465 | n1490) & (~x2 | (~n1491 & (~n1489 | ~n698)));
  assign n1489 = ~x3 & ~x0 & x1;
  assign n1490 = x1 ? ((x2 | x3) & (x0 | ~x2 | ~x3)) : ((~x2 | x3) & (~x0 | x2 | ~x3));
  assign n1491 = ~x1 & ((x6 & ~x7 & x4 & x5) | (x3 & ~x4 & ~x5 & ~x6 & x7));
  assign z082 = ~n1495 | (~x3 & (x2 ? ~n1494 : ~n1493));
  assign n1493 = (x6 | ((~x4 | x5 | x7) & (x0 | ~x1 | x4 | (~x5 ^ x7)))) & (~x5 | ~x6 | (x4 ? (x7 | (x0 ^ ~x1)) : ~x7));
  assign n1494 = x4 ? ((x6 | ~x7 | x0 | x5) & (~x5 | ((x1 | ~x6 | ~x7) & (x0 | (x6 ^ x7))))) : (x0 ? (x1 | ((x6 | x7) & (x5 | ~x6 | ~x7))) : ((x5 | x6 | x7) & (~x1 | ~x6 | (~x5 ^ x7))));
  assign n1495 = ~n1499 & (x6 ? (n1496 & (x7 | n1498)) : (n1497 & (~x7 | n1498)));
  assign n1496 = x2 ? (x0 ? (x1 | (x3 ? (x4 ^ x5) : (x4 | ~x5))) : ((x4 | x5 | x1 | x3) & (~x4 | ~x5 | ~x1 | ~x3))) : ((x3 | ~x4 | x5) & (~x3 | x4 | ~x5 | x0 | x1));
  assign n1497 = (x1 | ((~x4 | ((~x3 | ~x5 | x0 | x2) & (~x0 | ~x2 | (~x3 ^ x5)))) & (x2 | x4 | ((x3 | ~x5) & (x0 | ~x3 | x5))))) & (~x0 | x2 | x4 | ((x3 | ~x5) & (~x1 | ~x3 | x5)));
  assign n1498 = (x1 | (x2 ? ((x4 | ~x5 | x0 | x3) & (~x0 | (x3 ? (x4 | ~x5) : (~x4 | x5)))) : ((x3 | x4 | x5) & (x0 | ~x4 | (~x3 ^ x5))))) & (~x0 | x2 | x3 | ((x4 | x5) & (~x1 | ~x4 | ~x5)));
  assign n1499 = x3 & ((n664 & ~n1501) | (~x1 & ~n1500));
  assign n1500 = ((~x4 ^ ~x5) | (~x0 ^ x6) | (x2 ^ ~x7)) & ((x4 ? (x5 | x7) : (~x5 | ~x7)) | (x0 ? (x2 | ~x6) : (~x2 | x6))) & (~x2 | ~x4 | x5 | ~x6 | ~x7) & (x2 | x4 | ~x5 | x6 | x7);
  assign n1501 = ((x2 ? (~x4 | x5) : (x4 | ~x5)) | (~x6 ^ ~x7)) & ((x5 ? (x6 | ~x7) : (~x6 | x7)) | (x2 ^ ~x4)) & (x2 | x4 | x5 | x6 | ~x7);
  assign z083 = x2 ? (~n1506 | ~n1511) : (~n1503 | ~n1510);
  assign n1503 = x0 ? n1505 : n1504;
  assign n1504 = ((~x5 ^ x7) | ((~x1 | (x3 ? (~x4 | ~x6) : x6)) & (x4 | ((x3 | x6) & (x1 | ~x3 | ~x6))))) & (~x6 | ((~x1 | ((x4 | x5 | x7) & (~x5 | ~x7 | x3 | ~x4))) & (x3 | ~x4 | x5 | x7) & (x1 | ~x5 | ~x7 | (~x3 ^ ~x4)))) & (~x3 | x6 | (x4 ? (x5 | x7) : (~x5 | ~x7)));
  assign n1505 = x6 ? ((x3 | (x4 ? (x5 | x7) : (~x5 | ~x7))) & (x1 | ((~x3 | x5 | (~x4 ^ ~x7)) & (~x5 | (x7 ? x3 : ~x4))))) : (((~x5 ^ x7) | (x1 ? (x3 | ~x4) : x4)) & (~x1 | x3 | x4 | x5 | x7) & (x1 | ~x3 | ~x4 | ~x5 | ~x7));
  assign n1506 = ~n1507 & ~n1508 & (~n1489 | ~n698) & (x1 | n1509);
  assign n1507 = ~n620 & ((x3 & x4 & x5 & x0 & ~x1) | (~x0 & ((~x1 & ~x3 & ~x4 & ~x5) | (x1 & (x3 ? (~x4 & x5) : (x4 & ~x5))))));
  assign n1508 = ~n1115 & (x0 ? (~x1 & (x4 ? (x6 ^ ~x7) : (x6 & ~x7))) : (x1 ? (x4 ? (~x6 & ~x7) : (x6 & x7)) : (~x6 & (~x4 ^ x7))));
  assign n1509 = ((~x4 ^ ~x7) | ((x5 | x6 | ~x0 | x3) & (~x5 | ~x6 | x0 | ~x3))) & (x0 | ((x5 | ~x6 | x7 | x3 | ~x4) & (~x3 | ((~x6 | ~x7 | x4 | x5) & (x6 | x7 | ~x4 | ~x5))))) & (~x5 | x6 | ~x7 | ~x0 | ~x3 | x4);
  assign n1510 = ((~x1 ^ x4) | ((~x5 | ~x7 | x0 | x3) & (~x0 | ~x3 | x5 | x7))) & (((~x0 | ~x1 | x3 | x4) & (x0 | x1 | ~x3 | ~x4)) | (~x5 ^ x7)) & (~x0 | ~x5 | ~x7 | (x1 ? (x3 | ~x4) : (~x3 | x4))) & (x4 | x5 | x7 | x0 | x1 | ~x3);
  assign n1511 = (x3 | ((~x0 | x1 | x4 | x5 | ~x7) & (x0 | ~x5 | (x1 ? (x4 ^ x7) : (x4 | ~x7))))) & (x0 | ~x1 | ~x3 | (x4 ? (~x5 ^ x7) : (x5 | x7)));
  assign z084 = n1514 | ~n1517 | n1521 | (x5 ? ~n1520 : ~n1513);
  assign n1513 = x4 ? (x1 ? (x2 | ~x6 | (x0 & x3)) : (~x3 | (x0 ? (~x2 ^ ~x6) : (~x2 | x6)))) : ((x0 | ~x2 | (x1 ^ ~x6)) & (~x0 | ~x1 | x2 | ~x3 | x6));
  assign n1514 = ~x3 & (x5 ? ~n1515 : (n897 & ~n1516));
  assign n1515 = ((x2 ^ x6) | ((x4 | ~x7 | x0 | ~x1) & (~x4 | x7 | ~x0 | x1))) & (x1 | x4 | x6 | (x0 ? (~x2 | ~x7) : (x2 | x7)));
  assign n1516 = (x6 | ~x7 | x1 | ~x4) & (~x1 | x7 | (x4 ^ ~x6));
  assign n1517 = (n927 | n1518) & (~x3 | (~n1519 & (~n1176 | ~n686)));
  assign n1518 = (~x0 & ((~x5 & x6) | (~x2 & ~x3))) | (x1 & (~x5 | x6)) | (x0 & (x5 | ~x6) & (x2 | x3)) | (x2 & x3) | (~x5 & x6 & ~x2 & ~x3) | (~x1 & x5 & ~x6);
  assign n1519 = ~x0 & ~n599 & ((x2 & ~n1002) | (n1156 & n1148));
  assign n1520 = (x1 | ((~x3 | ((~x4 | ~x6 | x0 | ~x2) & (~x0 | (x2 ? (x4 | x6) : (~x4 | ~x6))))) & (x0 | x2 | ((~x4 | x6) & (x3 | x4 | ~x6))))) & (x0 | ~x1 | ~x2 | ~x3 | (~x4 ^ x6));
  assign n1521 = ~n592 & ~n1522;
  assign n1522 = x1 ? ((x3 | x5 | x6 | ~x0 | x2) & (~x6 | ((x2 | x3 | ~x5) & (x0 | (~x2 ^ x5))))) : (x2 ? (x0 ? ((~x3 | ~x5 | ~x6) & (x5 | x6)) : (~x5 | x6)) : ((x3 | x5 | ~x6) & (~x5 | x6 | ~x0 | ~x3)));
  assign z085 = n1524 | ~n1528 | ~n1532 | (~n912 & ~n1527);
  assign n1524 = ~x3 & (x7 ? ~n1526 : ~n1525);
  assign n1525 = x2 ? ((~x4 | x5 | ~x6 | x0 | x1) & ((x5 ^ x6) | (x0 ? (x1 | x4) : (~x1 | ~x4)))) : ((x0 | x4 | (x1 ? (x5 | x6) : (~x5 | ~x6))) & (~x4 | x5 | ~x6 | ~x0 | ~x1));
  assign n1526 = (x2 | ((x0 | ~x1 | ~x4 | x5 | x6) & (~x5 | ((~x4 | ~x6 | x0 | ~x1) & (~x0 | x1 | (~x4 ^ x6)))))) & (x1 | ~x2 | ((~x5 | ~x6 | ~x0 | ~x4) & (x5 | x6 | x0 | x4)));
  assign n1527 = x1 ? ((x3 | ~x7 | x0 | ~x2) & (x2 | x7 | (x0 ? (x3 | x4) : (~x3 ^ x4)))) : ((x0 | ~x2 | x3 | x4 | x7) & (~x3 | (x0 ? (x2 ? (~x4 | x7) : (x4 | ~x7)) : (~x4 | (~x2 ^ ~x7)))));
  assign n1528 = n1531 & (x0 | n1529) & (n800 | n1530);
  assign n1529 = (x7 | ((x2 | ((~x1 | ~x3 | ~x4 | x5) & (x1 | ~x5 | (~x3 ^ x4)))) & (~x1 | ~x2 | (x3 ? (~x4 | ~x5) : (x4 | x5))))) & (~x1 | ~x7 | ((x2 | x3 | x4 | ~x5) & (~x4 | x5 | ~x2 | ~x3)));
  assign n1530 = (~x3 | x4 | ~x6 | x0 | ~x1 | ~x2) & (x2 | ((x0 | ~x1 | x3 | x4 | ~x6) & (~x0 | x1 | ~x4 | (x3 ^ x6))));
  assign n1531 = (~x3 | x5 | x7 | x0 | x1 | ~x2) & (~x7 | ((x3 | (x0 ? (x1 ? (x2 | ~x5) : (~x2 | x5)) : (x1 | (x2 ^ x5)))) & (x0 | ~x1 | x2 | ~x3 | ~x5)));
  assign n1532 = (~x0 | n1533) & (~x3 | (n1535 & (x1 | n1534)));
  assign n1533 = (x2 | ~x3 | x4 | x5 | x7) & (x1 | ((~x5 | x7 | (x2 ? (~x3 ^ x4) : (x3 | x4))) & (x2 | x3 | x4 | x5 | ~x7)));
  assign n1534 = (x0 | ~x2 | x4 | ~x5 | x6 | ~x7) & (x7 | ((~x4 | ~x5 | ~x6 | x0 | ~x2) & (~x0 | x2 | (x4 ? (x5 | x6) : (~x5 | ~x6)))));
  assign n1535 = (x1 | ~x7 | (~x5 ^ ~x6) | (x0 ^ x2)) & (x0 | ~x1 | ~x2 | x5 | x6 | x7);
  assign z086 = (~x6 & ~n1550) | (x6 & ~n1549) | (~x3 & ~n1540) | (x3 & ~n1537);
  assign n1537 = (n620 | n1539) & (~n750 | ~n686) & (x1 | n1538);
  assign n1538 = (x0 & (x4 | (~x2 & x5))) | (x4 & ((x5 & x7) | (~x2 & (x5 | x7)))) | (~x6 & x7) | (x6 & ~x7) | (~x0 & x2 & ~x4 & ~x5);
  assign n1539 = (x2 | ((x0 | ~x1 | x4) & (~x4 | ~x5 | ~x0 | x1))) & (x0 | ~x1 | ((x4 | ~x5) & (~x2 | ~x4 | x5)));
  assign n1540 = ~n1542 & n1544 & (~x0 | n1541);
  assign n1541 = (x1 | ~x2 | ~x6 | (x4 ? (~x5 | ~x7) : (x5 | x7))) & (x6 | ((~x1 | x2 | ~x4 | x5 | ~x7) & (x1 | x4 | ~x5 | (x2 ^ x7))));
  assign n1542 = ~n620 & ((~x5 & n598 & x2 & x4) | (~x4 & ((x5 & n598) | (~x2 & (n598 | n1543)))));
  assign n1543 = x0 & x1;
  assign n1544 = (n1545 | n1548) & (n662 | n1547) & (~n686 | ~n1546);
  assign n1545 = x2 ? (x5 | x6) : (~x5 | ~x6);
  assign n1546 = x2 & ~x0 & ~x1;
  assign n1547 = (~x2 | x4 | x0 | ~x1) & (x2 | ~x4 | ~x0 | x1);
  assign n1548 = (~x4 | x7 | x0 | ~x1) & (x4 | ~x7 | ~x0 | x1);
  assign n1549 = (x1 | ~x3 | ((~x0 | ((~x4 | x5) & (x2 | x4 | ~x5))) & (~x4 | (x5 ? (x0 & ~x2) : x2)))) & (x0 | ~x1 | x3 | (x4 ? (~x2 & x5) : x2));
  assign n1550 = x4 ? ((x3 | ((~x0 | (x1 ? (x2 | ~x5) : ~x2)) & (x1 | (x2 ? ~x5 : x0)))) & (x0 | ~x1 | ~x3 | (x2 & ~x5))) : (x5 | ((x0 | x1 | ~x2 | ~x3) & (~x0 | x2 | (x1 ^ x3))));
  assign z087 = n1552 | ~n1554 | n1557 | n1561 | (~x2 & ~n1562);
  assign n1552 = ~x4 & ((n540 & n916 & n694) | (~x0 & ~n1553));
  assign n1553 = (~x7 | (x1 ^ x3) | (x2 ? (x5 | ~x6) : (~x5 | x6))) & (~x2 | ~x3 | x6 | x7 | (~x1 ^ x5));
  assign n1554 = (n620 | n1556) & (~x2 | n1555);
  assign n1555 = (x3 | ((x0 | ~x1 | x4 | x5 | ~x7) & (~x0 | x1 | ~x4 | ~x5 | x7))) & (x0 | x1 | (x4 ? (x5 | ~x7) : ((x5 | x7) & (~x3 | ~x5 | ~x7))));
  assign n1556 = (~x3 | ~x4 | ~x5 | x0 | x1 | ~x2) & (~x0 | x3 | ((x4 | ~x5 | x1 | ~x2) & (~x1 | x2 | ~x4 | x5)));
  assign n1557 = x4 & ((x5 & ~n1559) | (n1558 & ~n1560));
  assign n1558 = ~x0 & ~x5;
  assign n1559 = x0 ? (x1 | ((x2 | ~x3 | x6 | x7) & (~x6 | ~x7 | ~x2 | x3))) : (~x1 | x2 | x3 | (x6 ^ x7));
  assign n1560 = (x1 | x2 | ~x3 | ~x6 | x7) & (~x1 | ~x2 | (x3 ? (x6 | ~x7) : (~x6 | x7)));
  assign n1561 = ~n592 & (x0 ? ((x1 & ~x2 & ~x3 & x5) | (~x1 & ((x3 & ~x5) | (x2 & (x3 | ~x5))))) : ((x1 & (x2 ? x5 : (x3 & ~x5))) | (x2 & ~x3 & x5) | (~x1 & ~x2 & (x3 ^ ~x5))));
  assign n1562 = x0 ? ((x4 | ((x5 | (x1 ? (~x3 ^ x7) : (x3 | x7))) & (~x5 | x7 | x1 | ~x3))) & (x1 | ~x7 | ((~x4 | ~x5) & (x3 | (~x4 & ~x5))))) : (x1 ? (x7 | (x3 ^ (x4 & x5))) : ((x3 | ~x4 | ~x5 | x7) & (x5 | ~x7 | ~x3 | x4)));
  assign z088 = ~n1569 | (x3 ? ~n1566 : (x2 ? ~n1565 : ~n1564));
  assign n1564 = x5 ? ((~x6 | ~x7 | x0 | x4) & (~x0 | ~x4 | ((~x6 | x7) & (x1 | x6 | ~x7)))) : ((x6 | (x0 ? (x1 ? (x4 | ~x7) : (~x4 | x7)) : (x1 ? (~x4 | x7) : (x4 | ~x7)))) & (x0 | x1 | x4 | ~x6 | x7));
  assign n1565 = (x1 | ~x6 | (x0 ? (~x4 | (x5 ^ x7)) : (x4 | (~x5 ^ x7)))) & (x0 | ~x1 | ~x4 | x6 | (~x5 ^ x7));
  assign n1566 = ~n1567 & (~n724 | ((x5 | ~x7 | ~x2 | ~x4) & (x2 | (x4 ? (x5 | x7) : (~x5 | ~x7)))));
  assign n1567 = n658 & ((~x0 & (x4 ? (~x5 & ~n607) : (x5 & ~n1568))) | (x0 & x4 & x5 & ~n607));
  assign n1568 = ~x2 ^ ~x7;
  assign n1569 = ~n1570 & ~n1571 & ~n1573 & ~n1575 & (x1 | n1572);
  assign n1570 = ~x0 & ((x2 & ((x4 & x5 & ~x1 & ~x3) | (x1 & (x3 ? (x4 & x5) : (~x4 & ~x5))))) | (~x1 & ~x2 & ~x5 & (x3 ^ x4)));
  assign n1571 = n664 & ((~x3 & x4 & x6 & (x2 ^ x5)) | (~x2 & ~x5 & ~x6 & (x3 | ~x4)));
  assign n1572 = (~x4 | ~x5 | ~x6 | ~x0 | x2 | ~x3) & (~x2 | ((~x5 | ~x6 | x0 | ~x3) & (x3 | ((~x5 | x6 | x0 | x4) & (~x0 | ((x5 | x6) & (x4 | ~x5 | ~x6)))))));
  assign n1573 = ~n912 & (n1574 | (x1 & (n1415 | (n650 & n616))));
  assign n1574 = x4 & x3 & ~x2 & ~x0 & ~x1;
  assign n1575 = x0 & ~x1 & (x2 ? (x3 & ~x5) : (~x4 & x5));
  assign z089 = n1578 | ~n1583 | (n1123 & ~n1582) | (~n1577 & ~n1581);
  assign n1577 = x0 ^ ~x6;
  assign n1578 = x4 & (x1 ? ~n1580 : ~n1579);
  assign n1579 = (x0 | ~x3 | ~x5 | ~x6 | x7) & (x6 | (x3 ? (x5 | ~x7 | (x0 & ~x2)) : ((x0 | ~x2 | x5 | x7) & (~x0 | (x2 ? (~x5 | x7) : (x5 | ~x7))))));
  assign n1580 = (x3 | ((~x5 | ~x6 | ~x7 | ~x0 | x2) & (x0 | x5 | (x2 ? (~x6 | x7) : (x6 | ~x7))))) & (x5 | ~x6 | ~x7 | x0 | ~x3);
  assign n1581 = (x2 | (x7 ? ((x3 | x4 | x5) & (x1 | (~x3 ^ ~x4))) : ((~x3 | x4 | x5) & (~x4 | ~x5 | ~x1 | x3)))) & (x1 | ~x3 | (x4 ? (x5 ^ x7) : (~x5 | x7)));
  assign n1582 = (~x5 | x6 | ~x7 | x1 | ~x3) & (x3 | x7 | ((~x1 | ~x6 | (x2 ^ x5)) & (~x5 | x6 | (x1 & x2))));
  assign n1583 = ~n1584 & ~n1586 & ~n1588 & n1589 & (n824 | n1587);
  assign n1584 = ~x4 & ~n1585;
  assign n1585 = (x0 | ~x1 | x2 | ~x3 | ~x6 | ~x7) & (x1 | ((x3 | ~x6 | ~x7 | x0 | ~x2) & (~x0 | x2 | x6 | (x3 ^ x7))));
  assign n1586 = ~x3 & ((~x0 & ~x1 & ~x2 & x4 & ~x6) | (~x4 & ((~x0 & x1 & x2 & ~x6) | (x0 & x6 & (~x1 ^ ~x2)))));
  assign n1587 = (x0 | ~x1 | x2 | x3 | ~x4 | ~x6) & (~x0 | x1 | ((~x4 | ~x6 | x2 | x3) & (x4 | x6 | ~x2 | ~x3)));
  assign n1588 = n923 & ((x0 & x1 & ~x2 & ~x5 & x6) | (~x0 & x2 & x5 & (~x1 ^ x6)));
  assign n1589 = ~n1593 & (n1591 | ~n1592) & (~n1590 | ~n750);
  assign n1590 = x6 & x3 & ~x4;
  assign n1591 = (~x3 | x7) & (~x2 | x3 | ~x7);
  assign n1592 = x4 & (x0 ? (~x1 & x6) : (x1 & ~x6));
  assign n1593 = ~x6 & ~x5 & ~x4 & x3 & ~x0 & ~x1;
  assign z090 = ~n1607 | ~n1604 | n1601 | n1600 | n1595 | n1598;
  assign n1595 = ~x5 & ((n605 & ~n1597) | (x3 & ~n1596));
  assign n1596 = (x4 | x6 | ~x7 | ~x0 | ~x1 | x2) & (x1 | (x0 ? (x7 | ((~x4 | x6) & (~x2 | x4 | ~x6))) : (~x7 | ((x4 | ~x6) & (x2 | ~x4 | x6)))));
  assign n1597 = (x0 | x2 | ~x4 | ~x6 | x7) & (~x2 | ((x6 | x7 | x0 | x4) & ((~x0 ^ x7) | (~x4 ^ x6))));
  assign n1598 = n1599 & ((~x0 & x2 & ~x3 & ~x4 & x5) | (~x5 & ((~x0 & ~x2 & ~x3 & ~x4) | (x0 & x4 & (~x2 ^ ~x3)))));
  assign n1599 = ~x1 & x7;
  assign n1600 = ~x1 & ((~x4 & ~x5 & ~x7 & x0 & ~x2) | (~x0 & x5 & ((~x2 & ~x4 & x7) | (x4 & ~x7))));
  assign n1601 = ~n824 & (n1603 | (n1123 & (n539 | n1602)));
  assign n1602 = x3 & ~x1 & x2;
  assign n1603 = x4 & ~x3 & ~x2 & x0 & x1;
  assign n1604 = n1605 & (n927 | ((~x2 | x5 | x0 | ~x1) & (~x0 | x1 | ~x5)));
  assign n1605 = (~x4 | x5 | ~x7 | (~n924 & (x1 | n1606))) & (~x1 | x4 | ~x5 | x7 | n1606);
  assign n1606 = x0 ? (x2 | x3) : (~x2 | ~x3);
  assign n1607 = (n783 | n1608) & (~x5 | ~n664 | n1609);
  assign n1608 = (x5 | ((x0 | x1 | x2 | ~x3 | x7) & (~x0 | ~x7 | (x1 ? (x2 | x3) : (~x2 | ~x3))))) & (x0 | ~x1 | ~x5 | x7 | (~x2 ^ x3));
  assign n1609 = (x2 | x3 | ~x4 | ~x6 | x7) & (~x7 | ((~x3 | ~x4 | x6) & (~x2 | (~x4 ^ x6))));
  assign z091 = ~n1613 | (~x1 & (x0 ? ~n1611 : ~n1612));
  assign n1611 = (~x5 | x6 | ~x7 | ~x2 | x3 | x4) & (x2 | ((x3 | x4 | x5 | ~x6 | ~x7) & (~x3 | x6 | x7 | (~x4 ^ x5))));
  assign n1612 = (x5 | x6 | x7 | x2 | x3 | ~x4) & (~x2 | ~x6 | ((x3 | ~x4 | x5 | x7) & (~x3 | ~x7 | (~x4 ^ x5))));
  assign n1613 = (~n539 | n1616) & (x2 | n1614) & (~x2 | n1615);
  assign n1614 = (~x1 | ((x0 | ((x5 | ~x6) & (x6 | x7 | ~x3 | ~x5))) & (x3 | x5 | (x7 ? x6 : ~x0)))) & (x0 | ~x3 | x5 | x6 | (x1 & ~x7)) & (~x5 | ((~x6 | (x1 & (~x0 | x3 | ~x7))) & (x1 | ((x3 | ~x7) & (~x0 | (x3 & ~x7))))));
  assign n1615 = (~x6 | ((x0 | ~x1 | x5 | (x3 & ~x7)) & (x1 | ~x5 | (~x0 & (x3 | ~x7))))) & (x0 | (x1 ^ x5) | (x6 & (~x3 | x7))) & (x1 | x5 | x6 | (~x3 & x7));
  assign n1616 = (~x3 | ((~x0 | x4 | x5 | (x6 & x7)) & (~x5 | x6 | ~x7 | x0 | ~x4))) & (x0 | x3 | x6 | x7 | (~x4 ^ ~x5));
  assign z092 = ~n1619 | ~n1623 | ~n1626 | (~n662 & ~n1618);
  assign n1618 = (x1 | ((~x0 | (x2 ? (x3 | x4) : (~x3 | ~x4))) & (x3 | ~x5 | x0 | x2))) & (x0 | x2 | ((x3 | ~x4) & (~x1 | (x4 ? x5 : ~x3))));
  assign n1619 = ~n1622 & (~n1620 | ~n1621) & (~n924 | ~n1478);
  assign n1620 = ~x3 & x2 & x0 & ~x1;
  assign n1621 = ~x7 & ~x6 & x4 & ~x5;
  assign n1622 = ~x6 & ((x0 & ~x1 & x2 & x3) | (~x0 & (x1 ? (x2 & ~x3) : (~x2 & x3))));
  assign n1623 = ~n1624 & (x4 | (~n1625 & (~n1343 | ~n540 | ~n750)));
  assign n1624 = x6 & ((x0 & ~x1 & ~x2 & ~x3 & x4) | (~x0 & ((~x1 & x2 & x3 & x4) | (x1 & ~x2 & ~x3 & ~x4))));
  assign n1625 = n537 & n670 & (x0 ? x5 : (~x3 & ~x5));
  assign n1626 = (n620 | n1627) & (x1 | n1628);
  assign n1627 = x0 ? (x2 | ((x3 | x4) & (~x1 | (x3 & (x4 | x5))))) : (~x2 | ((x1 | (x4 ? x3 : ~x5)) & (~x3 | (~x1 & x4))));
  assign n1628 = (x0 | ~x2 | x3 | x4 | x5 | x6) & (~x0 | ((x2 | ~x3 | x4 | x5 | ~x6) & (~x2 | x3 | ~x4 | ~x5 | x6)));
  assign z093 = n1631 | ~n1633 | ~n1634 | (x0 ? ~n1630 : ~n1632);
  assign n1630 = (x1 | ((x2 | x3 | x4 | x5 | x7) & (~x7 | ((~x2 | ~x4 | (~x3 ^ x5)) & (x4 | x5 | x2 | ~x3))))) & (~x1 | x2 | ~x3 | x4 | x5 | x7);
  assign n1631 = ~x1 & (x0 ? (x2 ? (~x4 & (~x3 ^ x7)) : (x4 & (x3 ^ x7))) : ((~x3 & x4 & ~x7) | (x2 & x3 & (~x4 ^ x7))));
  assign n1632 = (x4 | ((x1 | x3 | ((~x5 | x7) & (~x2 | x5 | ~x7))) & (~x1 | ~x2 | ~x3 | ~x5 | x7))) & (~x1 | x2 | ~x3 | ~x4 | (x5 ^ x7));
  assign n1633 = (~x1 | ((x0 | ((~x2 | (x3 ? (~x4 | x7) : ~x7)) & (x4 | ((x3 | ~x7) & (x2 | ~x3 | x7))))) & (x2 | x3 | x7 | (~x0 & ~x4)))) & (x0 | x1 | x2 | ~x3 | ~x7);
  assign n1634 = x2 ? n1635 : ((x7 | n1637) & (~n565 | ~n586));
  assign n1635 = (~n1229 | ~n1163) & (x5 | n1636);
  assign n1636 = (x1 | ~x4 | ((~x0 | x3 | (x6 ^ x7)) & (x6 | x7 | x0 | ~x3))) & (x0 | ~x1 | ~x3 | x4 | (~x6 ^ x7));
  assign n1637 = (x0 | ~x1 | ~x3 | ~x4 | ~x5 | x6) & (x1 | x4 | ((x5 | ~x6 | x0 | x3) & (~x0 | ~x5 | (~x3 ^ ~x6))));
  assign z094 = ~n1643 | (x1 ? ~n1641 : ~n1639);
  assign n1639 = (x6 | n1640) & (~n1020 | (x0 ? (~x3 | ~x7) : (x3 | x7)));
  assign n1640 = (~x4 | x5 | ~x7 | x0 | ~x2 | ~x3) & (x2 | ((~x5 | ((~x0 | (x3 ? (x4 | ~x7) : (~x4 | x7))) & (x0 | x3 | x4 | x7))) & (x0 | x3 | x4 | x5 | ~x7)));
  assign n1641 = x0 ? (~n563 | ~n1621) : n1642;
  assign n1642 = (~x2 | x3 | x4 | ~x5 | ~x6 | x7) & (x2 | ((~x6 | x7 | x4 | x5) & (~x3 | ~x4 | ~x5 | x6 | ~x7)));
  assign n1643 = x2 ? (n1644 & n1647) : (n1645 & n1646);
  assign n1644 = (x1 | (x0 ? (x3 ? (x4 | x5) : (~x4 | ~x5)) : (x3 ? (~x4 | ~x5) : (~x4 ^ x5)))) & (x0 | ~x1 | (x3 ? (~x4 ^ x5) : (x4 | x5)));
  assign n1645 = (~x0 | x1 | x4 | ~x5 | ~x6) & (x0 | (x1 ? ((x4 | x5 | x6) & (~x5 | ~x6 | ~x3 | ~x4)) : (x5 | (x3 ? (~x4 | x6) : (x4 | ~x6)))));
  assign n1646 = x0 ? (x1 ? (x3 | x4) : (~x4 | (~x3 & x5))) : (x1 ? (x3 | ~x4) : (~x3 | x4));
  assign n1647 = (~x4 | x5 | ~x6 | ~x0 | x1 | x3) & (x0 | (~x1 ^ x4) | (x3 ? (x5 | ~x6) : (~x5 | x6)));
  assign z095 = ~n1656 | ~n1653 | n1652 | n1649 | n1651;
  assign n1649 = ~x5 & ((n814 & n543 & n1546) | (~x2 & ~n1650));
  assign n1650 = x1 ? (~x7 | ((x0 | x4 | ~x6) & (~x4 | x6 | ~x0 | x3))) : (x7 | ((x3 | ~x4 | ~x6) & (~x0 | ((~x4 | ~x6) & (x3 | x4 | x6)))));
  assign n1651 = ~x2 & ((x0 & x1 & ~x3 & ~x4 & ~x5) | (~x0 & ((x1 & (x3 ? (~x4 & x5) : (x4 & ~x5))) | (~x4 & ~x5 & ~x1 & x3))));
  assign n1652 = ~n912 & ((~x0 & x1 & x2 & x3 & ~x4) | (x4 & (x0 ? (~x3 & (~x1 ^ ~x2)) : (~x1 & x3))));
  assign n1653 = ~n1654 & (x6 | ~n629 | n1655);
  assign n1654 = x2 & (((~x3 ^ x5) & (x0 ? (~x1 & ~x4) : (x1 & x4))) | (~x0 & ~x1 & ~x4 & (x3 ^ x5)));
  assign n1655 = (~x0 | x1 | ~x3 | ~x4) & (x0 | x3 | (~x1 ^ x4));
  assign n1656 = (x2 | n1657) & (~x5 | (~n1659 & (x1 | n1658)));
  assign n1657 = (~x5 | ((~x6 | ((x0 | ~x1 | ~x3 | ~x4) & (x1 | ((x3 | x4) & (~x0 | (x3 & x4)))))) & (x0 | ~x1 | x3 | x4 | x6))) & (x1 | ~x4 | x5 | x6 | (~x0 & x3));
  assign n1658 = x7 ? ((~x0 | x2 | x3 | ~x4 | x6) & ((x2 ? (~x4 | ~x6) : (x4 | x6)) | (x0 ^ x3))) : ((x0 ? (~x2 | x3) : (x2 | ~x3)) | (~x4 ^ ~x6));
  assign n1659 = n664 & ((~x4 & x6 & (x2 ? (x3 ^ x7) : (~x3 & ~x7))) | (~x2 & x4 & ~x6 & (~x3 ^ x7)));
  assign z096 = n1662 | ~n1666 | (x4 ? (x6 ? ~n1661 : ~n1665) : (x6 ? ~n1665 : ~n1661));
  assign n1661 = x1 ? ((x2 | x3 | x7) & (~x5 | ((x2 | x3) & (x0 | x7 | (x2 & x3))))) : (((x5 ^ x7) | (~x2 & (x0 | ~x3))) & (~x3 | x7 | x0 | ~x2) & (x5 | ~x7 | (~x0 & x2 & x3)));
  assign n1662 = ~x3 & (x2 ? (x5 & ~n1663) : (~n1664 | (~x5 & ~n1663)));
  assign n1663 = (~x0 | x1 | x4 | ~x6 | ~x7) & (~x4 | x6 | x7 | x0 | ~x1);
  assign n1664 = (x0 | ((~x1 | ~x4 | ~x5 | x6 | ~x7) & (x1 | x4 | x5 | ~x6 | x7))) & (~x5 | ~x6 | x7 | ~x0 | ~x1 | x4);
  assign n1665 = (x0 | ~x1 | ((~x2 | (x5 ^ x7)) & (x5 | ~x7 | (x2 & x3)))) & (x1 | ((x2 | ~x5 | x7) & (~x0 | x3 | ((~x5 | x7) & (x2 | (~x5 & x7))))));
  assign n1666 = x5 ? (n607 | n1668) : (n1669 & (~n758 | n1667));
  assign n1667 = (x4 | x6 | x7 | ~x0 | x2) & (x0 | ((~x2 | x4 | ~x6 | ~x7) & (x6 | x7 | x2 | ~x4)));
  assign n1668 = (~x3 | x4 | ~x0 | x1) & (x0 | (x1 ? (~x3 | ~x4) : (x3 | x4)));
  assign n1669 = (~x3 | ~x4 | ~x7 | x0 | x1 | ~x2) & (~x0 | x2 | ((~x4 | ~x7 | ~x1 | x3) & (x4 | x7 | x1 | ~x3)));
  assign z097 = n1673 | ~n1675 | (x5 ? (x7 ? ~n1671 : ~n1672) : (x7 ? ~n1672 : ~n1671));
  assign n1671 = (x3 | ((~x0 | ((x1 | ~x2 | x6) & (~x1 | x2 | x4 | ~x6))) & (~x2 | ((x1 | ~x4 | ~x6) & (x0 | (~x6 & (~x1 | x4))))))) & (~x2 | ~x6 | (x0 ? (x1 | ~x3) : ~x1)) & (x2 | ((x1 | ~x3 | ~x4 | x6) & (x0 | ((~x3 | x6) & (x1 | ~x4 | (~x3 & x6))))));
  assign n1672 = (x2 | ((x3 | ((x0 | ~x6 | (~x1 & x4)) & (x6 | (~x0 & (~x1 | x4))))) & (~x0 | x1 | ~x6 | (~x3 & ~x4)))) & (x0 | ~x2 | ~x3 | x6 | (x1 & ~x4));
  assign n1673 = ~n1674 & (x2 ? n691 : n723);
  assign n1674 = (x0 | ~x1 | x3 | ~x4 | x6) & (x1 | x4 | (x0 ? (~x3 | x6) : (x3 ^ x6)));
  assign n1675 = ~n1676 & ~n1678 & ~n1679 & ~n1681 & (~n698 | ~n754);
  assign n1676 = ~x6 & ~n1677;
  assign n1677 = (x0 | ~x1 | x2 | x3 | ~x4 | x5) & (~x0 | x1 | ~x3 | (x2 ? ~x5 : (x4 | x5)));
  assign n1678 = ~n885 & ((x0 & ~x2 & ~x3 & x5 & x6) | (~x0 & ((x2 & ~x3 & x5 & ~x6) | (~x5 & x6 & ~x2 & x3))));
  assign n1679 = ~x0 & ~n1680 & ((~x2 & ~x5 & x6 & x7) | (~x6 & ~x7 & x2 & x5));
  assign n1680 = x1 ? (~x3 | x4) : (x3 | ~x4);
  assign n1681 = x6 & n538 & ((~x0 & n985) | (n597 & n610));
  assign z098 = n1683 | ~n1686 | ~n1691 | ~n1694 | (~n620 & ~n1685);
  assign n1683 = ~x3 & ((~x5 & ~n1684) | (n534 & n587));
  assign n1684 = (x2 | ((~x0 | ~x4 | (x1 ? (x6 | x7) : (~x6 | ~x7))) & (x0 | x1 | x4 | x6 | ~x7))) & (x0 | ~x2 | ~x6 | ~x7 | (x1 ^ x4));
  assign n1685 = x0 ? (x1 ? (x2 | (x3 ? (x4 | x5) : ~x4)) : (x3 | (x4 & x5))) : ((x1 | ((x2 | (x3 ? x4 : (~x4 | ~x5))) & (~x3 | (x4 ? ~x2 : ~x5)))) & (x2 | ~x3 | (x4 ? ~x1 : ~x5)));
  assign n1686 = ~n1689 & (~x2 | ~n664 | n1687) & (x2 | n1577 | n1688);
  assign n1687 = x3 ? (~x4 | x6) : (x4 | ~x6);
  assign n1688 = x1 ? (x3 | x4) : (~x3 | ~x4);
  assign n1689 = x5 & n904 & (x0 ? (x2 & n540) : (~x2 & n1690));
  assign n1690 = x7 & ~x4 & x6;
  assign n1691 = x3 ? (x4 | (x5 ? n1693 : n1692)) : (~x4 | (x5 ? n1692 : n1693));
  assign n1692 = (x0 | x6 | (x1 ^ ~x2)) & (~x0 | x1 | ~x2 | ~x6);
  assign n1693 = (~x2 | ~x6 | ~x7 | ~x0 | x1) & (x0 | x6 | x7 | (x1 ^ ~x2));
  assign n1694 = x6 ? (~x7 | n1696) : (n1695 & (x7 | n1696));
  assign n1695 = (x3 | ~x4 | x5 | x0 | x1 | x2) & (x4 | ~x5 | ((x2 | ~x3 | ~x0 | x1) & (x0 | (x1 ? (~x2 | ~x3) : (x2 | x3)))));
  assign n1696 = (x1 | ((x0 | ~x2 | x3 | x4 | ~x5) & (~x0 | ~x3 | x5 | (x2 ^ x4)))) & (x0 | ~x1 | ~x2 | (x3 ? (x4 | x5) : (~x4 | ~x5)));
  assign z099 = n1700 | ~n1702 | (x1 ? ~n1698 : (n1706 | ~n1707));
  assign n1698 = x0 ? (~n563 | ~n762) : n1699;
  assign n1699 = (~x5 | ((x6 | ~x7 | x2 | x4) & (~x3 | ((~x6 | x7 | x2 | x4) & (~x2 | x6 | (~x4 ^ ~x7)))))) & (x3 | ~x4 | x5 | (x2 ? (~x6 ^ x7) : (~x6 | ~x7)));
  assign n1700 = ~n906 & (x1 ? (x0 ? (~x2 & n597) : (x2 ? n597 : n1701)) : ((x2 & n1701) | (~x0 & ~x2 & n597)));
  assign n1701 = x4 & x5;
  assign n1702 = (x1 | n1705) & (n592 | n1703) & (n627 | n1704);
  assign n1703 = x1 ? ((x3 | ~x5 | ~x0 | x2) & (x0 | (x2 ? (x3 | ~x5) : x5))) : ((~x2 | ~x3 | x5) & (x3 | ~x5 | x0 | x2));
  assign n1704 = (~x0 | x1 | x2 | ~x3 | ~x7) & (x0 | ~x2 | (x1 ? (~x3 | ~x7) : (x3 | x7)));
  assign n1705 = (x2 | ((x5 | x7 | ~x0 | x4) & (x0 | ~x4 | ~x7 | (~x3 & x5)))) & (~x0 | x4 | x7 | (x3 & (~x2 | ~x5)));
  assign n1706 = n1365 & ((x3 & ~x4 & ~x7 & ~x0 & x2) | (x0 & x4 & (x2 ? (x3 & x7) : (~x3 & ~x7))));
  assign n1707 = (n662 | n1708) & (n927 | n1709);
  assign n1708 = (~x4 | x5 | ~x0 | x3) & (x0 | x2 | ~x3 | x4 | ~x5);
  assign n1709 = (x0 | ~x2 | x3 | x5 | ~x6) & (~x0 | x2 | ~x3 | ~x5 | x6);
  assign z100 = ~n1715 | (~n783 & ~n1721) | (~x1 & ~n1713) | (x1 & ~n1711);
  assign n1711 = x0 ? (~n563 | ~n1166) : n1712;
  assign n1712 = (x3 | x4 | ~x5 | x6 | x7) & (x2 | ~x4 | x5 | ~x6 | (x3 ^ ~x7));
  assign n1713 = (~x2 | ~x3 | n1714) & (x0 | x2 | x3 | x4 | n1226);
  assign n1714 = (x0 | x4 | ~x5 | x6 | ~x7) & (~x4 | ((~x0 | (x5 ? (~x6 | ~x7) : (x6 | x7))) & (~x6 | x7 | x0 | x5)));
  assign n1715 = ~n1718 & ~n1719 & (x3 ? (n1716 | n1720) : n1717);
  assign n1716 = x4 ? (x5 | x6) : (~x5 | ~x6);
  assign n1717 = (~x4 | ((~x1 | ((x5 | ~x6 | x0 | ~x2) & (~x5 | x6 | ~x0 | x2))) & (~x0 | ((x2 | x5 | ~x6) & (x1 | ((x5 | ~x6) & (~x2 | ~x5 | x6))))))) & (x0 | x1 | x4 | (~x5 ^ x6));
  assign n1718 = ~x1 & ((x0 & ~x4 & ((~x3 & ~x5) | (x2 & x3 & x5))) | (~x3 & x4 & x5 & (~x0 | ~x2)));
  assign n1719 = x1 & ~x3 & ((~x2 & ~x4 & ~x5) | (~x0 & (~x4 ^ x5)));
  assign n1720 = x0 & (x1 | x2);
  assign n1721 = (x1 | (x0 ? (~x5 | (x2 ? (x3 | x7) : (~x3 | ~x7))) : (x5 | (x2 ? (x3 | ~x7) : (~x3 | x7))))) & (~x3 | ~x5 | ~x7 | x0 | ~x1 | ~x2);
  assign z101 = ~n1724 | (x1 & (x0 ? (n665 & n559) : ~n1723));
  assign n1723 = (x3 | ((x4 | ~x5 | x6 | ~x7) & (x5 | ((x2 | ~x4 | (x6 ^ x7)) & (~x6 | x7 | ~x2 | x4))))) & (~x5 | x6 | ((~x3 | ~x4 | x7) & (~x2 | (~x4 ^ x7))));
  assign n1724 = n1727 & (x1 | (x2 ? (x6 | n1726) : n1725));
  assign n1725 = (~x5 | ((x4 | ((~x6 | ~x7 | x0 | x3) & (~x0 | (x3 ? (x6 | ~x7) : (~x6 | x7))))) & (~x0 | ~x3 | ~x4 | (x6 ^ x7)))) & (x0 | x5 | (x4 ? ((x6 | x7) & (~x3 | ~x6 | ~x7)) : (x6 | ~x7)));
  assign n1726 = (x0 | ~x3 | ~x4 | ~x5 | x7) & (~x7 | (x0 ? (x3 ? (~x4 | x5) : (x4 | ~x5)) : (x4 | (x3 ^ x5))));
  assign n1727 = n1731 & (x0 ? n1728 : n1729) & (n927 | n1730);
  assign n1728 = (x4 | ~x5 | ((x2 | x3 | x6) & (x1 | ~x3 | (x2 ^ ~x6)))) & (~x1 | x2 | x3 | ~x4 | ~x6);
  assign n1729 = x5 ? ((x3 | x4 | ~x6 | x1 | ~x2) & (x2 | ((~x4 | x6 | x1 | ~x3) & (~x1 | (x3 ? (x4 | ~x6) : (~x4 | x6)))))) : ((x1 | x4 | (x2 ? (~x3 | x6) : ~x6)) & (~x4 | ~x6 | ~x1 | ~x2));
  assign n1730 = x0 ? ((~x1 | x2 | x3 | x5 | x6) & (~x5 | ~x6 | x1 | ~x2)) : (~x6 | (x1 ? (~x3 | (x2 ^ x5)) : (~x2 | x5)));
  assign n1731 = (x1 | (x0 ? (x5 | (x4 ^ x6)) : (~x5 | (x3 ? (x4 | ~x6) : (~x4 | x6))))) & (x0 | ~x1 | x4 | ((x5 | x6) & (x3 | ~x5 | ~x6)));
  assign z102 = ~n1738 | (x4 ? ~n1735 : (x0 ? ~n1733 : ~n1734));
  assign n1733 = (x2 & (x1 | (x3 & ~x6))) | (x1 & (x5 | (~x6 & ~x7))) | (~x2 & (x3 ? x6 : (~x6 & x7))) | (x5 & ~x7) | (~x5 & x7 & (~x1 | x6));
  assign n1734 = (x3 | (x5 ^ x7) | (x1 ? x6 : (x2 | ~x6))) & (~x2 | ((x6 | ~x7 | ~x3 | ~x5) & (~x1 | ((~x3 | ~x5 | ~x7) & (x5 | x6 | x7)))));
  assign n1735 = x0 ? (x1 | n1737) : n1736;
  assign n1736 = (~x2 | (x5 ^ x7) | ((~x3 | x6) & (~x1 | (~x3 & x6)))) & (x5 | ~x6 | x7 | x1 | x2 | x3) & (~x1 | ~x3 | ~x5 | x6 | ~x7);
  assign n1737 = (x2 | ~x3 | (x5 ? ~x7 : (x6 | x7))) & (~x2 | ~x5 | ~x6 | ~x7) & (x5 | x7 | ((x3 | ~x6) & (~x2 | (x3 & ~x6))));
  assign n1738 = (x2 | n1741) & (n800 | n1739) & (n1099 | n1740);
  assign n1739 = (x6 | ((~x0 | ((x1 | ~x2 | ~x3 | ~x4) & (~x1 | x2 | x3))) & (~x1 | x2 | x3 | ~x4) & (x0 | x1 | (x2 & (x3 | x4))))) & (x0 | ~x6 | (x2 ? (x1 & (x3 | x4)) : ((~x3 | ~x4) & (~x1 | (~x3 & ~x4)))));
  assign n1740 = (x1 | ((~x0 | ~x2 | ~x5 | x6) & (x0 | (x2 ? (x5 | x6) : (~x5 | ~x6))))) & (x0 | ~x1 | ~x2 | x5 | ~x6);
  assign n1741 = (~x1 | ((~x5 | ~x6 | ~x0 | x3) & (x0 | x5 | (x3 ? x6 : (x4 | ~x6))))) & (~x0 | x1 | (x3 ? (x5 | ~x6) : (~x5 | x6)));
  assign z103 = ~n1747 | (~x2 & (n1744 | n1746 | (n1743 & n1621)));
  assign n1743 = x3 & ~x0 & x1;
  assign n1744 = ~x3 & ~n1745;
  assign n1745 = (~x5 | ~x6 | ~x7 | x0 | ~x1) & (x6 | ((x7 | ((x0 | ~x1 | x4 | x5) & (~x0 | ~x5 | (x1 ^ ~x4)))) & (x4 | x5 | ~x7 | x0 | x1)));
  assign n1746 = ~n662 & ((x3 & ~x4 & ~x0 & x1) | (x0 & ~x1 & ~x3 & ~n627));
  assign n1747 = ~n1749 & (n620 | n1751) & (x1 ? n1748 : n1752);
  assign n1748 = (~x0 | x2 | x3 | x4 | x5 | x6) & (x0 | (x2 ? (x3 ? (~x4 | ~x6) : (x4 | x6)) : (~x4 | (x3 ? (~x5 | x6) : (x5 | ~x6)))));
  assign n1749 = x2 & ((n565 & n1743) | (~x1 & ~n1750));
  assign n1750 = (x4 & (x3 | (x0 & ~x5 & ~x7))) | (~x6 & x7) | (x6 & ~x7) | (~x4 & (~x3 | (~x0 & x5)));
  assign n1751 = (~x1 | ((x0 | (x2 ? (~x3 ^ x4) : (x3 | x4))) & (x2 | x3 | (x4 ? ~x0 : ~x5)))) & (x2 | ((~x4 | ~x5 | x1 | x3) & (~x3 | ((x1 | x4) & (~x0 | x5 | (x1 & x4))))));
  assign n1752 = x3 ? ((x0 | (x2 ? (~x5 | x6) : (~x4 | ~x6))) & (~x4 | (x2 ? x6 : (~x5 | ~x6)))) : ((x0 | x2 | x6 | (~x4 ^ x5)) & (x4 | ~x6 | (~x2 & (~x0 | x5))));
  assign z104 = ~n1758 | (~x3 & ~n1754) | (x1 & ~n1757);
  assign n1754 = (n620 | n1756) & (~x0 | ~n670 | ~n1163) & (x0 | n1755);
  assign n1755 = (x1 | ~x2 | x4 | ~x5 | x6 | ~x7) & (x2 | ((x1 | ~x4 | x5 | x6 | ~x7) & (~x1 | ~x5 | ~x6 | (~x4 ^ x7))));
  assign n1756 = (~x0 | ((~x4 | x5 | x1 | ~x2) & (~x1 | x2 | x4 | ~x5))) & (x2 | x4 | x5 | x0 | ~x1);
  assign n1757 = (x0 | ~x2 | ~x3 | x4 | x5 | x7) & (x2 | ((x4 | ((~x0 | x5 | (~x3 ^ x7)) & (~x5 | x7 | x0 | x3))) & (x0 | ~x4 | ~x7 | (x3 ^ x5))));
  assign n1758 = n1760 & ~n1761 & (~n1317 | n1762) & (x1 | n1759);
  assign n1759 = x3 ? ((x5 ^ x7) | (x0 ? (x2 | ~x4) : (~x2 | x4))) : (x0 ? ((~x5 | x7 | ~x2 | ~x4) & (x2 | x4 | (~x5 ^ x7))) : ((x5 | ~x7 | ~x2 | x4) & (x2 | ~x4 | ~x5 | x7)));
  assign n1760 = (x7 | ((x0 | (x2 ? (x3 | ~x4) : (~x3 | x4))) & (x3 | ~x4 | ~x0 | x2))) & (x0 | ~x2 | ~x7 | ((~x3 | ~x4) & (~x1 | x3 | x4)));
  assign n1761 = ~x1 & ((~x4 & ~x7 & x0 & x3) | (x7 & (x3 ^ ~x4) & (~x0 ^ x2)));
  assign n1762 = (x2 | ~x4 | x5 | x6 | x7) & (~x1 | ((~x2 | x4 | ~x5 | (x6 ^ x7)) & (x2 | ~x4 | x5 | ~x6 | ~x7)));
  assign z105 = ~n1766 | (n735 & ~n1764) | (~x1 & ~n1765);
  assign n1764 = (~x1 | x2 | x3 | ~x4 | ~x5 | x6) & (x1 | (x2 ? ((x5 | ~x6 | x3 | x4) & (~x3 | (x4 ? (~x5 | ~x6) : (x5 | x6)))) : ((~x5 | x6 | ~x3 | x4) & (x3 | ~x4 | x5 | ~x6))));
  assign n1765 = (x6 | ((~x5 | (x0 ? (~x3 | ~x4) : (x2 ? (~x3 | x4) : (x3 | ~x4)))) & (~x0 | ((x4 | x5 | x2 | ~x3) & (~x2 | (x3 ? ~x4 : (x4 | x5))))))) & (~x0 | ~x4 | ~x6 | (x2 ? x3 : ~x5));
  assign n1766 = n1771 & (x0 | (~n1768 & n1770 & (~x4 | n1767)));
  assign n1767 = ((~x3 ^ x6) | ((x5 | ~x7 | x1 | x2) & (~x5 | x7 | ~x1 | ~x2))) & (x1 | ~x2 | x7 | (x3 ? (x5 | ~x6) : (~x5 | x6))) & (~x5 | x6 | ~x7 | ~x1 | x2 | x3);
  assign n1768 = n690 & (x1 ? (~x7 & ~n1545) : n1769);
  assign n1769 = x7 & (x2 ? (x5 & x6) : (~x5 & ~x6));
  assign n1770 = (x5 | (x2 ? (x3 | ~x4) : (x4 | (~x3 ^ x6)))) & (x2 | ~x4 | ((~x5 | ~x6) & (~x3 | (~x5 & ~x6))));
  assign n1771 = (n1772 | ~n1774) & (~n694 | ~n1773) & (n1716 | n1606);
  assign n1772 = x3 ? (x5 | ~x6) : (~x5 | x6);
  assign n1773 = x6 & ~x5 & ~x3 & x4;
  assign n1774 = (x2 ^ ~x4) & (~x0 ^ ~x1);
  assign z106 = n1776 | ~n1781 | (x1 ? ~n1779 : ~n1780);
  assign n1776 = ~x0 & (x5 ? ~n1777 : ~n1778);
  assign n1777 = x2 ? ((x4 | x6 | x7 | ~x1 | x3) & (~x4 | ((~x6 | x7 | x1 | ~x3) & (~x7 | (x1 ? (~x3 ^ x6) : (x3 | x6)))))) : (x4 | ((x6 | x7 | x1 | ~x3) & (~x6 | (x1 ? (~x3 ^ x7) : (x3 | x7)))));
  assign n1778 = (~x2 | ((~x4 | ~x6 | ~x7 | x1 | ~x3) & (x4 | ((x6 | x7 | x1 | ~x3) & (~x1 | (x3 ? (~x6 | x7) : (x6 | ~x7))))))) & (x1 | x2 | ~x4 | ~x7 | (~x3 ^ x6));
  assign n1779 = (x2 | x3 | ~x4 | ~x5 | ~x6) & (x0 | ((x2 | ((x4 | ~x5 | x6) & (~x3 | ((~x5 | x6) & (~x4 | x5 | ~x6))))) & (x3 | x5 | (x4 ? ~x2 : ~x6))));
  assign n1780 = x0 ? (x4 ? (x2 ? (x5 | (~x3 ^ x6)) : (~x5 | (~x3 & ~x6))) : ((x3 | ~x5 | x6) & (x5 | ~x6 | ~x2 | ~x3))) : (x2 ? ((x5 | x6 | x3 | x4) & (~x3 | ~x5 | (x4 & x6))) : (x3 ? (x5 | ~x6) : (~x5 | x6)));
  assign n1781 = (n824 | n1784) & (n846 | n1783) & (~n738 | n1782);
  assign n1782 = x4 ? ((x2 | x5 | (x3 ? (x6 | x7) : (~x6 | ~x7))) & (x6 | x7 | x3 | ~x5)) : ((x3 | ~x5 | ~x6 | x7) & (~x7 | ((~x5 | x6 | x2 | ~x3) & (~x2 | x5 | (~x3 ^ x6)))));
  assign n1783 = x0 ? (x2 | x4 | (~x1 ^ x3)) : (~x2 | (x1 ? ~x3 : (x3 | ~x4)));
  assign n1784 = (~x1 | x2 | x3 | ~x4 | x6) & (x1 | ~x2 | ~x6 | (x0 ? (~x3 | ~x4) : (x3 | x4)));
  assign z107 = ~n1787 | (~x0 & (x1 ? ~n1786 : (n563 & n698)));
  assign n1786 = ((x6 ^ x7) | ((x4 | ~x5 | x2 | ~x3) & (~x2 | (x3 ? (x4 | x5) : (~x4 | ~x5))))) & (x2 | ~x3 | ~x4 | x5 | x6 | x7) & (~x2 | (x3 ? (~x4 | ((~x6 | x7) & (~x5 | x6 | ~x7))) : (x4 | (~x6 ^ x7))));
  assign n1787 = n1789 & ~n1792 & (x3 | n1791) & (~x2 | n1788);
  assign n1788 = (x4 | ~x5 | x6 | x1 | ~x3) & (x0 | ~x1 | ((x3 | ~x4 | x5 | x6) & (~x5 | ~x6 | ~x3 | x4)));
  assign n1789 = (x2 | n1790) & (n1323 | ((~x1 | x2 | x4 | x5) & (x1 | ~x4 | (~x2 ^ x5))));
  assign n1790 = (~x3 | ~x6 | ((x1 | x4 | x5) & (x0 | ~x1 | ~x4))) & (x1 | x3 | x4 | x6 | (~x0 & ~x5));
  assign n1791 = x4 ? ((x2 | (x1 ? ((x6 | ~x7) & (x5 | ~x6 | x7)) : ((x6 | x7) & (x5 | ~x6 | ~x7)))) & (x1 | ~x2 | ~x5 | (~x6 ^ x7))) : ((~x1 | x2 | ~x5 | ~x6 | x7) & (x1 | ((~x5 | ~x6 | ~x7) & (~x2 | (x6 ^ x7)))));
  assign n1792 = n904 & (x4 ? ((~x6 & x7 & ~x2 & ~x5) | (x2 & ((x5 & ~x6 & ~x7) | (x6 & x7)))) : ((x6 ^ x7) & (x2 ^ x5)));
  assign z108 = n1795 | n1798 | n1800 | (~x2 & ~n1794);
  assign n1794 = (~x3 | ((x4 | x5 | x7) & (~x5 | (x0 & x1) | (~x4 ^ x7)))) & (x3 | (x4 ? (x5 | ~x7) : (~x5 | x7))) & (x4 | x5 | x7 | (~x0 & ~x1));
  assign n1795 = ~x3 & ((~n1116 & ~n1796) | (x1 & ~n1797));
  assign n1796 = (x0 | x1 | x4 | x5 | x7) & (~x5 | (x0 & x1) | (~x4 ^ x7));
  assign n1797 = (x0 | ~x2 | x4 | x5 | x6 | x7) & (~x0 | x2 | ~x5 | ~x6 | (~x4 ^ x7));
  assign n1798 = x2 & ~n1799 & (x4 ? ((x5 & x7) | (~x3 & ~x5 & ~x7)) : ((~x5 & x7) | (x3 & x5 & ~x7)));
  assign n1799 = x0 & x1;
  assign n1800 = ~x5 & n814 & ~n1799 & (x2 ? (x6 ^ ~x7) : (x6 ^ x7));
  assign z109 = ~n1805 | n1802 | n1804;
  assign n1802 = ~x2 & ((n559 & n1229) | (x1 & ~n1803));
  assign n1803 = (x0 | x4 | x5 | x6 | x7) & (~x0 | x3 | ((~x4 | (x6 ? ~x5 : ~x7)) & (~x5 | ~x6 | ~x7) & (x5 | (x4 & x6))));
  assign n1804 = ~x6 & n597 & (x0 ? (~x1 & ~x3) : ((~x3 & x7) | (~x1 & x3 & ~x7)));
  assign n1805 = n1799 | (x3 ? ((~x4 | x5 | ~x6) & (~x5 | ((x6 | x7) & (x4 | (x6 & x7))))) : ((~x6 | (x5 ? (~x4 & ~x7) : x4)) & (~x4 | x6 | (x5 & ~x7))));
  assign z110 = n1813 | (~x5 & (n1808 | n1811 | (~x2 & ~n1807)));
  assign n1807 = (~x0 | ~x1 | ((x4 | x6) & (x3 | ~x4 | ~x6))) & (x6 | ~x7 | ~x3 | x4) & (~x4 | ((x0 | (x6 ? ~x3 : x7)) & (x1 | ~x3 | (~x6 & x7))));
  assign n1808 = ~n1809 & ((~n783 & ~n857) | (n598 & (n641 | n1810)));
  assign n1809 = ~x2 ^ ~x3;
  assign n1810 = x7 & ~x4 & ~x6;
  assign n1811 = n1812 & ((~x1 & ((x4 & x6) | (x0 & ~x4 & ~x6))) | (~x0 & (~x4 ^ (x6 | ~x7))));
  assign n1812 = x2 & ~x3;
  assign n1813 = (~x4 | (~x6 ^ ~x7)) & (x4 | (~x6 ^ x7)) & x5 & (~n1799 | n720);
  assign z111 = n1815 | n1818 | n1819 | ~n1820 | (~x4 & ~n1817);
  assign n1815 = ~x7 & ((~n912 & ~n1816) | (n750 & n1773));
  assign n1816 = (x2 | ((x1 | ~x3) & (x0 | (~x3 & ~x4)))) & (x0 | ((~x2 | x3 | x4) & (x1 | (x3 & x4))));
  assign n1817 = (x5 | x7 | (x0 ? (x1 ? (x2 | ~x3) : ~x2) : (~x1 | (~x2 ^ ~x3)))) & (~x0 | x1 | ~x5 | ~x7 | (~x2 & ~x3));
  assign n1818 = ~x2 & ((~x0 & x5 & x7) | (~x3 & ((x5 & x7) | (x0 & ~x5 & ~x7))));
  assign n1819 = x4 & n738 & ((n723 & n665) | (x2 & ~n824));
  assign n1820 = ~n1821 & (~n698 | ~n685) & (x0 | ~x2 | ~n723);
  assign n1821 = ~x7 & ~x5 & x4 & x3 & ~x0 & x2;
  assign z112 = n1823 | ~n1825 | ~n1826 | (~x7 & n616 & ~n1824);
  assign n1823 = ~x6 & (x0 ? ((x3 & ~x7 & ~x1 & x2) | (x1 & ~x2 & ~x3)) : (x2 & (x1 ? (x3 & ~x7) : (~x3 & x7))));
  assign n1824 = (x1 | ~x3 | x4 | x5 | ~x6) & (~x1 | x3 | ~x4 | (~x5 ^ x6));
  assign n1825 = (~x3 | ((x1 | ((x6 | ~x7) & (x2 | ~x6 | x7))) & (~x6 | x7 | x0 | x2))) & (x3 | x6 | ~x0 | x1) & (x0 | ((~x1 | x6 | ~x7) & (~x6 | x7 | x1 | x3)));
  assign n1826 = x0 ? (x2 | n1828) : (n1827 & (x2 | ~n605 | ~n1231));
  assign n1827 = (~x4 | ((~x1 | x2 | x3 | ~x6 | x7) & (x1 | x6 | (x2 ? (~x3 | x7) : (x3 | ~x7))))) & (~x1 | x3 | x4 | x7 | (x2 ^ x6));
  assign n1828 = (x4 | x5 | x6 | ~x1 | ~x3) & (~x5 | ~x6 | x7 | x1 | x3 | ~x4);
  assign z113 = n1830 | n1832 | ~n1833 | n1837 | (~x7 & ~n1836);
  assign n1830 = ~x0 & ((x7 & ~n1831) | (n1449 & n544 & n1602));
  assign n1831 = (x4 | ~x5 | x6 | x1 | ~x2 | ~x3) & (x3 | ((x1 | x2 | x4 | x5 | ~x6) & (~x1 | ((~x5 | ~x6 | x2 | x4) & (x5 | x6 | ~x2 | ~x4)))));
  assign n1832 = ~x0 & ((~x1 & x2 & x3 & x4 & ~x7) | (~x3 & ((~x2 & x4 & x7) | (x1 & ~x4 & (x2 ^ ~x7)))));
  assign n1833 = (x7 | ((x0 | ~x1 | ~x2 | ~x3) & (~x0 | (x1 ? (x2 | x3) : ~x2)))) & n1834 & (~x7 | ((x1 | x2 | ~x3) & (x0 | ((x2 | ~x3) & (x1 | ~x2 | x3)))));
  assign n1834 = (~n568 | ~n1476) & (x3 | ~n534 | ~n1835);
  assign n1835 = ~x4 & ~x7;
  assign n1836 = (~x0 | x2 | x5 | (x1 ? (~x3 | x4) : (x3 | ~x4))) & (x3 | ~x4 | ~x5 | x0 | ~x1 | ~x2);
  assign n1837 = n1599 & ((n651 & n1838) | (n1123 & ~n1839));
  assign n1838 = x5 & ~x3 & x4;
  assign n1839 = x2 ? (~x3 | x5) : (x3 | ~x5);
  assign z114 = n1842 | ~n1845 | n1847 | (~x1 & (~n1841 | ~n1848));
  assign n1841 = (x3 | ~x4 | x0 | x2) & (~x3 | (x0 ? (~x2 | x4) : (x2 ^ x4)));
  assign n1842 = n1843 & ((n1812 & n1844) | (n665 & n672));
  assign n1843 = ~x5 & ~x0 & x1;
  assign n1844 = x7 & x4 & x6;
  assign n1845 = x0 ? (x1 | x3 | (~x2 & ~n597 & ~n1846)) : (~x1 | (~x2 ^ ~x3));
  assign n1846 = ~x7 & ~x6 & ~x4 & x5;
  assign n1847 = ~x0 & ((x1 & x2 & ~x3 & x4 & x5) | (~x1 & ~x2 & (x3 ? (x4 & ~x5) : (~x4 & x5))));
  assign n1848 = (x0 | x4 | ~x6 | (x2 ? (~x3 | ~x5) : (x3 | x5))) & (~x0 | ~x2 | ~x3 | ~x4 | x5 | x6);
  assign z115 = n1850 | n1852 | ~n1854 | (n539 & ~n1853);
  assign n1850 = ~x2 & ((~x4 & ~n1851) | (n943 & n958));
  assign n1851 = (~x1 | ((~x0 | x3 | ~x5 | ~x6 | x7) & (x0 | x5 | (x3 ? (x6 | ~x7) : (~x6 | x7))))) & (~x0 | x1 | ((~x6 | x7 | ~x3 | x5) & (x3 | ~x5 | x6 | ~x7)));
  assign n1852 = ~x3 & ((~x0 & x5 & (x1 ? (x2 & x4) : ~x4)) | (~x4 & ((~x1 & x2) | (~x2 & ~x5 & x0 & x1))) | (~x1 & x4 & ((~x2 & ~x5) | (x0 & (~x2 | ~x5)))));
  assign n1853 = (~x0 | x3 | x4 | ~x5 | x6) & (x0 | ((x3 | x4 | x5 | x6) & (~x3 | (x4 ? (~x5 | x6) : (x5 | ~x6)))));
  assign n1854 = ~n1856 & (~x4 | ~n1812 | n1857) & (x1 | n1855);
  assign n1855 = (~x6 | (x0 ? ((x2 | x3 | x4 | ~x5) & (~x4 | x5 | ~x2 | ~x3)) : (x4 | (x2 ? (~x3 | ~x5) : (x3 | x5))))) & (x2 | x6 | ((x0 | x3 | ~x4 | ~x5) & (~x0 | ~x3 | x4 | x5)));
  assign n1856 = x3 & ((x4 & x5 & ~x1 & x2) | (~x0 & ((x1 & ~x2 & x4 & ~x5) | ((x2 | x5) & (x1 ^ x4)))));
  assign n1857 = (~x5 | x6 | x7 | ~x0 | x1) & (x0 | x5 | (x1 ? (~x6 | ~x7) : (x6 | x7)));
  assign z116 = x2 ? ~n1864 : (~n1859 | ~n1861 | (~x5 & ~n1860));
  assign n1859 = ((~x1 & x6) | ((x0 | x4 | ~x5) & (~x4 | x5 | ~x0 | x3))) & (x1 | ((~x3 | x6 | ((x4 | ~x5) & (x0 | (x4 & ~x5)))) & (x4 | ~x5 | ~x6 | (~x0 & x3)))) & (x0 | ~x3 | ~x6 | (~x4 ^ ~x5));
  assign n1860 = (~x4 | (x0 ? (x1 | (x3 ? (x6 | ~x7) : (~x6 | x7))) : (~x1 | x3 | (~x6 ^ x7)))) & (x0 | x4 | ((x1 | x3 | ~x6 | x7) & (x6 | ~x7 | ~x1 | ~x3)));
  assign n1861 = ~n1863 & (n1862 | (x0 ? (x1 ? (x3 | ~x5) : (~x3 | x5)) : (x3 | x5)));
  assign n1862 = x4 ? (x6 | x7) : (~x6 | ~x7);
  assign n1863 = n723 & n605 & (x0 ? n642 : n641);
  assign n1864 = ~n1866 & n1868 & (x7 ? (~n923 | n1867) : n1865);
  assign n1865 = (~x4 | ~x5 | ~x6 | x0 | x1 | x3) & (x4 | (((~x3 ^ x5) | (x0 ? (x1 | ~x6) : (~x1 | x6))) & (x0 | x1 | x3 | x5 | ~x6)));
  assign n1866 = ~x1 & ((~x0 & x5 & (x3 ? (~x4 & x6) : (x4 & ~x6))) | ((~x4 ^ x6) & (x0 ? (x3 ^ x5) : (~x3 & ~x5))));
  assign n1867 = (x0 | x5 | (x1 ^ x6)) & (~x5 | x6 | ~x0 | x1);
  assign n1868 = x0 ? (x1 | (x3 ? (~x4 | ~x5) : (x4 | x5))) : ((~x3 | ~x4 | x5) & (~x1 | ((~x4 | ~x5 | x6) & (x3 | (~x4 ^ ~x5)))));
  assign z117 = ~n1870 | n1877 | (~x1 & ~n1874);
  assign n1870 = (~x3 | n1873) & (x3 | n1871) & (n824 | n1872);
  assign n1871 = (x4 | ((x6 | (x0 ? (x5 | (x1 ^ ~x2)) : (~x5 | (x1 & x2)))) & (x0 | ~x6 | (x1 ? (~x2 | ~x5) : (x2 | x5))))) & (~x5 | ((~x4 | x6 | x0 | ~x1) & (~x0 | ((x2 | ~x4 | ~x6) & (x1 | ((~x4 | ~x6) & (x2 | (~x4 & ~x6))))))));
  assign n1872 = (x3 | (x0 ? ((x1 | x2 | x4 | x6) & ((x1 ^ ~x2) | (~x4 ^ x6))) : ((x1 | ~x4 | ~x6) & (x4 | x6 | ~x1 | ~x2)))) & (x0 | ~x3 | (x1 ? (~x4 | ~x6) : ((~x4 | x6) & (~x2 | x4 | ~x6))));
  assign n1873 = (x1 | (x0 ? (x4 ? (x5 | ~x6) : (~x5 | x6)) : (x4 | ((x5 | x6) & (x2 | ~x5 | ~x6))))) & (x0 | ~x1 | x5 | (~x4 ^ x6));
  assign n1874 = (~x0 | n1876) & (n1875 | ((~x2 | ~x4 | x6) & (x0 | (~x4 & (~x2 | ~x6)))));
  assign n1875 = x3 ? (~x5 | x7) : (x5 | ~x7);
  assign n1876 = (x2 | ~x4 | ((~x6 | ~x7 | x3 | x5) & (x6 | x7 | ~x3 | ~x5))) & (~x3 | x4 | ~x6 | (~x5 ^ x7));
  assign n1877 = x1 & ((n1415 & n1166) | (~x0 & ~n1878));
  assign n1878 = (~x3 | x4 | x6 | (~x5 ^ x7)) & (~x6 | ((x3 | ~x7 | (x4 ? x5 : x2)) & (~x5 | x7 | ~x3 | ~x4)));
  assign z118 = n1883 | ~n1885 | (~x2 & (n1881 | (n1880 & n762)));
  assign n1880 = x3 & ~x0 & ~x1;
  assign n1881 = ~x3 & ~n1882;
  assign n1882 = (x1 | ((x0 | ~x4 | x5 | x6 | ~x7) & (~x0 | ~x5 | (x4 ? (~x6 | x7) : (x6 | ~x7))))) & (x0 | ~x1 | ((x5 | (x6 ^ x7)) & (x7 | (x4 ? x6 : (~x5 | ~x6)))));
  assign n1883 = ~n927 & ~n1884;
  assign n1884 = x0 ? ((x2 | x3 | (x1 ? (~x5 | x6) : (x5 | ~x6))) & (x1 | ~x5 | x6 | (~x2 & ~x3))) : ((x1 | ~x5 | ~x6) & (x5 | (~x2 & ~x3) | (x1 ^ x6)));
  assign n1885 = ~n1889 & ~n1890 & (~n1886 | ~n1887) & (n592 | n1888);
  assign n1886 = ~x6 & (x3 ? (~x4 & ~x5) : (x4 & x5));
  assign n1887 = ~x2 & x0 & ~x1;
  assign n1888 = ((~x2 & ~x3) | (x0 ? (x1 | ~x6) : (~x1 | x6))) & (x5 | ~x6 | x1 | ~x2) & (~x0 | x2 | x3 | (x1 ? ~x6 : (x5 | x6)));
  assign n1889 = ~x6 & ((~x0 & ~x1 & x4 & x5) | (x0 & ~x4 & ~x5 & (~x1 ^ ~x2)));
  assign n1890 = ~x0 & x6 & ((x1 & x4 & x5) | (~x1 & ~x2 & ~x4 & ~x5));
  assign z119 = n1892 | ~n1895 | n1896 | n1898 | (n664 & ~n1894);
  assign n1892 = ~x1 & ((~x2 & ~n1893) | (x7 & ~n846 & ~x0 & x2));
  assign n1893 = x6 ? ((~x0 | x3 | x4 | ~x5 | x7) & (x0 | ((~x5 | ~x7) & (~x3 | x4 | x5 | x7)))) : (x0 ? (x3 | ((x5 | x7) & (~x4 | ~x5 | ~x7))) : (x5 | ~x7));
  assign n1894 = (x6 & (~x5 | x7)) | (x7 & (x2 | x3 | x4)) | (x5 & ~x6) | (~x4 & ~x7 & ~x2 & ~x3);
  assign n1895 = (x5 | (((~x2 & ~x3) | (x0 ? (x1 | x7) : (~x1 | ~x7))) & (~x0 | x2 | x3 | (x1 ^ ~x7)))) & (x0 | x1 | ~x5 | x7 | (~x2 & ~x3));
  assign n1896 = n539 & (x0 ? (x3 & n1897) : (~x3 & ~n1002));
  assign n1897 = ~x7 & ~x4 & ~x5;
  assign n1898 = ~n912 & ((~x2 & ~x3 & (x0 ? (x1 & x7) : (~x1 & ~x7))) | (x0 & ~x1 & x7 & (x2 | x3)));
  assign z120 = ~n1904 | (~x2 & (n1900 | (~x0 & ~n1903)));
  assign n1900 = x0 & ((n1902 & n770) | (n1901 & n769));
  assign n1901 = x7 & x5 & x6;
  assign n1902 = ~x7 & ~x5 & ~x6;
  assign n1903 = (x3 | ((x1 | ~x6) & (~x5 | x6 | x7 | ~x1 | x4))) & (x1 | x4 | ~x6 | (x5 & ~x7));
  assign n1904 = x6 ? (x7 ? n1905 : n1906) : (x7 ? n1906 : n1905);
  assign n1905 = (~x0 | (x1 ? (x2 | x3) : ~x3)) & (~x1 | x2 | x3 | x4 | x5) & (x1 | (~x2 & (~x3 | ~x4)));
  assign n1906 = x0 ? (x1 | x2 | x3 | (x4 & x5)) : (~x1 | (~x2 & ~x3 & ~x4));
  assign z121 = n1909 | n1910 | (n1148 & ~n1908) | (~n1115 & n1911);
  assign n1908 = (~x0 | ~x1 | ~x3 | x5 | x6 | ~x7) & (x0 | x1 | ((~x6 | x7 | x3 | x5) & (~x3 | ~x5 | (x6 ^ x7))));
  assign n1909 = x7 & (x1 ? (~x0 | (~x2 & ~x3)) : (x0 | x2 | (x3 & x4)));
  assign n1910 = ~x7 & x4 & ~x3 & ~x2 & ~x0 & ~x1;
  assign n1911 = ~x7 & ~x4 & ~x2 & ~x0 & ~x1;
  assign z122 = ~n1917 | (~x4 & (~n1914 | n1916 | (n1913 & ~n1915)));
  assign n1913 = x7 & ~x0 & ~x6;
  assign n1914 = (x0 | x1 | x2 | x3 | x5 | ~x6) & (~x3 | ((~x0 | ~x1 | x2 | x5 | x6) & (x0 | ~x5 | (x1 ? (~x2 | ~x6) : (x2 | x6)))));
  assign n1915 = (x1 | x2 | x3 | x5) & (~x1 | ~x2 | ~x3 | ~x5);
  assign n1916 = n694 & n544 & n1343;
  assign n1917 = (~x0 | (x1 & (x2 | x3))) & (~x3 | ((x0 | ~x1 | ~x2 | ~x4) & (x1 | x2 | x4 | x5))) & (x1 | x2 | x3 | (~x4 & ~x5));
  assign z123 = n1919 | n1920 | n1921 | ~n1925 | (x6 & ~n1923);
  assign n1919 = ~x0 & ((~x2 & ~x3 & ~x4 & (~x1 ^ ~x5)) | (x3 & ((x4 & x5 & ~x1 & x2) | (~x4 & (x1 ? (x2 ^ x5) : (~x2 & ~x5))))));
  assign n1920 = n1148 & ((x3 & ~x5 & ~x6 & x0 & x1) | (~x0 & (x1 ? (x3 ? (~x5 & x6) : (x5 & ~x6)) : (x3 ? (x5 & ~x6) : (~x5 & x6)))));
  assign n1921 = ~n1922 & ~x6 & n1123;
  assign n1922 = (x1 | x2 | x3 | x5 | ~x7) & (~x1 | ~x3 | (x2 ? (~x5 | x7) : (x5 | ~x7)));
  assign n1923 = x0 ? n1924 : ((~n828 | ~n1602) & (~n1082 | ~n745));
  assign n1924 = (x1 | ~x2 | x3 | ~x4 | ~x5 | ~x7) & (~x1 | x2 | ~x3 | x4 | x5 | x7);
  assign n1925 = x0 ? (x1 ? (x2 | x3) : (~x2 | ~x3)) : ((x1 | x2 | x3 | ~x4) & (~x1 | (x2 ? x3 : (~x3 | ~x4))));
  assign z124 = (n648 & ~n1929) | (~x2 & ~n1930) | n1927 | (x2 & ~n1931);
  assign n1927 = ~x4 & ((n537 & n708 & n534) | (x1 & ~n1928));
  assign n1928 = (x0 | ~x2 | ((~x6 | ~x7 | x3 | x5) & (x6 | x7 | ~x3 | ~x5))) & (x2 | ((~x5 | ~x6 | ~x7 | x0 | x3) & (x5 | ((x6 | x7 | x0 | ~x3) & (~x0 | (x3 ? (~x6 | x7) : (x6 | ~x7)))))));
  assign n1929 = (~x2 | ((~x0 | x3 | ~x5 | ~x6 | x7) & (x0 | x5 | (x3 ? (~x6 | x7) : (x6 | ~x7))))) & (~x0 | x2 | ~x5 | x6 | (~x3 ^ ~x7));
  assign n1930 = (~x0 | ((~x3 | ((~x5 | ~x6 | x1 | ~x4) & (x5 | x6 | ~x1 | x4))) & (~x1 | x3 | (~x5 & ~x6)))) & (x3 | ((~x1 & x5) ? x0 : ~x4)) & (x0 | x1 | x4 | (x5 ? x6 : ~x3));
  assign n1931 = (~x3 & ((x1 & ~x4 & ~x5) | (~x0 & ~x1 & (~x4 | (~x5 & ~x6))))) | (x4 & ((x5 & (x3 | (x0 & x6))) | (x3 & (x1 | x6)))) | (x1 & x3 & x5) | (x0 & (x1 | x3));
  assign z125 = n1934 | ~n1935 | ~n1939 | (n735 & ~n1933);
  assign n1933 = (x1 | ~x2 | x3 | ~x4 | ~x5 | ~x6) & (x2 | ((x1 | ~x3 | ~x4 | ~x5 | x6) & (x4 | ((~x5 | ~x6 | x1 | x3) & (~x1 | x5 | (~x3 ^ ~x6))))));
  assign n1934 = x0 & ((x1 & ~x2 & ~x3 & x4 & x5) | (~x1 & ((~x2 & ~x4 & (~x3 ^ x5)) | (x4 & ((x3 & ~x5) | (x2 & (x3 | ~x5)))))));
  assign n1935 = ~n1938 & (~x2 | ((~n664 | n759) & (n1936 | ~n1937)));
  assign n1936 = x0 ? (x3 | ~x5) : (~x3 | x5);
  assign n1937 = ~x1 & (~x4 ^ ~x6);
  assign n1938 = ~x0 & ((~x4 & ((x3 & ~x5 & (x1 ^ ~x2)) | (~x1 & x2 & (~x3 | x5)))) | (x1 & x4 & ((~x3 & x5) | (~x2 & (~x3 | x5)))));
  assign n1939 = (x2 | n1940) & (x0 | (~n1942 & (x1 | n1941)));
  assign n1940 = ((x3 ? (x4 | x6) : (~x4 | ~x6)) | (x0 ? (~x1 | x5) : (x1 | ~x5))) & (x4 | ~x5 | x6 | ~x0 | x1 | x3) & (x0 | ((x1 | x3 | x4 | x5 | ~x6) & (~x1 | ((~x5 | x6 | x3 | x4) & (x5 | ~x6 | ~x3 | ~x4)))));
  assign n1941 = (x2 | x3 | x4 | x5 | x6 | ~x7) & (~x4 | (x3 ^ x6) | (x2 ? (x5 | x7) : (~x5 | ~x7)));
  assign n1942 = n1943 & (x2 ? (x3 ? (x5 & ~x6) : (~x5 & x6)) : (x3 ? (~x5 & ~x6) : (x5 & x6)));
  assign n1943 = ~x7 & x1 & ~x4;
  assign z126 = ~n1950 | (x4 ? (n1949 | (x7 & ~n1948)) : ~n1945);
  assign n1945 = x2 ? (~n664 | n1947) : n1946;
  assign n1946 = (x3 | ((~x0 | x7 | (x1 ? (x5 | x6) : (~x5 | ~x6))) & (~x7 | ((x0 | (x1 ? (~x5 | ~x6) : (x5 | x6))) & (x5 | ~x6 | ~x0 | x1))))) & (~x1 | ~x3 | ((x0 | x6 | (x5 ^ x7)) & (~x6 | x7 | ~x0 | x5)));
  assign n1947 = (~x3 | ~x5 | x6 | x7) & (x3 | ~x6 | (x5 ^ x7));
  assign n1948 = (x1 | ((~x2 | (x0 ? (x3 ? (~x5 | x6) : (x5 | ~x6)) : (~x5 | (x3 ^ x6)))) & (x0 | x2 | x5 | (x3 ^ x6)))) & (x3 | ~x5 | ~x6 | ~x0 | x2) & (x0 | ~x1 | ~x2 | ~x3 | x5 | x6);
  assign n1949 = n873 & ((x5 & ((x0 & (x2 ? (~x3 & x6) : ~x6)) | (~x2 & ((~x3 & ~x6) | (~x0 & x3 & x6))))) | (~x0 & x2 & ~x5 & (~x3 ^ x6)));
  assign n1950 = ~n1953 & n1955 & (x2 ? n1952 : n1951);
  assign n1951 = (~x3 | ((~x0 | x5 | (x1 & (x4 | x6))) & (x0 | x1 | ~x4 | ~x5 | x6))) & (x0 | ((x1 | x3 | x5 | ~x6) & (~x1 | ~x4 | ~x5 | (x3 & ~x6))));
  assign n1952 = (x0 | ~x1 | x3 | x4 | x5 | x6) & (x1 | ((x0 | x3 | ~x5 | (x4 & ~x6)) & (~x3 | ((~x0 | ~x5 | ~x6) & (x5 | x6 | x0 | x4)))));
  assign n1953 = ~n912 & (n1954 | (n1317 & (x1 ? n710 : n1148)));
  assign n1954 = ~x4 & ~x3 & x2 & x0 & ~x1;
  assign n1955 = (n1716 | n1957) & (n1958 | (~n1956 & (~x2 | n1099)));
  assign n1956 = ~x4 & ~x2 & ~x3;
  assign n1957 = (~x0 | ~x1 | x2 | x3) & (x0 | ~x3 | (x1 ^ ~x2));
  assign n1958 = (x0 | ~x1 | x5) & (~x5 | x6 | ~x0 | x1);
  assign z127 = ~n1962 | (~x5 & (x3 ? ~n1961 : ~n1960));
  assign n1960 = (x6 | x7 | ((x0 | (x1 ? (~x2 | x4) : ~x4)) & (x1 | ~x2 | ~x4) & (~x0 | x2 | x4))) & (x1 | ~x4 | ~x6 | ~x7 | (x0 & x2));
  assign n1961 = (~x6 | ~x7 | (x0 ? (x1 | (~x2 & ~x4)) : (~x1 | x4))) & (x0 | x6 | x7 | ((~x2 | ~x4) & (~x1 | x2 | x4)));
  assign n1962 = ~n1966 & (n620 | n1963) & (x3 ? n1964 : n1965);
  assign n1963 = x0 ? (x3 ? (x4 | x5 | (x1 ^ ~x2)) : ((x2 | ~x4 | ~x5) & (x1 | (x2 & ~x4)))) : ((x1 | ~x3 | ~x4) & (x3 | x4 | ~x1 | ~x2));
  assign n1964 = ((x2 & ~x5) | ((x4 | ~x6 | ~x0 | x1) & (~x4 | x6 | x0 | ~x1))) & (x0 | x1 | x4 | x6);
  assign n1965 = (x4 | (x0 ? (x6 | (x1 ? (x2 | ~x5) : ~x2)) : (~x6 | (x1 & x2)))) & (~x1 | ~x4 | ((x5 | x6 | ~x0 | x2) & (x0 | ~x6)));
  assign n1966 = x5 & ((~n662 & ~n1968) | (n677 & n1967));
  assign n1967 = ~x7 & ~x6 & ~x3 & x4;
  assign n1968 = (~x3 | ~x4 | ~x0 | x1) & (x0 | ((~x1 | ~x3 | x4) & (x3 | ~x4 | x1 | ~x2)));
  assign z128 = n1971 | n1974 | n1975 | ~n1976 | (~x4 & ~n1970);
  assign n1970 = (x2 | (x0 ? (x1 | (x3 ? (x5 | ~x7) : (~x5 | x7))) : (~x1 | (~x3 ^ x7)))) & (x1 | ~x2 | x5 | ~x7 | (~x0 ^ x3));
  assign n1971 = ~x1 & ((n629 & ~n1973) | (~x2 & ~n1972));
  assign n1972 = (~x7 | ((~x5 | x6 | x0 | x4) & (x3 | ((~x0 | x5 | (x4 ^ x6)) & (~x5 | ~x6 | x0 | ~x4))))) & (~x0 | x7 | ((x3 | ~x4 | ~x5 | ~x6) & (x5 | (x3 ? (x4 ^ x6) : (~x4 ^ x6)))));
  assign n1973 = (~x0 | (x4 ? (~x6 ^ x7) : ((x6 | x7) & (~x3 | ~x6 | ~x7)))) & (~x3 | x7 | (~x4 ^ ~x6));
  assign n1974 = ~x0 & ((x4 & ((~x1 & ~x2 & x5 & ~x7) | (x1 & x7 & (~x2 | x5)))) | (x1 & x2 & ~x4 & x5 & ~x7));
  assign n1975 = ~n592 & ((x5 & ((~x1 & x2) | (x0 & (x1 ? (~x2 & ~x3) : x3)))) | (~x0 & ~x1 & ~x5 & (~x2 | ~x3)));
  assign n1976 = (~n750 | ~n1979) & (~n694 | ~n1897) & (~n1977 | n1978);
  assign n1977 = x1 & ~x5;
  assign n1978 = ((~x4 ^ x6) | ((x0 | ~x2 | x7) & (x3 | ~x7 | ~x0 | x2))) & (x0 | ((x2 | x3 | x4 | x6 | x7) & (~x4 | ~x6 | ~x7 | ~x2 | ~x3)));
  assign n1979 = x7 & ~x5 & ~x3 & x4;
  assign z129 = x1 ? ~n1983 : (x3 ? ~n1981 : ~n1982);
  assign n1981 = (~x6 | ((~x0 | (x5 & (~x2 | ~x4 | x7))) & (x0 | x2 | x4 | ~x5 | ~x7) & (x5 | (~x2 & ~x4)))) & (x0 | x2 | x5 | x7) & (x6 | (x5 ? ((~x2 | x7) & (~x0 | (~x2 & x7))) : (~x7 | (x0 & x2))));
  assign n1982 = x5 ? ((x2 | (x0 ? (x4 | x6) : (~x6 | ~x7))) & (~x0 | x6 | (x7 & (~x2 | ~x4)))) : ((~x2 | (x0 & (x4 | ~x7))) & (~x0 | ~x6) & (x0 | (x7 ? x6 : ~x4)));
  assign n1983 = n1985 & (x0 | n1984);
  assign n1984 = (~x5 | ~x6 | ~x7 | x2 | x3 | x4) & (x6 | (x2 ? (~x3 | ~x7 | (~x4 ^ ~x5)) : (x3 | x7 | (~x4 ^ x5))));
  assign n1985 = (x2 | ((x0 | ~x3 | x5) & (x3 | ((x5 | ~x6 | ~x7) & (~x0 | ~x5 | (x6 & x7)))))) & (x0 | ((x6 | x7 | ~x2 | ~x5) & (x5 | (~x6 & (x3 | ~x7)))));
  assign z130 = x2 ? ~n1993 : (~n1988 | (~x6 & ~n1987));
  assign n1987 = x0 ? ((~x1 | ~x3 | x4 | x5 | x7) & (x1 | ~x7 | (~x3 & (~x4 | ~x5)))) : ((x1 | ~x3 | ~x4 | x5 | x7) & (~x1 | x3 | (x4 ? (x5 | x7) : ~x7)));
  assign n1988 = ~n1990 & ~n1991 & n1992 & (~n544 | (~n1229 & ~n1989));
  assign n1989 = ~x5 & ~x4 & ~x3 & ~x0 & x1;
  assign n1990 = ~x0 & ((~x1 & x3 & x4 & x5 & ~x6) | (~x3 & ((~x5 & x6 & ~x1 & ~x4) | (x1 & x5 & (x4 ^ x6)))));
  assign n1991 = ~n662 & ((~x3 & (x0 ? x1 : (~x1 & x4))) | (~x0 & ~x1 & ~x4 & (x3 | x5)));
  assign n1992 = (x0 | ~x1 | ~x3 | x6) & (~x0 | x1 | x3 | ~x6 | (x4 & x5));
  assign n1993 = n1994 & ~n1995 & (~x6 | n1996);
  assign n1994 = x0 ? (x1 | ~x6 | (x4 ? (x3 & ~x7) : ~x3)) : ((~x1 | ~x3 | ~x4 | ~x6) & (x1 | x3 | x6));
  assign n1995 = (~x0 | (~x1 & ~x3)) & (x1 | x3 | (x0 & ~x4)) & (~x6 | ~x7) & (x6 | x7) & (~x1 | ~x3 | ~x4);
  assign n1996 = (~x0 | x1 | ((~x5 | ~x7 | x3 | x4) & (x5 | x7 | ~x3 | ~x4))) & (x4 | ~x5 | ~x7 | x0 | ~x1 | ~x3);
  assign z131 = ~n1999 | (~x6 & ((n1176 & n753) | (x7 & ~n1998)));
  assign n1998 = (x4 | ((x0 | ~x1 | ~x2 | ~x3 | ~x5) & (~x0 | ((x3 | ~x5 | x1 | ~x2) & (~x3 | x5 | ~x1 | x2))))) & (x0 | x2 | ~x4 | x5 | (~x1 ^ x3));
  assign n1999 = ~n2002 & n2004 & ~n2005 & (x0 | (~n2000 & n2001));
  assign n2000 = x1 & ((~x2 & ~x3 & ~x4 & x7) | (x4 & ~x7 & x2 & x3));
  assign n2001 = x1 ? ((x2 | x3 | ~x4 | ~x5 | x7) & (~x2 | ~x3 | x4 | x5 | ~x7)) : (x2 | ~x5 | (x3 ? (~x4 | x7) : (x4 | ~x7)));
  assign n2002 = n2003 & (n1144 | (x3 & n746));
  assign n2003 = x2 & x0 & ~x1;
  assign n2004 = x1 ? ((x3 | ~x7 | ~x0 | x2) & (x0 | (x2 ? (x3 | ~x7) : (~x3 | x7)))) : (x3 ? ((~x0 | (x2 ? (x4 | x7) : ~x7)) & (~x7 | (x2 ? x0 : x4))) : ((x0 | (x2 ? x7 : (~x4 | ~x7))) & (x7 | (x2 ? ~x4 : ~x0))));
  assign n2005 = ~x7 & n1120 & n897 & (x1 ? (~x3 & x4) : (x3 ^ ~x4));
  assign z132 = n2007 | n2012 | ~n2013 | (~x0 & ~n2011);
  assign n2007 = x5 & ((~n2008 & n2010) | (~x1 & ~n2009));
  assign n2008 = x2 ? (~x6 | x7) : (x6 | ~x7);
  assign n2009 = (~x4 | ~x6 | ~x7 | x0 | x2 | x3) & (~x2 | ((x0 | x3 | x4 | x6 | ~x7) & (~x0 | x7 | (x3 ? (~x4 | x6) : (x4 | ~x6)))));
  assign n2010 = ~x4 & x3 & ~x0 & x1;
  assign n2011 = (x4 | ((x1 | x2 | x3 | x5 | ~x6) & (~x5 | ((~x1 | ~x3 | (x2 ^ ~x6)) & (x3 | ~x6 | x1 | ~x2))))) & (x2 | ~x4 | x5 | x6 | (~x1 ^ x3));
  assign n2012 = n541 & ((x3 & ~x5 & ~x6 & x1 & ~x2) | (~x1 & ((x2 & (x3 ? (~x5 & x6) : (x5 & ~x6))) | (~x2 & ~x3 & ~x5 & x6))));
  assign n2013 = ~n2015 & ~n2016 & n2018 & (~n2014 | n2017);
  assign n2014 = ~x5 & ~x2 & ~x4;
  assign n2015 = x2 & (x0 ? (~x1 & (x3 ? (x4 ^ x5) : (~x4 & ~x5))) : ((x4 & x5 & ~x1 & x3) | (x1 & (x3 ? (~x4 & ~x5) : (x4 & x5)))));
  assign n2016 = ~x2 & (x0 ? (~x3 & x4) : (x1 ? (x3 ^ ~x4) : (x3 & ~x4)));
  assign n2017 = (~x0 | ~x1 | ~x3 | ~x6 | x7) & (x0 | x1 | x3 | x6 | ~x7);
  assign n2018 = x1 | ((x3 | ~x4 | x0 | ~x2) & (~x0 | x2 | ~x5 | (~x3 ^ ~x4)));
  assign z133 = n2020 | n2024 | n2026 | ~n2027 | (x6 & ~n2023);
  assign n2020 = ~x4 & (x1 ? ~n2021 : ~n2022);
  assign n2021 = (x0 | ~x2 | ~x3 | (x5 ? (~x6 | x7) : (x6 | ~x7))) & (x2 | ((x0 | ~x3 | ~x5 | x6 | x7) & (x5 | ((x6 | ~x7 | x0 | x3) & (~x0 | ~x6 | (~x3 ^ x7))))));
  assign n2022 = (~x5 | x6 | ~x7 | x0 | x2 | ~x3) & (x3 | ((x0 | x2 | x5 | x6 | ~x7) & (~x2 | ((~x0 | (x5 ? (~x6 | x7) : (x6 | ~x7))) & (x6 | x7 | x0 | ~x5)))));
  assign n2023 = x3 ? (~x5 | ((x1 | x2 | x4) & (x0 | (x1 ^ x4)))) : (x5 | ((x0 | ~x1 | (x2 ^ x4)) & (x1 | ((~x2 | x4) & (~x0 | x2 | ~x4)))));
  assign n2024 = x4 & ((n537 & n1343 & n924) | (~x1 & ~n2025));
  assign n2025 = (x0 | x2 | x3 | (x5 ? (~x6 | x7) : (x6 | ~x7))) & (~x2 | ((x0 | x3 | x5 | ~x6 | ~x7) & (~x0 | ~x3 | ~x5 | x6 | x7)));
  assign n2026 = ~n1115 & ((~x0 & (x1 ? (~x4 & x6) : (x4 & ~x6))) | (~x1 & x4 & x6 & (x0 | x2)) | (~x2 & ~x6 & (x1 ^ x4)));
  assign n2027 = ~n2029 & (x0 ? n2028 : (x6 | n2030));
  assign n2028 = (~x1 | x2 | x3 | ~x5 | ~x6) & (x1 | x6 | (x2 ? (~x3 ^ x5) : (x3 | x5)));
  assign n2029 = ~x0 & ((x1 & x2 & x3 & x5 & ~x6) | (~x1 & ~x2 & ~x3 & ~x5 & x6));
  assign n2030 = (x3 | x4 | x5 | x1 | ~x2) & (~x1 | ~x4 | ((x3 | x5) & (x2 | ~x3 | ~x5)));
  assign z134 = ~n2034 | (~x0 & (x3 ? ~n2033 : ~n2032));
  assign n2032 = (x2 | ((x1 | (x4 ? (x6 | x7) : (~x6 | ~x7))) & (x4 | ((~x5 | ~x6 | ~x7) & (x6 | x7 | ~x1 | x5))))) & (~x1 | ~x2 | (x5 ? (x4 ? (~x6 | x7) : (x6 | ~x7)) : (~x6 | ~x7)));
  assign n2033 = (~x5 | ~x6 | ~x7 | x1 | x2 | x4) & (~x2 | ((~x5 | x6 | ~x7 | x1 | x4) & (~x6 | ((x1 | ((x5 | ~x7) & (~x4 | ~x5 | x7))) & (~x1 | ~x4 | x5 | x7)))));
  assign n2034 = n2036 & ~n2040 & (n620 | n2039) & (~n738 | n2035);
  assign n2035 = (~x4 | x7 | ((~x2 | ((x5 | ~x6) & (~x3 | ~x5 | x6))) & (x3 | x5 | ~x6) & (x2 | ~x5 | (x3 ^ x6)))) & (x2 | ~x3 | ~x7 | ((x5 | ~x6) & (x4 | ~x5 | x6)));
  assign n2036 = (x2 | n2038) & (n846 | n2037) & (~n1546 | ~n921);
  assign n2037 = (x0 | ~x1 | x2 | ~x3 | ~x4 | x7) & (x1 | ((~x0 | x4 | ~x7 | (~x2 ^ ~x3)) & (x3 | ~x4 | x7 | x0 | ~x2)));
  assign n2038 = x4 ? ((x3 | ((~x0 | ~x5 | (x1 ^ ~x6)) & (x5 | x6 | x0 | ~x1))) & (x0 | x1 | ~x3 | x5 | x6)) : (~x6 | ((x0 | ~x3 | x5) & (~x0 | ~x1 | x3 | ~x5)));
  assign n2039 = x0 ? ((x2 | x5 | (x1 ? x4 : (~x3 | ~x4))) & (x1 | x4 | ~x5 | (~x2 & x3))) : ((~x1 | ((x4 | ~x5 | ~x2 | ~x3) & (x2 | (x3 ? (~x4 | x5) : ~x5)))) & (x1 | x2 | x3 | x4 | x5) & (~x4 | ((~x2 | x3 | x5) & (x1 | (~x2 ^ x5)))));
  assign n2040 = ~n1307 & ((x0 & ~x5 & (x2 ? ~x1 : ~x3)) | (~x0 & ((x3 & x5) | (x1 & (x5 | (x2 & x3))))) | (~x1 & x5 & (x2 ^ x3)));
  assign z135 = (x7 & (n2042 | (x5 & ~n2043))) | ~n2045 | (~x5 & ~x7 & ~n2044);
  assign n2042 = ~n912 & ((~x1 & ((x0 & (x2 ? (~x3 & ~x4) : (x3 & x4))) | (x3 & x4 & ~x0 & x2))) | (~x0 & x1 & x2 & (x3 ^ x4)));
  assign n2043 = (~x0 | x1 | x2 | x3 | x4 | ~x6) & (x0 | ((x1 | ~x2 | x3 | x4 | ~x6) & (x2 | ((x3 | x4 | x6) & (~x6 | (x1 ? (~x3 ^ x4) : (~x3 | ~x4)))))));
  assign n2044 = (~x3 | x4 | ~x6 | ~x0 | x1 | x2) & (x0 | (x2 ? (~x6 | (x1 ? (x3 | x4) : (~x3 ^ x4))) : (x1 ? (x3 ? (~x4 | ~x6) : (x4 | x6)) : (x3 ? (x4 | x6) : (~x4 ^ x6)))));
  assign n2045 = n2048 & (x1 | n2046) & (x2 | n2047);
  assign n2046 = (~x5 | ~x6 | ~x7 | ~x0 | ~x2 | ~x3) & (x3 | ((~x2 | ((x6 | ~x7 | x0 | x5) & (x7 | (x0 ? (~x5 ^ ~x6) : (~x5 | x6))))) & (x0 | x2 | ~x6 | (~x5 ^ x7))));
  assign n2047 = x0 ? ((~x1 | ((x3 | ~x5 | ~x7) & (x5 | x7 | ~x3 | x4))) & (~x5 | ~x7 | x3 | ~x4) & (x1 | (x3 ? (x4 ? (x5 | x7) : (~x5 | ~x7)) : (x4 | (~x5 ^ x7))))) : ((~x4 | ~x5 | ~x7 | ~x1 | ~x3) & ((~x5 ^ x7) | (x1 ? (x3 | ~x4) : ~x3)));
  assign n2048 = (n800 | n2051) & (~x2 | n2050) & (~x1 | n2049);
  assign n2049 = (x5 | ~x6 | x7 | ~x0 | x2 | x3) & (x0 | ~x3 | ((x6 | ~x7 | x2 | x5) & (x7 | (x2 ? (~x5 ^ ~x6) : (~x5 | x6)))));
  assign n2050 = (x1 | ((~x7 | (~x0 ^ x5) | (~x3 ^ x4)) & (~x3 | x7 | (x0 ? (x4 | ~x5) : (~x4 | x5))))) & (x0 | ~x1 | ((x5 | ~x7 | ~x3 | ~x4) & (x3 | (x4 ? (x5 | x7) : (~x5 | ~x7)))));
  assign n2051 = (~x0 | x1 | ~x2 | ~x3 | ~x4 | x6) & (x2 | x3 | ((x4 | ~x6 | x0 | ~x1) & (~x0 | x6 | (~x1 ^ x4))));
  assign z136 = ~n2053 | n2061 | (~x2 & ~n2060);
  assign n2053 = n2056 & (x6 ? (x7 ? n2054 : n2055) : (x7 ? n2055 : n2054));
  assign n2054 = (x0 | (x1 ? ((x2 | ~x3 | x4 | x5) & (x3 | ~x4 | (~x2 & ~x5))) : ((~x3 | ~x4 | ~x5) & (x4 | x5 | ~x2 | x3)))) & (x1 | ~x4 | (x2 ? (~x3 | x5) : ((~x3 | ~x5) & (~x0 | x3 | x5))));
  assign n2055 = (~x4 | ((x3 | (x0 ? (x1 ? (x2 | x5) : ~x2) : (x1 | ~x5))) & (x0 | ~x1 | ~x3 | (~x2 & ~x5)))) & (x2 | x4 | ((x1 | ~x3 | x5) & (x3 | ~x5 | ~x0 | ~x1)));
  assign n2056 = x2 ? (n2057 & (x1 | ~x6 | n2059)) : (~x6 | n2058);
  assign n2057 = (~x4 | ~x5 | ~x6 | ~x0 | x1 | ~x3) & (x4 | ((x1 | (~x3 ^ x6) | (~x0 & ~x5)) & (x0 | ~x1 | (x3 ? ~x6 : (~x5 | x6)))));
  assign n2058 = ((x3 ? (~x4 | x5) : (x4 | ~x5)) | (x0 ? (x1 | ~x7) : (~x1 | x7))) & (x1 | x3 | ((x5 | ~x7 | x0 | x4) & (~x5 | x7 | ~x0 | ~x4)));
  assign n2059 = (~x4 | x5 | x7 | x0 | x3) & (~x0 | ~x3 | x4 | ~x5 | ~x7);
  assign n2060 = x3 ? ((x5 | x6 | x1 | ~x4) & (x4 | (x1 ? (x0 ? (x5 | x6) : (~x5 | ~x6)) : (~x5 | x6)))) : (x6 ? ((~x1 | x4 | x5) & (x0 | x1 | (~x4 ^ x5))) : ((~x4 | x5 | x0 | ~x1) & (~x0 | (x4 ? ~x5 : x1))));
  assign n2061 = ~x6 & ((n750 & n1144) | (~x1 & ~n2062));
  assign n2062 = (x4 | ~x5 | x7 | x0 | x2 | x3) & (~x2 | ((~x0 | x7 | (x3 ? (~x4 | ~x5) : (x4 | x5))) & (x0 | ~x3 | x4 | x5 | ~x7)));
  assign z137 = ~n2067 | (x2 & (~n2065 | (~x1 & ~n2064)));
  assign n2064 = (~x5 | x6 | ~x7 | ~x0 | x3 | ~x4) & (x0 | x5 | ((~x3 | x4 | ~x6 | x7) & (x3 | (x4 ? (x6 ^ x7) : (x6 | ~x7)))));
  assign n2065 = x7 ? ((x6 | n2066) & (~x3 | ~x5 | n786)) : ((~x6 | n2066) & (x3 | x5 | n786));
  assign n2066 = (x3 | x4 | x5 | x0 | ~x1) & (~x3 | ~x4 | ~x5 | ~x0 | x1);
  assign n2067 = x2 ? n2071 : (n2070 & (x1 ? n2068 : n2069));
  assign n2068 = (~x0 | x3 | x4 | ~x5 | x6 | x7) & (x5 | ~x6 | ~x7 | x0 | ~x3 | ~x4);
  assign n2069 = (x3 | ~x5 | ((x6 | x7 | x0 | ~x4) & (x4 | (x0 ? (x6 ^ x7) : (~x6 ^ x7))))) & (~x0 | ~x3 | x5 | (x4 ? (x6 ^ x7) : (x6 | ~x7)));
  assign n2070 = x4 ? ((x1 | ~x5 | ~x7) & (x0 | (x5 ^ x7)) & (~x0 | x3 | ((x5 | ~x7) & (~x1 | ~x5 | x7)))) : ((x1 | ((x0 | x5 | ~x7) & (~x3 | ~x5 | x7))) & (x0 | ((~x1 | ~x5 | x7) & (~x3 | x5 | ~x7))) & (~x1 | x3 | x5 | x7) & (~x0 | ((x3 | x5 | x7) & (~x1 | ((x5 | x7) & (x3 | ~x5 | ~x7))))));
  assign n2071 = (x0 & (x1 | (x5 & x7))) | (~x5 & ((~x3 & ~x7) | (~x0 & ~x1 & (~x3 | ~x7)))) | (x4 & ~x7) | (x7 & (~x4 | (x1 & x3 & x5)));
  assign z139 = ~n2074 | (~x3 & (x6 ? (~x7 & ~n577) : ~n2073));
  assign n2073 = (x4 | ((x1 | ((~x0 | (x2 ? (~x5 | ~x7) : (x5 | x7))) & (~x5 | x7 | x0 | ~x2))) & (x0 | ~x1 | x2 | ~x5 | x7))) & (~x4 | x5 | ~x7 | ~x0 | ~x1 | x2);
  assign n2074 = n581 & n584 & (x6 ? (x7 ? n579 : n2075) : (x7 ? n2075 : n579));
  assign n2075 = x1 ? (x3 | (x0 ? (x2 | x4) : (~x4 | (~x2 & x5)))) : (x0 ? ((~x4 | ~x5 | x2 | ~x3) & (x4 | x5 | ~x2 | x3)) : ((~x3 | x4 | (~x2 & x5)) & (~x4 | ~x5 | x2 | x3)));
  assign z140 = ~n590 | n2078 | (~x2 & (n596 | (x4 & ~n2077)));
  assign n2077 = (x3 | x5 | ~x7 | (~x1 ^ x6)) & (x7 | ((~x0 | ((~x5 | x6 | x1 | ~x3) & (~x1 | x3 | x5 | ~x6))) & (x1 | x3 | x5 | x6) & (~x3 | ~x5 | ~x6 | x0 | ~x1)));
  assign n2078 = n601 & (((~x4 ^ x7) & (x6 ? ~x1 : n664)) | (~x4 & x7 & (x6 ? n664 : ~x1)));
  assign z141 = (~n607 & ~n2080) | ~n2085 | (~x3 & (n2081 | ~n2082));
  assign n2080 = (x0 | x3 | x4 | x5 | x6) & (~x3 | ((~x0 | x1 | ~x4 | ~x5 | x6) & (x0 | ((~x5 | x6 | ~x1 | ~x4) & (x5 | ~x6 | x1 | x4)))));
  assign n2081 = n641 & (x2 ? (n738 & ~n824) : (n1156 & n664));
  assign n2082 = ~n2084 & (~n924 | ~n1846) & (~n1901 | ~n2083);
  assign n2083 = x4 & ~x0 & x2;
  assign n2084 = ~x2 & ((x6 & ~x7 & x4 & x5) | (x0 & ~x4 & ~x5 & ~x6 & x7));
  assign n2085 = (~x2 | n2087) & (~n588 | ~n686) & (x2 | n2086);
  assign n2086 = (x3 & ((x0 & (x1 | (x4 & ~x6))) | ~x5 | (x1 & x4 & ~x6))) | (~x5 & ~x6) | (~x3 & x5 & x6) | (~x0 & x1 & ((x4 & ~x5) | (~x3 & ~x4 & ~x6)));
  assign n2087 = (~x0 & ~x4 & (x6 ? ~x5 : ~x3)) | (x5 & (x3 | x4 | ~x6)) | (x0 & x1) | (~x3 & ~x5 & x6);
  assign z142 = n2090 | ~n2092 | n2101 | n2102 | (n738 & ~n2089);
  assign n2089 = (~x5 | x6 | x7 | ~x2 | x3 | ~x4) & (x2 | ((x3 | x4 | x5 | x6 | ~x7) & (~x6 | ((~x5 | x7 | ~x3 | ~x4) & (x3 | (x4 ? (~x5 | ~x7) : (x5 | x7)))))));
  assign n2090 = ~n627 & (x0 ? (~x1 & ~n2091) : (x1 ? (x3 & ~x6) : (~x3 & x6)));
  assign n2091 = x2 ? (~x3 | x6) : (x3 | ~x6);
  assign n2092 = ~n2094 & ~n2097 & ~n2098 & n2099 & (x0 | n2093);
  assign n2093 = (x5 | ~x6 | x7 | x1 | x3 | x4) & (~x1 | ~x3 | ~x4 | ~x5 | x6 | ~x7);
  assign n2094 = n2096 & (x0 ? n2095 : n1449);
  assign n2095 = x4 & ~x5;
  assign n2096 = ~x2 & (x1 ? (~x3 & x6) : (x3 & ~x6));
  assign n2097 = ~n630 & (x0 ? (~x1 & n814) : (x1 & n1956));
  assign n2098 = ~n1875 & ((x0 & ~x1 & x2 & n641) | (~x0 & (x1 ? (~x2 & n641) : (x2 & n642))));
  assign n2099 = ~n2100 & ((x0 & (x1 ^ ~x2)) | (n633 & (~x1 | ~x2 | ~n1773)));
  assign n2100 = ~x6 & x4 & x3 & ~x0 & ~x1;
  assign n2101 = ~n622 & ((~x3 & ~x6 & ((x1 & ~x2) | (~x0 & (x1 | ~x2)))) | (~x0 & x3 & x6 & (~x1 | x2)));
  assign n2102 = ~x4 & ((x0 & ~x1 & ~x2 & x3 & ~x6) | (~x3 & x6 & (x0 ? (~x1 ^ ~x2) : (x1 & x2))));
  assign z143 = (x7 & ~n2104) | (~x4 & ~n2108) | (~x7 & ~n2110) | (x4 & ~n2109);
  assign n2104 = (n783 | n2107) & (x5 | n2106) & (~x5 | ~n732 | n2105);
  assign n2105 = (~x1 | x2 | x4 | x6) & (x1 | ~x2 | ~x4 | ~x6);
  assign n2106 = x0 ? ((x1 | ~x2 | x3 | ~x4 | ~x6) & (~x1 | x2 | ~x3 | x4 | x6)) : (~x1 | x3 | (x2 ? (x4 | x6) : (~x4 | ~x6)));
  assign n2107 = (x0 | x1 | ~x2 | ~x3 | ~x5) & (x5 | ((x2 | ~x3 | x0 | ~x1) & (~x0 | (x1 ? (x2 | x3) : (~x2 | ~x3)))));
  assign n2108 = x5 ? (x7 | (((~x2 & ~x3) | (x0 ^ ~x1)) & (x2 | x3 | (~x0 ^ ~x1)))) : (~x7 | ((x0 | (~x2 ^ ~x3)) & (x1 | (x0 & (x2 | x3)))));
  assign n2109 = (~x3 | ((x2 | ~x7 | ~x0 | x1) & (x0 | x5 | x7))) & (~x0 | ((x1 | ~x5 | ~x7) & (x5 | x7 | x2 | x3))) & (x0 | ((~x1 | ~x5 | ~x7) & (~x2 | x5 | x7))) & (x2 | ((x3 | ~x5 | ~x7) & (x1 | ((~x5 | ~x7) & (x3 | x5 | x7)))));
  assign n2110 = (~n924 | ~n2112) & (~n1937 | (~n2114 & (n2111 | n2113)));
  assign n2111 = x0 ^ ~x5;
  assign n2112 = ~x6 & ~x5 & ~x3 & x4;
  assign n2113 = ~x2 & ~x3;
  assign n2114 = x5 & ~x3 & x0 & ~x2;
  assign z144 = ~n2126 | n2125 | ~n2122 | n2121 | n2116 | n2119;
  assign n2116 = ~x2 & ((n1489 & n983) | n2117 | (~x3 & ~n2118));
  assign n2117 = x0 & ((~x1 & ~x3 & x4 & x5 & x6) | (x1 & x3 & ~x4 & ~x5 & ~x6));
  assign n2118 = (~x5 | x6 | ~x7 | ~x0 | x1 | ~x4) & (x0 | x5 | ((~x4 | x6 | x7) & (~x1 | x4 | ~x6 | ~x7)));
  assign n2119 = ~x1 & ~n2120;
  assign n2120 = (~x5 | ~x6 | ~x7 | ~x0 | ~x2 | ~x3) & (x6 | ((x7 | ((x3 | ~x5 | ~x0 | x2) & ((x2 ^ ~x3) | (~x0 ^ x5)))) & (x2 | ~x7 | ((~x0 | ~x3 | ~x5) & (x5 | (x0 & x3))))));
  assign n2121 = ~x0 & ((x1 & ((x2 & x3 & ~x5) | (x5 & x6 & ~x2 & ~x3))) | (~x5 & x6 & x2 & x3) | (~x1 & ((~x5 & x6 & ~x2 & ~x3) | (x5 & ~x6 & x2 & x3))));
  assign n2122 = ~n2123 & (n2124 | (x1 ? (x2 | x5) : (~x2 | ~x5)));
  assign n2123 = (x2 ^ x3) & ((x5 & x6 & x0 & ~x1) | (~x0 & ~x5 & (~x1 ^ ~x6)));
  assign n2124 = (~x0 | ~x3 | x4 | ~x6 | x7) & (x0 | x3 | ~x4 | x6 | ~x7);
  assign n2125 = n1156 & n1812 & ((x4 & ~x6 & x0 & ~x1) | (~x0 & (x1 ? (x4 & x6) : (~x4 & ~x6))));
  assign n2126 = x1 ? ((~x6 | n2128) & (x2 | x3 | x6 | ~n2127)) : (~n2127 | (x2 ? (~x3 | x6) : (x3 | ~x6)));
  assign n2127 = x0 & ~x5;
  assign n2128 = (x3 | x5 | x7 | x0 | ~x2) & (x2 | (~x5 ^ ~x7) | (~x0 ^ x3));
  assign z145 = n2131 | ~n2132 | n2134 | n2137 | (~n620 & ~n2130);
  assign n2130 = (~x0 | ((~x3 | ~x4 | ~x5 | x1 | ~x2) & (~x1 | x2 | x3))) & (~x1 | ((x2 | x4 | x5) & (x0 | (x3 ? x2 : x4))));
  assign n2131 = x2 & ((x4 & ~x6 & ~x0 & ~x1) | ((x3 ^ x4) & ((~x1 & ~x6) | (~x0 & x1 & x6))));
  assign n2132 = (~x4 | ((~x3 | n2133) & (x6 | ~n897 | ~x1 | x3))) & (x3 | ((x4 | n2133) & (x1 | ~x6 | ~n897)));
  assign n2133 = (~x0 | x1 | x2 | (x6 ^ x7)) & (~x5 | ~x6 | ~x7 | x0 | ~x1 | ~x2);
  assign n2134 = x2 & ((n2135 & n1743) | (~x6 & n738 & ~n2136));
  assign n2135 = x6 & x4 & ~x5;
  assign n2136 = x3 ? (~x4 | x5) : (x4 | ~x5);
  assign n2137 = ~n2138 & ~x1 & ~n662;
  assign n2138 = (x0 | (x2 ? (x3 | x4) : ~x3)) & (~x2 | x3 | x4 | x5) & (x2 | ((~x3 | x4) & (~x0 | x3 | ~x4)));
  assign z146 = ~n2142 | (x5 & (x2 ? ~n2140 : (n664 & n2141)));
  assign n2140 = (~x0 | x1 | x3 | x4 | x6 | x7) & (x0 | ((~x1 | x3 | x4 | (x6 ^ x7)) & (~x3 | ~x4 | ((x6 | ~x7) & (~x1 | ~x6 | x7)))));
  assign n2141 = ~x3 & x7 & (~x4 ^ ~x6);
  assign n2142 = ~n2144 & ~n2145 & (x5 ? (n1403 | ~n2003) : n2143);
  assign n2143 = x4 ? (~x7 | ((x1 | ~x2 | ~x3) & (x0 | ((~x2 | ~x3) & (~x1 | x2 | x3))))) : (x7 | ((~x2 | x3 | x0 | ~x1) & (~x0 | (x1 ? (x2 | ~x3) : (~x2 | x3)))));
  assign n2144 = x2 & ((x7 & (~x0 | ~x1) & (x3 ^ x4)) | (~x0 & ~x1 & ~x3 & ~x4 & ~x7));
  assign n2145 = ~x2 & ((~x0 & ((x3 & ~x7) | (~x1 & ~x3 & x7))) | (~x7 & (x3 ? ~x1 : (x0 | (x1 & ~x4)))));
  assign z147 = ~n2148 | (~x2 & ((~x3 & ~n2147) | (n1229 & n1621)));
  assign n2147 = (x1 | x6 | ((~x0 | ~x4 | (x5 ^ x7)) & (x5 | ~x7 | x0 | x4))) & (x0 | ~x1 | ~x5 | ~x6 | (~x4 ^ ~x7));
  assign n2148 = ~n2151 & n2152 & (~n538 | n2150) & (x0 | n2149);
  assign n2149 = (~x4 | ~x5 | ~x6 | ~x1 | ~x2 | ~x3) & (x4 | ((x1 | ~x2 | ~x3 | x5 | x6) & (x3 | ((x5 | ~x6 | x1 | x2) & (~x1 | ~x5 | (x2 ^ x6))))));
  assign n2150 = (~x5 | x6 | ~x7 | ~x0 | x3 | x4) & (x0 | ~x3 | ~x6 | (x4 ? (~x5 | ~x7) : (x5 | x7)));
  assign n2151 = ~n1446 & (x3 ? (n730 & n664) : (n1365 & n738));
  assign n2152 = (~x0 | ((x2 | x3 | x4) & (~x4 | ~x5 | x1 | ~x2))) & ((x0 & x1) | (x2 ? (x3 | ~x4) : (~x3 | x4))) & (x2 | x5 | ((~x1 | x3 | x4) & (x0 | x1 | ~x3)));
  assign z148 = ~n2158 | ~n2163 | (x0 ? (~x1 & ~n2162) : ~n2154);
  assign n2154 = x4 ? ((~n2155 | ~n742) & (n1429 | n2156)) : n2157;
  assign n2155 = ~x7 & x5 & ~x6;
  assign n2156 = x1 ? (x2 | x3) : (~x2 | ~x3);
  assign n2157 = (~x1 | x2 | x3 | ~x5 | (x6 ^ x7)) & (x5 | ~x6 | ~x7 | x1 | ~x2 | ~x3);
  assign n2158 = (~x6 | n2161) & (n868 | n2160) & (x1 | x6 | n2159);
  assign n2159 = ((x3 ? (x4 | ~x5) : (~x4 | x5)) | (~x0 ^ ~x2)) & (x3 | x4 | x5 | (x0 ^ ~x2));
  assign n2160 = (~x2 | ~x3 | ~x6 | x0 | ~x1) & (~x0 | x2 | x6 | (~x1 ^ x3));
  assign n2161 = x0 ? (x1 | ((x2 | ~x4 | x5) & (x4 | ~x5 | ~x2 | x3))) : (~x1 | ((x2 | ~x3 | ~x4 | x5) & (x4 | ~x5 | ~x2 | x3)));
  assign n2162 = (~x5 | x6 | ~x7 | ~x2 | x3 | x4) & (x2 | ((~x6 | x7 | x4 | x5) & (~x4 | ((~x6 | x7 | ~x3 | ~x5) & (x5 | x6 | ~x7)))));
  assign n2163 = x2 ? ((~x4 | x5 | x0 | x3) & (~x3 | (x0 ? (x1 | (x4 ^ x5)) : (x4 | ~x5)))) : ((x3 | ((x4 | ~x5 | x0 | x1) & (~x0 | ~x4 | (x1 ^ ~x5)))) & (x0 | ((~x1 | x4 | x5) & (~x3 | (x4 ^ x5)))));
  assign z149 = n2165 | ~n2168 | n2173 | (x0 & ~n2172);
  assign n2165 = ~x7 & (x3 ? ~n2167 : ~n2166);
  assign n2166 = (~x6 | (x0 ? ((~x1 | x2 | ~x4 | x5) & (x4 | ~x5 | x1 | ~x2)) : (x4 | ((x2 | ~x5) & (~x1 | ~x2 | x5))))) & (~x5 | x6 | (x0 ? (x1 ? (x2 | x4) : (~x2 | ~x4)) : (x1 | (~x2 ^ x4))));
  assign n2167 = (x0 | ~x1 | ~x4 | (x2 ? (x5 | ~x6) : (~x5 | x6))) & (x4 | ((x5 | ((x2 | ~x6 | x0 | x1) & (~x0 | (x1 ? (x2 | x6) : (~x2 | ~x6))))) & (x0 | ~x1 | ~x2 | ~x5 | x6)));
  assign n2168 = (x0 | n2169) & (n846 | (n2170 & n2171));
  assign n2169 = (~x1 | (x2 ? ((x3 | ~x4 | ~x5 | x6) & (x5 | ~x6 | ~x3 | x4)) : (x4 ? (x5 | ~x6) : (x6 | (x3 ^ x5))))) & (x2 | x3 | ~x4 | x5 | ~x6) & (x1 | ((~x2 | ~x3 | x4 | ~x5 | x6) & ((~x3 ^ ~x4) | (x2 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n2170 = x0 ? ((~x3 | x4 | x1 | ~x2) & (~x1 | x2 | x3 | ~x4)) : ((x1 | x2 | ~x3 | x4) & (~x2 | (x1 ? (~x3 ^ ~x4) : (x3 | ~x4))));
  assign n2171 = (~x4 | (((~x2 ^ x7) | (x0 ? (x1 | ~x3) : (~x1 | x3))) & (x0 | x1 | ~x3 | (~x2 ^ ~x7)))) & (x0 | ~x1 | x2 | ~x3 | x4 | x7);
  assign n2172 = (~x1 | x2 | x3 | x4 | x5 | ~x6) & (x1 | ((x6 | (x2 ? (x3 ? (~x4 | ~x5) : (x4 | x5)) : (x4 | ~x5))) & (~x4 | ~x6 | ((x3 | x5) & (x2 | (x3 & x5))))));
  assign n2173 = x7 & ((n1121 & n690 & n924) | (~x1 & ~n2174));
  assign n2174 = (~x2 | ((x4 | ~x5 | x6 | ~x0 | x3) & (x0 | ((x3 | ~x4 | ~x5 | x6) & (x5 | ~x6 | ~x3 | x4))))) & (~x0 | x2 | ((x4 | x5 | ~x6) & (x3 | ~x4 | x6)));
  assign z150 = n2177 | n2180 | (~n2176 & ~n2185) | (~n662 & ~n2186);
  assign n2176 = x4 ? (~x6 | x7) : (x6 | ~x7);
  assign n2177 = x5 & (x3 ? ~n2179 : ~n2178);
  assign n2178 = (x4 | (x0 ? (x1 | ~x6 | (~x2 ^ ~x7)) : (~x1 | (x2 ? x7 : (x6 | ~x7))))) & (x1 | ~x4 | x6 | (~x7 & (~x0 | x2)));
  assign n2179 = (~x6 | x7 | x1 | x4) & (x0 | ~x4 | x6 | ~x7 | (x1 ^ ~x2));
  assign n2180 = ~x5 & ((x2 & ~n2182) | (~n2181 & ~n2183) | (~x2 & ~n2184));
  assign n2181 = x3 ? (x6 | ~x7) : (~x6 | x7);
  assign n2182 = (x1 | x3 | x4 | ~x6 | x7) & (x0 | ~x1 | ((x3 | x6 | ~x7) & (~x6 | x7 | ~x3 | x4)));
  assign n2183 = (x1 | ~x2 | ~x4) & (~x0 | ~x1 | x2 | x4);
  assign n2184 = (x0 | ((~x6 | x7 | x3 | x4) & (~x1 | ((x4 | ~x6 | x7) & (x3 | ~x4 | x6 | ~x7))))) & (x1 | ~x4 | x6 | ~x7 | (~x0 & ~x3));
  assign n2185 = x1 ? ((x3 | ~x5 | ~x0 | x2) & (x0 | ~x3 | (x2 & ~x5))) : ((~x2 | (~x3 ^ x5)) & (x3 | (x5 ? x0 : x2)));
  assign n2186 = x5 ? ((x0 | ~x1 | ((x3 | ~x4) & (x2 | ~x3 | x4))) & (x1 | ((x2 | x3 | x4) & (~x3 | (~x2 & ~x4))))) : ((~x0 | x2 | (x1 ? (x3 | ~x4) : x4)) & (x0 | (x1 ? ((~x2 | x3 | x4) & (~x3 | ~x4)) : (x3 | ~x4))) & (x1 | ((~x3 | x4) & (~x2 | x3 | ~x4))));
  assign z151 = ~n2188 | (x1 ? ~n2193 : (x3 ? ~n2191 : ~n2192));
  assign n2188 = (n662 | n2190) & (n1465 | (x2 ? n1799 : n2189));
  assign n2189 = x0 ^ ~x3;
  assign n2190 = (~x2 & ((~x1 & x4) | (~x0 & (x4 | (~x1 & ~x3 & ~x5))))) | (x2 & ((~x4 & x5) | (x0 & x1))) | (x0 & (x3 ? x1 : (~x4 & x5))) | (x4 & ~x5) | (~x4 & x5 & x1 & ~x3);
  assign n2191 = x5 ? ((x6 | ~x7 | x2 | ~x4) & (~x0 | ((~x4 | x6 | ~x7) & (x2 | x4 | ~x6 | x7)))) : ((x0 | ~x2 | x4 | ~x6 | x7) & (x2 | (x4 ? (~x6 | x7) : (x6 | ~x7))));
  assign n2192 = (x5 | ((x0 | ((x2 | x4 | ~x7) & (~x4 | ~x6 | x7))) & (~x6 | x7 | ((~x2 | ~x4) & (~x0 | x2 | x4))))) & (x6 | ~x7 | ~x4 | ~x5) & (~x0 | ((~x2 | x4 | ~x5 | ~x6 | ~x7) & (x2 | ((~x5 | x6 | ~x7) & (~x4 | x7 | (~x5 & x6))))));
  assign n2193 = (x4 | n2194) & (n630 | ((x2 | x3 | x4) & (x0 | ~x4 | (x2 & x3))));
  assign n2194 = (~x5 | ~x6 | ~x7 | x0 | x3) & (x2 | ((~x0 | ~x3 | x5 | ~x6 | x7) & (x0 | ((x3 | ~x5 | ~x6) & (x6 | ~x7 | ~x3 | x5)))));
  assign z152 = ~n2201 | (x2 ? ~n2196 : (x0 ? ~n2200 : ~n2199));
  assign n2196 = x0 ? (x1 | n2198) : n2197;
  assign n2197 = (x4 | ((~x1 | ~x6 | x7 | (x3 ^ x5)) & (~x5 | x6 | ~x7 | (x1 & ~x3)))) & (~x7 | ((~x3 | x5 | ~x6) & (~x4 | ((x5 | ~x6) & (x3 | ~x5 | x6)))));
  assign n2198 = (x3 | x4 | x5 | ~x6 | x7) & (~x7 | ((~x4 | ~x5 | x6) & (~x3 | (~x5 ^ x6))));
  assign n2199 = (x4 | ((x1 | ~x3 | x5 | x6 | ~x7) & (~x1 | x3 | (x5 ? (~x6 | ~x7) : (x6 | x7))))) & (x7 | ((~x4 | ~x5 | x6) & (~x3 | (~x5 ^ x6))));
  assign n2200 = (x5 | ((~x6 | x7 | x1 | ~x3) & (x6 | ((~x1 | (x3 ? (x4 | ~x7) : (~x4 | x7))) & (x1 | ~x3 | ~x4 | ~x7))))) & (x1 | ~x5 | ((~x3 | x6 | x7) & (~x6 | ~x7 | x3 | ~x4)));
  assign n2201 = ~n2203 & ~n2204 & n2206 & (n846 | n2202);
  assign n2202 = x2 ? (~x3 | x7 | ((x1 | ~x4) & (x0 | (x1 & ~x4)))) : ((x4 | ((~x3 | ~x7 | x0 | ~x1) & (~x0 | ((x3 | x7) & (x1 | ~x3 | ~x7))))) & (x0 | x3 | ~x7 | (x1 & ~x4)));
  assign n2203 = ~n857 & ((x2 & ~x5 & ~x7 & (~x3 ^ ~x4)) | (x7 & ((~x4 & x5 & x2 & ~x3) | (~x2 & (x3 ? (x4 & x5) : (~x4 & ~x5))))));
  assign n2204 = n563 & ((n738 & n828) | (n2205 & (n1119 | n1123)));
  assign n2205 = x5 & ~x7;
  assign n2206 = (x3 | x5 | ~x7 | ~x0 | ~x1 | x2) & (x0 | x1 | ((~x5 | ~x7 | x2 | ~x3) & (x5 | x7 | ~x2 | x3)));
  assign z153 = ~n2213 | (x2 ? ~n2208 : (x5 ? ~n2212 : ~n2211));
  assign n2208 = (n846 | n2210) & (~x0 | ~n605 | ~n678) & (x0 | n2209);
  assign n2209 = x5 ? (x6 | ((~x3 | x4 | x7) & (~x1 | x3 | ~x4 | ~x7))) : ((x4 | ((~x6 | ~x7 | x1 | x3) & (~x1 | x7 | (x3 ^ x6)))) & (x1 | ~x3 | ~x4 | x6 | ~x7));
  assign n2210 = (x3 | x4 | x7 | ~x0 | x1) & (~x3 | ~x4 | ~x7 | x0 | ~x1);
  assign n2211 = x0 ? (x1 ? (x7 | (x3 ? (x4 | ~x6) : (~x4 | x6))) : (~x4 | ~x7 | (~x3 ^ x6))) : ((x1 | ~x3 | x4 | x6 | ~x7) & (x3 | ((~x4 | ~x6 | x7) & (~x1 | x4 | (x6 ^ x7)))));
  assign n2212 = (x0 | ~x1 | x3 | x4 | ~x6 | x7) & (x1 | ((x6 | (x0 ? (x3 ? (x4 | x7) : (~x4 | ~x7)) : (x3 | (~x4 ^ x7)))) & (x0 | ~x3 | ~x6 | (~x4 ^ x7))));
  assign n2213 = n2217 & (n662 | n2216) & (x2 ? n2215 : n2214);
  assign n2214 = (~x4 | x6 | ~x7 | x0 | x3) & (x1 | (x0 ? ((x3 | ~x4 | ~x6 | x7) & (x6 | ~x7 | ~x3 | x4)) : (x4 | x7 | (~x3 ^ x6))));
  assign n2215 = (x1 | (x6 ? ((~x0 | x4 | (~x3 ^ x7)) & (x3 | x7 | (x0 & ~x4))) : (~x7 | ((~x3 | x4) & (x0 | x3 | ~x4))))) & (x0 | ((x3 | ~x4 | ~x6 | x7) & (~x3 | x6 | ((x4 | ~x7) & (~x1 | ~x4 | x7)))));
  assign n2216 = (x3 | x4 | ~x0 | x2) & (~x3 | ~x4 | ((x1 | x2) & (x0 | (x1 & x2))));
  assign n2217 = x0 ? (~x4 | ((x3 | ~x6 | ~x1 | x2) & (~x3 | x6 | x1 | ~x2))) : (~x1 | x4 | (x2 ? (x3 | ~x6) : (~x3 | x6)));
  assign z154 = ~n2224 | (x3 ? ~n2219 : (x1 ? ~n2223 : ~n2222));
  assign n2219 = x1 ? n2220 : n2221;
  assign n2220 = (~x0 | x2 | x4 | x5 | x6 | ~x7) & (x0 | ~x2 | ~x4 | ~x5 | ~x6 | x7);
  assign n2221 = x4 ? ((~x0 | x2 | x5 | x6 | ~x7) & (x0 | (x2 ? (x5 | (~x6 ^ x7)) : (~x5 | (x6 ^ x7))))) : ((x7 | ((x0 | (x2 ? (x5 | x6) : (~x5 | ~x6))) & (x5 | x6 | ~x0 | x2))) & (~x0 | ~x6 | ~x7 | (x2 ^ x5)));
  assign n2222 = (~x7 | ((~x5 | ((x0 | ~x2 | x4 | x6) & (~x0 | (x2 ? (~x4 | x6) : (x4 | ~x6))))) & (x0 | x2 | x5 | (x4 ^ x6)))) & (~x6 | x7 | ((~x0 | ~x4 | ~x5) & (x0 | x2 | x4 | x5)));
  assign n2223 = (x5 | (((~x4 ^ ~x7) | (x0 ? (x2 | ~x6) : (~x2 | x6))) & (~x0 | x2 | ~x4 | x6 | x7))) & (x0 | x2 | ~x5 | (x4 ? (x6 ^ x7) : (x6 | ~x7)));
  assign n2224 = ~n2225 & ~n2226 & ~n2228 & (x3 | n2227);
  assign n2225 = ~n592 & ((x0 & ~x1 & ~x2 & x3 & x5) | (~x0 & ((x1 & (x2 ? (~x3 & x5) : x3)) | (~x2 & x3 & ~x5) | (~x1 & x2 & (x3 ^ ~x5)))));
  assign n2226 = ~n927 & (x0 ? ((x1 & ~x2 & ~x3 & x5) | (~x1 & (x3 ? x2 : ~x5))) : ((~x1 & ~x2 & ~x3 & x5) | (x3 & ~x5 & x1 & x2)));
  assign n2227 = (x1 | ~x5 | ((~x4 | x7 | x0 | ~x2) & (~x0 | x4 | (~x2 ^ ~x7)))) & (x0 | x5 | ((x2 | ~x4 | x7) & (~x1 | (x2 ? (x4 | ~x7) : x7))));
  assign n2228 = x7 & n650 & n616 & (x1 ^ ~x5);
  assign z155 = n2230 | n2234 | n2239 | ~n2240 | (~x5 & ~n2233);
  assign n2230 = ~x2 & (x0 ? ~n2231 : ~n2232);
  assign n2231 = (~x6 | (x1 ? ((~x5 | ~x7 | x3 | ~x4) & (~x3 | x4 | x5 | x7)) : (x7 | (x3 ? (~x4 | x5) : (x4 | ~x5))))) & (~x1 | x3 | x4 | x6 | (x5 ^ x7));
  assign n2232 = (x1 | ((x5 | ~x6 | x7 | x3 | ~x4) & (x6 | ((x3 | x4 | x5 | ~x7) & (~x3 | (x4 ? (x5 | ~x7) : (~x5 | x7))))))) & (x5 | ~x6 | ~x7 | ~x1 | ~x3 | x4);
  assign n2233 = (~x3 | x4 | x6 | ~x0 | x2) & (~x6 | ((x0 | ~x1 | ~x4 | (~x2 ^ ~x3)) & (x1 | ((x0 | x2 | ~x3 | ~x4) & (~x0 | x3 | (x2 ^ x4))))));
  assign n2234 = x2 & ((n586 & n1166) | n2236 | (~x0 & ~n2235));
  assign n2235 = (x5 | ~x6 | x7 | ~x1 | x3 | ~x4) & ((x1 ^ ~x3) | ((x6 | x7 | x4 | x5) & (~x6 | ~x7 | ~x4 | ~x5)));
  assign n2236 = ~n800 & ((x0 & ~x1 & x3 & n2237) | (~x0 & (x1 ? (x3 & n2238) : (~x3 & n2237))));
  assign n2237 = ~x4 & x6;
  assign n2238 = x4 & ~x6;
  assign n2239 = n1121 & ((~x0 & x1 & ~x2 & ~x3 & x4) | (~x1 & (x0 ? (x2 ? (x3 ^ x4) : (~x3 & ~x4)) : (x2 ? (~x3 & ~x4) : (x3 & x4)))));
  assign n2240 = ~n2242 & ~n2243 & (~n534 | ~n1838) & (n2241 | n1475);
  assign n2241 = x3 ? (~x4 | ~x5) : (x4 | x5);
  assign n2242 = ~x0 & ((~x1 & x2 & ~x3 & x4 & x5) | (x3 & ~x4 & (x1 ? (x2 ^ x5) : (~x2 & ~x5))));
  assign n2243 = ~n1716 & ((~x0 & ~x1 & ~x2 & ~x3) | ((x1 ^ x3) & (x0 ^ x2)));
  assign z156 = ~n2247 | ~n2252 | (~n1041 & ~n2245) | (~x0 & ~n2246);
  assign n2245 = x1 ? ((x5 | ~x7 | x2 | x3) & (x0 | (x2 ? (~x3 | x7) : (x3 | ~x5)))) : ((~x3 | x5 | ~x7 | x0 | ~x2) & ((x5 ^ x7) | (x0 ? (~x2 | x3) : (x2 | ~x3))));
  assign n2246 = x1 ? ((~x2 | x3 | x4 | ~x5 | x6) & (~x4 | x5 | ~x6 | x2 | ~x3)) : ((x2 | x3 | x4 | ~x5 | x6) & (~x2 | ((x3 | ~x4 | ~x6) & (~x5 | x6 | ~x3 | x4))));
  assign n2247 = x1 ? n2248 : (n2250 & (~x0 | (n2249 & n2251)));
  assign n2248 = (x0 | ((~x5 | ~x6 | ~x7 | x2 | ~x3) & (~x2 | x5 | (x3 ? (~x6 | ~x7) : (x6 | x7))))) & (~x0 | x2 | x3 | x6 | x7);
  assign n2249 = x2 ? (x6 | x7 | (x3 ? (x4 | x5) : (~x4 | ~x5))) : (~x4 | ~x6 | ~x7 | (x3 & ~x5));
  assign n2250 = (x5 | ~x6 | ~x7 | ~x0 | ~x2 | x3) & (x0 | ~x3 | x6 | x7 | (~x2 ^ x5));
  assign n2251 = (~x2 | ~x3 | ~x4 | ~x6) & (x2 | x4 | x6 | (~x3 & x5));
  assign n2252 = (n620 | n2253) & (x0 | (x1 ? n2254 : n2255));
  assign n2253 = (x3 | (((x1 ^ x4) | (x0 ? (x2 | ~x5) : ~x2)) & (x1 | x2 | ~x4 | (x0 & x5)))) & (x0 | ~x1 | x2 | x4 | x5) & (~x3 | (x1 ? (x2 | x4 | (x0 & x5)) : ((~x0 | (~x2 ^ x4)) & (~x4 | ~x5 | x0 | ~x2))));
  assign n2254 = (x5 | x6 | x7 | x2 | x3 | ~x4) & (~x5 | ~x6 | ~x7 | ~x2 | ~x3 | x4);
  assign n2255 = (~x2 | x3 | x4 | x5 | x6 | x7) & (x2 | ~x7 | ((~x3 | x4 | x5 | ~x6) & (x3 | (x4 ? (~x5 | ~x6) : (x5 | x6)))));
  assign z157 = n2261 | ~n2264 | (x2 & (~n2257 | ~n2260));
  assign n2257 = x4 ? n2259 : n2258;
  assign n2258 = (x1 | ((x7 | ((~x5 | x6 | x0 | ~x3) & (~x6 | (x0 ? (~x3 ^ x5) : (x3 | x5))))) & (~x0 | ~x3 | x5 | x6 | ~x7))) & (x0 | ~x1 | ((~x6 | ~x7 | x3 | x5) & (~x3 | x6 | (x5 ^ x7))));
  assign n2259 = (~x0 | x1 | ~x3 | x5 | x6 | x7) & (x0 | x3 | ((x6 | ~x7 | x1 | ~x5) & (~x1 | x5 | (~x6 ^ x7))));
  assign n2260 = ((x0 ? (x1 | ~x4) : (~x1 | x4)) | (x3 ? (x5 | ~x7) : (x5 ^ x7))) & (~x0 | x1 | x3 | x4 | x5 | ~x7) & (x0 | ((~x4 | ((x1 | x3 | x5 | ~x7) & (x7 | (x1 ? (~x3 ^ x5) : (~x3 | ~x5))))) & (x1 | x4 | ~x5 | (~x3 ^ ~x7))));
  assign n2261 = ~x2 & (x3 ? ~n2263 : ~n2262);
  assign n2262 = (~x5 | x6 | ~x7 | x0 | x4) & (~x4 | ((~x0 | ~x6 | ((~x5 | x7) & (x1 | x5 | ~x7))) & (x0 | ~x1 | x5 | x6 | x7)));
  assign n2263 = (x0 | ~x1 | ~x4 | ~x5 | ~x6 | x7) & (x1 | ((x5 | ~x6 | ~x7 | x0 | ~x4) & (~x0 | ((x6 | x7 | x4 | x5) & (~x6 | ~x7 | ~x4 | ~x5)))));
  assign n2264 = (x2 | n2267) & (n927 | n2266) & (n662 | n2265);
  assign n2265 = (x3 | x4 | ~x5 | ~x0 | ~x1 | x2) & (x0 | ((x1 | x2 | x3 | ~x4 | ~x5) & (~x1 | ((~x4 | ~x5 | ~x2 | ~x3) & (x2 | x4 | (x3 ^ x5))))));
  assign n2266 = x0 ? ((x1 | ~x2 | ~x3 | ~x5) & (~x1 | x2 | x3 | x5)) : (~x3 | (x1 ? (x2 | x5) : (~x2 ^ x5)));
  assign n2267 = x1 ? ((~x4 | ~x7 | x0 | x3) & (~x0 | ~x3 | x4 | x5 | x7)) : ((x4 | ~x5 | x7 | ~x0 | x3) & ((~x4 ^ x7) | (x5 & (~x0 | ~x3))));
  assign z158 = n2269 | ~n2272 | n2275 | n2278 | (~n2189 & ~n2271);
  assign n2269 = ~x0 & ~n2270;
  assign n2270 = x5 ? (x1 ? ((x3 | x4 | x6) & (~x4 | ~x6 | x2 | ~x3)) : (~x3 | (x4 ? x6 : x2))) : ((~x6 | ((~x1 | ((x3 | ~x4) & (~x2 | ~x3 | x4))) & (x3 | x4 | (x1 & x2)))) & (x1 | ~x2 | x3 | ~x4 | x6));
  assign n2271 = (x2 | (x1 ? ((~x6 | x7 | x4 | x5) & (x6 | ~x7 | ~x4 | ~x5)) : (x5 | (x4 ? (~x6 | ~x7) : (x6 | x7))))) & (x1 | ~x2 | ((x4 | ~x5 | x6 | ~x7) & (~x4 | x7 | (~x5 ^ ~x6))));
  assign n2272 = (n846 | n2273) & (~n738 | n2274);
  assign n2273 = (x3 | ((~x0 | (x1 ? x2 : (~x2 | x4))) & (x0 | x1 | x2 | ~x4))) & (x0 | ~x3 | (x1 ? (x2 ^ x4) : (~x2 | x4)));
  assign n2274 = x3 ? ((~x2 | ((x5 | ~x6) & (x4 | ~x5 | x6))) & (x5 | ((x4 | ~x6) & (x2 | ~x4 | x6)))) : (~x5 | (x4 ? x6 : x2));
  assign n2275 = ~x4 & (n2277 | (~n846 & ~n2276 & ~x0 & x7));
  assign n2276 = x1 ? (~x2 | ~x3) : (x2 | x3);
  assign n2277 = ~n800 & ((x0 & ~x1 & ~x2 & x3 & ~x6) | (~x0 & x2 & ~x3 & (~x1 ^ x6)));
  assign n2278 = x4 & ((~x1 & ~n2279) | (~x6 & n664 & ~n2280));
  assign n2279 = (~x0 | ~x2 | ~x3 | x5 | x6 | ~x7) & (~x6 | (x5 ^ x7) | (x0 ? (x2 | ~x3) : (~x2 | x3)));
  assign n2280 = (~x5 | x7 | ~x2 | x3) & (x2 | x5 | (~x3 ^ x7));
  assign z159 = ~n2282 | ~n2296 | (~n846 & ~n2295) | (x2 & ~n2294);
  assign n2282 = ~n2283 & n2287 & ~n2291 & ~n2293 & (x0 | n2284);
  assign n2283 = ~n1361 & ((~x3 & ~x5 & ~x6 & ~x0 & x2) | (~x2 & (x0 ? (x3 ? (~x5 & ~x6) : (x5 & x6)) : (x6 & (x3 ^ ~x5)))));
  assign n2284 = (~n709 | n2286 | x6 | ~x7) & (~x6 | x7 | ~n1701 | ~n2285);
  assign n2285 = ~x3 & x1 & x2;
  assign n2286 = x2 ? (~x3 | ~x4) : (x3 | x4);
  assign n2287 = (n2289 | n2290) & (~n698 | ~n1476) & (~n924 | ~n2288);
  assign n2288 = ~x7 & ~x6 & x3 & ~x4;
  assign n2289 = x2 ? (x5 | ~x6) : (~x5 | x6);
  assign n2290 = (~x0 | x1 | x3 | x4) & (x0 | (x1 ? (x3 | ~x4) : (~x3 | x4)));
  assign n2291 = ~n1019 & ((~x0 & x2 & ~x3 & ~n945) | (~x2 & ((x3 & ~n2292) | (x0 & ~x3 & ~n945))));
  assign n2292 = x0 ? (x1 | x7) : (~x1 | ~x7);
  assign n2293 = ~n783 & ((~x0 & ~x1 & x2 & ~x3 & x7) | (x0 & ~x2 & (x1 ? (~x3 & ~x7) : (x3 & x7))));
  assign n2294 = x0 ? (x1 | ((~x4 | ~x5 | x6) & (x5 | ~x6 | ~x3 | x4))) : (~x1 | ~x3 | (x4 ? (x5 | ~x6) : (~x5 | x6)));
  assign n2295 = (~x2 | (x0 ? (x1 | (x3 ? (x4 | x7) : (~x4 | ~x7))) : (~x1 | ~x3 | (~x4 ^ x7)))) & (x0 | x2 | x3 | x7 | (~x1 ^ x4));
  assign n2296 = x6 ? (x7 ? n2297 : n2298) : (x7 ? n2298 : n2297);
  assign n2297 = (x3 | ~x4 | x5 | ~x0 | x1 | x2) & (x0 | ((x1 | x2 | ~x3 | ~x4 | x5) & (~x5 | ((x1 | (x2 ? (~x3 | ~x4) : (x3 | x4))) & (x3 | x4 | ~x1 | ~x2)))));
  assign n2298 = (x0 | ~x1 | x2 | ~x4 | x5) & (x1 | ((x0 | x2 | ~x3 | x4 | x5) & (~x2 | ((~x0 | (x3 ? (~x4 | x5) : (x4 | ~x5))) & (x4 | ~x5 | x0 | ~x3)))));
  assign z160 = ~n2307 | (x3 ? (~n2301 | (~x0 & ~n2300)) : ~n2302);
  assign n2300 = x2 ? ((x1 | ~x4 | ~x5 | x6 | x7) & (~x6 | ((x5 | x7 | x1 | ~x4) & (~x1 | x4 | (x5 ^ x7))))) : ((x1 | x4 | x5 | x6 | ~x7) & (~x1 | ~x5 | (x4 ? (x6 | ~x7) : (~x6 | x7))));
  assign n2301 = (~x0 | x1 | (x2 ? ~n686 : (~x7 | n850))) & (x0 | ~x1 | ~x2 | x7 | n850);
  assign n2302 = (n2305 | ~n2306) & (n912 | n2303) & (~n1421 | n2304);
  assign n2303 = (~x4 | ((x0 | x1 | ~x2 | ~x7) & (~x0 | (x1 ? (x2 | ~x7) : (~x2 | x7))))) & (x0 | ((x1 | x2 | x7) & (x4 | ~x7 | ~x1 | ~x2)));
  assign n2304 = (x0 | ~x2 | x4 | x6 | ~x7) & (~x0 | ~x4 | ~x6 | (x2 ^ x7));
  assign n2305 = (~x0 | ~x4 | x6 | x7) & (x0 | (x4 ? (x6 | ~x7) : (~x6 | x7)));
  assign n2306 = ~x5 & x1 & ~x2;
  assign n2307 = ~n2310 & ~n2311 & (n846 | n2308) & (x0 | n2309);
  assign n2308 = x3 ? ((~x2 ^ ~x7) | (x0 ? (x1 | x4) : (~x1 | ~x4))) : ((x0 | x1 | ~x2 | x4 | x7) & (x2 | ((x0 | ~x7 | (~x1 ^ x4)) & (x4 | x7 | ~x0 | ~x1))));
  assign n2309 = x3 ? ((x1 | ~x5 | (x2 ? ~x7 : (~x4 | x7))) & (x2 | x5 | ~x7 | (~x1 & ~x4))) : (x7 | ((~x2 | ~x4 | x5) & (~x1 | (~x2 ^ x5))));
  assign n2310 = ~n906 & (x1 ? ((~x4 & ~x5 & x0 & ~x2) | (x4 & x5 & ~x0 & x2)) : (x0 ? (x2 ? (~x4 & x5) : (x4 & ~x5)) : (~x4 & (x2 ^ x5))));
  assign n2311 = n738 & (((x3 ? (x4 & x7) : (~x4 & ~x7)) & (x2 ^ x5)) | (x2 & x3 & x4 & x5 & ~x7) | (~x5 & x7 & ~x2 & ~x4));
  assign z161 = n2313 | n2316 | ~n2321 | ~n2330 | (~n620 & ~n2320);
  assign n2313 = x1 & ((n559 & n2314) | (~x0 & ~n2315));
  assign n2314 = x3 & x0 & ~x2;
  assign n2315 = (~x5 | ~x6 | ~x7 | x2 | x3 | x4) & (~x4 | ((~x3 | ((x6 | ~x7 | x2 | x5) & (~x2 | ~x5 | (x6 ^ x7)))) & (x2 | x3 | x5 | ~x6 | ~x7)));
  assign n2316 = ~x1 & ((n2317 & n698) | n2319 | (x2 & ~n2318));
  assign n2317 = ~x3 & ~x0 & ~x2;
  assign n2318 = (~x0 | x3 | x4 | ~x5 | ~x6 | x7) & (x0 | ((~x3 | ~x4 | ~x5 | x6 | ~x7) & (x3 | x4 | x5 | ~x6 | x7)));
  assign n2319 = ~n662 & ((~x0 & ((x2 & ~x3 & x4 & x5) | (~x4 & ~x5 & ~x2 & x3))) | (x0 & x2 & x3 & ~x4 & x5));
  assign n2320 = ((~x2 ^ x5) | ((~x3 | x4 | x0 | ~x1) & (x3 | ~x4 | ~x0 | x1))) & (x3 | x4 | x5 | ~x0 | ~x1 | x2) & (x0 | x1 | ((x4 | ~x5 | x2 | x3) & (~x4 | x5 | ~x2 | ~x3)));
  assign n2321 = ~n2323 & ~n2324 & ~n2325 & n2329 & (n557 | n2322);
  assign n2322 = x2 ? (x3 | x6) : (~x3 | ~x6);
  assign n2323 = ~x1 & ((~x0 & ~x2 & ~x3 & x4 & x6) | (x3 & ~x6 & (x0 ? (x2 & x4) : (x2 ^ x4))));
  assign n2324 = ~n627 & ((x2 & x3 & x6 & ~x0 & x1) | (x0 & ~x2 & ~x3 & (~x1 ^ x6)));
  assign n2325 = n2328 & ((n537 & n2327) | (n2326 & n540));
  assign n2326 = ~x2 & x4;
  assign n2327 = x2 & ~x4;
  assign n2328 = ~x3 & ~x0 & x1;
  assign n2329 = (~n814 | ~n534 | ~n540) & (~n924 | ~n1112);
  assign n2330 = (x4 | x6 | n2332) & (~x6 | (n2331 & (~x4 | n2332)));
  assign n2331 = (x0 | ~x1 | x2 | x3 | x4 | x5) & (x1 | ~x2 | (x0 ? (x3 ? (x4 | x5) : (~x4 | ~x5)) : (~x5 | (~x3 ^ ~x4))));
  assign n2332 = (x3 | (x0 ? (x2 | (x1 ? (~x5 | ~x7) : (x5 | x7))) : (~x2 | (x1 ? (~x5 | x7) : (x5 | ~x7))))) & (x1 | x2 | ~x3 | (x0 ? (x5 | ~x7) : (~x5 | x7)));
  assign z162 = n2334 | n2339 | (~n800 & ~n2338) | (~n824 & ~n2337);
  assign n2334 = ~x0 & (x1 ? ~n2335 : ~n2336);
  assign n2335 = x2 ? ((x6 | ~x7 | x4 | x5) & (x3 | (x4 ? (x6 | x7) : (~x6 | ~x7)))) : ((~x3 | ~x4 | ~x5 | ~x6 | x7) & (x3 | x6 | (x4 ? ~x7 : (~x5 | x7))));
  assign n2336 = x4 ? (x2 ? (~x7 | (~x3 ^ x6)) : (x7 | (x6 ? x3 : ~x5))) : ((~x3 | (x2 ? (~x5 | x7) : (x6 | ~x7))) & (x2 | ~x7 | (~x5 ^ x6)));
  assign n2337 = x4 ? ((x2 | (x0 ? (x3 | (~x1 & x6)) : (x1 | ~x3))) & (x0 | ~x2 | (~x1 ^ (~x3 & ~x6)))) : ((x0 | ((x2 | x3 | ~x6) & (~x1 | (x2 & (x3 | x6))))) & (x1 | ~x2 | (~x0 & (~x3 | ~x6))));
  assign n2338 = x2 ? ((x3 | ~x4 | ~x0 | x1) & (x0 | ((x4 | ~x6 | ~x1 | ~x3) & (x1 | (x3 ? (~x4 | ~x6) : x4))))) : (x0 ? (x4 | (x1 ? (x3 | ~x6) : x6)) : (~x1 | ~x4 | (~x3 ^ x6)));
  assign n2339 = x0 & ((~n592 & ~n2340) | n2342 | (~x2 & ~n2341));
  assign n2340 = (~x1 | x2 | x3 | ~x5 | x6) & (x1 | ~x2 | ~x3 | x5 | ~x6);
  assign n2341 = (x4 | ((x1 | ~x6 | x7) & (x6 | ~x7 | ~x1 | x5))) & (x1 | ~x4 | ~x7 | (x5 & (x3 | ~x6) & (~x3 | x6)));
  assign n2342 = n2205 & n538 & (x3 ? x4 : (~x4 & ~x6));
  assign z163 = ~n2352 | (~x2 & (~n2345 | (~x1 & ~n2344)));
  assign n2344 = (x0 | ~x3 | x4 | ~x5 | ~x6 | x7) & (x3 | ((x5 | ~x6 | x7 | x0 | x4) & (x6 | ((~x5 | x7 | ~x0 | ~x4) & (x0 | x5 | (~x4 ^ x7))))));
  assign n2345 = ~n2346 & n2350 & ((~x0 & ~n723) | n2349 | (x0 & ~n691));
  assign n2346 = ~n2348 & (n2347 | (n690 & n543));
  assign n2347 = x3 & (x4 ? (x6 & ~x7) : (~x6 & x7));
  assign n2348 = x0 ? (x1 | ~x5) : (~x1 | x5);
  assign n2349 = (~x4 | x6 | x1 | x3) & (x4 | ~x6 | ~x1 | ~x3);
  assign n2350 = (~x0 | ~x1 | x3 | n2351) & (x0 | (x1 ? (x3 | ~n1846) : (~x3 | n2351)));
  assign n2351 = (~x4 | ~x5 | x6 | x7) & (x4 | x5 | ~x6 | ~x7);
  assign n2352 = x2 ? (n2353 & n2358) : n2357;
  assign n2353 = (x1 | n2355) & (x0 | ~x1 | (~n2356 & (n2354 | n1307)));
  assign n2354 = ~x3 ^ ~x5;
  assign n2355 = (((x0 | x4 | ~x5 | ~x6) & (~x0 | ~x4 | x5 | x6)) | (x3 ^ ~x7)) & (x5 | ~x6 | x7 | ~x0 | ~x3 | x4) & ((x4 ? (~x6 | ~x7) : (x6 | x7)) | (x0 ? (x3 | ~x5) : (~x3 | x5)));
  assign n2356 = x7 & ~x6 & x5 & ~x3 & ~x4;
  assign n2357 = (~x1 | ((x0 | (x4 ? (x3 ? (x5 ^ x6) : (~x5 | x6)) : (x5 | ~x6))) & (x3 | ((~x4 | x5 | ~x6) & (~x5 | x6 | ~x0 | x4))))) & (~x0 | ~x3 | x4 | x5 | x6) & (x1 | ((~x3 | ((~x5 | x6 | ~x0 | ~x4) & (x0 | (x4 ? (x5 | ~x6) : (~x5 | x6))))) & (x3 | ~x5 | ~x6) & (~x0 | x4 | (x5 ^ x6))));
  assign n2358 = (x1 | (x5 ? ((x0 | (x3 ? x6 : (~x4 | ~x6))) & (~x3 | (x6 ? ~x0 : ~x4))) : ((~x0 | (x3 ? (x4 | x6) : ~x6)) & (x3 | (x6 ? x4 : x0))))) & (x0 | ~x1 | (x3 ? (x5 | (~x4 & ~x6)) : (~x5 | (~x4 ^ x6))));
  assign z164 = ~n2365 | (x2 ? ~n2360 : (x4 ? ~n2363 : ~n2364));
  assign n2360 = x0 ? (x1 | n2362) : n2361;
  assign n2361 = x1 ? ((x3 | x4 | ~x5 | ~x6 | x7) & (~x3 | ((x6 | ~x7 | x4 | x5) & (~x4 | ~x6 | (~x5 ^ x7))))) : (x3 ? (~x4 | x7 | (~x5 ^ x6)) : (x4 | (x5 ? (x6 | ~x7) : ~x6)));
  assign n2362 = (~x5 | x6 | ~x3 | x4) & (~x6 | ((x3 | ~x4 | x5 | x7) & (~x3 | (x4 ? (~x5 | ~x7) : (x5 | x7)))));
  assign n2363 = x3 ? ((x1 | (x0 ? (~x6 | (~x5 ^ x7)) : (x5 | x6))) & (x0 | ~x1 | x7 | (~x5 ^ x6))) : ((x0 | x1 | ~x5 | ~x6 | x7) & (~x0 | ~x1 | x5 | x6 | ~x7));
  assign n2364 = (~x5 | ~x6 | x7 | x0 | x1 | ~x3) & (x3 | x6 | (x0 ? (~x1 | ~x7) : (x1 ? (~x5 | x7) : (x5 | ~x7))));
  assign n2365 = (~x1 | n2368) & (n662 | n2366) & (x1 | n2367);
  assign n2366 = x4 ? (x5 ? ((~x1 | x2 | x3) & (x0 | x1 | (x2 & x3))) : ((x1 | x2 | x3) & (~x0 | (x2 ? x1 : x3)))) : (x0 ? (x1 | (x3 ? x2 : ~x5)) : ((~x2 | ~x3 | x5) & (~x1 | (~x2 & x5))));
  assign n2367 = x0 ? ((x6 | ~x7 | x4 | x5) & (~x4 | ((~x6 | x7 | ~x2 | ~x5) & (x2 | (x5 ? (x6 | ~x7) : (~x6 | x7)))))) : (x2 ? ((x4 | ~x5 | ~x6 | x7) & (~x4 | x6 | ~x7)) : (x4 | (x5 ? (x6 | ~x7) : (~x6 | x7))));
  assign n2368 = (x2 | ((x5 | ~x6 | x7 | ~x0 | x4) & (x0 | ((x4 | ~x5 | ~x6 | x7) & (~x4 | x6 | ~x7))))) & (x0 | ~x4 | ((~x2 | x5 | ~x6 | x7) & (~x5 | x6 | ~x7)));
  assign z165 = n2370 | n2373 | (~n2181 & ~n2377) | (~n662 & ~n2376);
  assign n2370 = ~x0 & (x6 ? ~n2371 : ~n2372);
  assign n2371 = (x5 | ((~x3 | (x1 ? (x2 ? (~x4 | ~x7) : x7) : (x2 ? x7 : (~x4 | ~x7)))) & (x4 | ((~x1 | x2 | x7) & (x3 | ~x7 | x1 | ~x2))))) & (~x3 | ~x5 | (x1 ? (x2 ? x7 : (~x4 | ~x7)) : (x2 ? (~x4 | ~x7) : x7)));
  assign n2372 = (~x4 | ((x5 | ((x1 | ~x2 | ~x3 | x7) & (~x1 | ((x3 | ~x7) & (x2 | ~x3 | x7))))) & (x1 | ~x5 | (x2 ? (x3 | ~x7) : (~x3 | x7))))) & (~x2 | ((x1 | x3 | x4 | x5 | ~x7) & (~x1 | ~x3 | ~x5 | x7))) & (~x5 | ((x2 | x3 | x4 | ~x7) & (~x1 | ((x3 | x4 | ~x7) & (x2 | ((x4 | ~x7) & (x3 | (x4 & ~x7))))))));
  assign n2373 = x0 & ((n538 & ~n2375) | (~x2 & ~n2374));
  assign n2374 = (~x4 | ((x5 | ~x7 | x1 | ~x3) & (x3 | ((~x6 | ~x7 | x1 | ~x5) & (~x1 | ((~x6 | x7) & (x5 | x6 | ~x7))))))) & (x1 | ((~x3 | ~x5 | x7) & (x4 | (x5 ? (~x6 | x7) : (x6 | ~x7)))));
  assign n2375 = (~x4 | ((~x5 | x6 | ~x7) & (~x3 | x5 | x7))) & (~x3 | ~x6 | (x5 ^ x7)) & (x3 | x4 | x5 | x6 | ~x7);
  assign n2376 = (x3 | ((~x0 | (x1 ? (x2 | ~x5) : x5)) & (~x4 | x5 | x1 | ~x2) & (x0 | (x1 ? (x2 ? ~x5 : (~x4 | x5)) : (x2 | ~x5))))) & (x4 | ((~x3 | x5 | x1 | ~x2) & (x0 | x2 | (x1 ? (~x3 | x5) : ~x5))));
  assign n2377 = (x4 | ((~x0 | ~x1 | x2 | x5) & (x1 | ~x2 | ~x5))) & (x0 | (x1 ? (x2 ? x5 : (~x4 | ~x5)) : (x2 ^ x5)));
  assign z166 = ~n2381 | (~x2 & ((~x7 & ~n2379) | (x0 & x7 & ~n2380)));
  assign n2379 = (x1 | ((x0 | x3 | x4 | x5 | ~x6) & (~x0 | ~x4 | (x3 ? ~x6 : (~x5 | x6))))) & (x0 | ~x1 | x5 | (x3 ? (~x4 | ~x6) : (x4 | x6)));
  assign n2380 = (~x1 | x3 | x4 | ~x5 | x6) & (x1 | ((~x5 | x6 | x3 | ~x4) & (~x3 | ~x6 | (~x4 & ~x5))));
  assign n2381 = ~n2382 & (n620 | n2386) & (x4 ? n2385 : n2387);
  assign n2382 = x2 & ((~x4 & ~n2383 & ~x0 & x1) | (~x1 & (~n2384 | (x0 & ~n2383))));
  assign n2383 = (x3 | x5 | x6 | x7) & (~x3 | ~x5 | ~x6 | ~x7);
  assign n2384 = (x0 | ~x3 | ~x4 | ~x5 | ~x6 | x7) & (~x0 | ((~x6 | ((x3 | x4 | x5 | ~x7) & (~x3 | (x4 ? x5 : (~x5 | x7))))) & (x3 | x6 | ((~x5 | x7) & (~x4 | x5 | ~x7)))));
  assign n2385 = (x0 | ((~x2 | (x3 ? (x5 | ~x6) : x6)) & (x3 | ~x5 | x6) & (~x3 | ~x6 | (~x7 & (x2 | ~x5))))) & (x2 | x3 | x5 | x6 | (~x0 & x7));
  assign n2386 = (~x0 | x3 | ~x4 | ~x5 | (x1 ^ ~x2)) & (~x3 | ((x0 | (x4 & (x1 | x2 | x5))) & (x4 | ((x2 | x5) & (x1 | (x2 & x5))))));
  assign n2387 = (x2 | ((x0 | ~x3 | x5 | x6 | x7) & (x3 | ((x5 | ~x6 | ~x7) & (~x0 | x6 | x7))))) & (x0 | x3 | ((~x6 | ~x7) & (~x5 | x6 | x7)));
  assign z167 = ~n2391 | (~x0 & (x3 ? ~n2389 : ~n2390));
  assign n2389 = x6 ? ((~x1 | ~x2 | ~x5 | (~x4 ^ x7)) & (x2 | x5 | ((x4 | x7) & (x1 | ~x4 | ~x7)))) : ((~x5 | ~x7 | ~x2 | ~x4) & (x2 | x5 | ((~x4 | x7) & (x1 | x4 | ~x7))));
  assign n2390 = (~x4 | ((~x6 | ~x7 | x2 | x5) & (x6 | ((x1 | ~x2 | x5 | x7) & (~x1 | (x2 ? (~x5 | ~x7) : (x5 | x7))))))) & (x1 | x4 | x5 | (x2 ? (~x6 | x7) : (x6 | ~x7)));
  assign n2391 = (~n2392 | n2395) & (x2 | n2394) & (~x2 | n2393);
  assign n2392 = x5 & x0 & ~x1;
  assign n2393 = (x1 | (x4 ? (~x7 | (x5 & (x0 | x3))) : ((~x3 | x5 | x7) & (~x0 | ((x5 | x7) & (~x3 | ~x5 | ~x7)))))) & (x0 | (x4 ? (x5 | ~x7) : (x7 | (~x1 & ~x5))));
  assign n2394 = (~x3 | ((~x5 | x7 | x1 | x4) & (~x4 | ~x7 | x0 | ~x1))) & (~x4 | ((x0 | ((~x5 | ~x7) & (x1 | x3 | x5 | x7))) & (~x7 | ((x1 | x3 | ~x5) & (~x0 | x5 | (x1 & x3)))) & (~x0 | ~x1 | x3 | ~x5 | x7))) & (x4 | ((~x0 | ((x5 | x7) & (~x1 | x3 | ~x5 | ~x7))) & (x7 | ((x0 | ~x5) & (~x1 | x3 | x5)))));
  assign n2395 = x7 ? ((x2 | ((x4 | ~x6) & (~x3 | ~x4 | x6))) & (x3 | ((x4 | ~x6) & (~x2 | ~x4 | x6)))) : ((x3 | x4 | x6) & (~x2 | (~x4 ^ ~x6)));
  assign z168 = n2398 | ~n2399 | n2400 | n2404 | (~x0 & ~n2397);
  assign n2397 = (x1 | ((x2 | ~x5 | x6) & (~x2 | x3 | x5 | ~x6))) & (x5 | ~x6 | x2 | ~x3) & (~x1 | ((~x4 | ~x5 | ~x6 | ~x2 | ~x3) & (x5 | ((x2 | ~x4 | ~x6) & (x6 | (x2 ^ (x3 | x4)))))));
  assign n2398 = n738 & (x5 ? (x6 & (x2 | (~x3 & ~x4))) : (~x6 & ((x2 & (~x3 | ~x4)) | (~x3 & ~x4) | (~x2 & x3 & x4))));
  assign n2399 = x0 ? (x2 | ((~x1 | x3 | ~x5) & (x4 | x5 | x1 | ~x3))) : (~x2 | x5 | (x1 ? (x3 | x4) : ~x3));
  assign n2400 = ~x1 & (n2401 | n2402 | (~x0 & n871 & n587));
  assign n2401 = ~n1116 & (x0 ? (x3 & ((x4 & ~x5 & ~x7) | (x5 & x7))) : (~x3 & (x5 ^ x7)));
  assign n2402 = n610 & n691 & (n2403 | (x2 & n2237));
  assign n2403 = ~x6 & ~x2 & x4;
  assign n2404 = x1 & ((n559 & n1415) | (~x0 & ~n2405));
  assign n2405 = ((x3 ^ ~x4) | ((x6 | x7 | x2 | ~x5) & (~x2 | ~x6 | (x5 ^ x7)))) & (x2 | x5 | ((~x3 | x6 | ~x7) & (x3 | x4 | ~x6 | x7)));
  assign z169 = n2407 | n2410 | n2412 | ~n2413 | (~n620 & ~n2409);
  assign n2407 = ~x0 & ((n1386 & n837) | (x4 & ~n2408));
  assign n2408 = (~x5 | ~x6 | x7 | x1 | x2 | ~x3) & (~x2 | ((~x5 | x6 | ~x7 | x1 | x3) & (~x1 | x5 | (x3 ? (x6 | x7) : (~x6 | ~x7)))));
  assign n2409 = (~x5 | ((~x0 | x1 | ~x2 | ~x3) & (x0 | ~x1 | x2 | x3 | ~x4))) & (x1 | (x0 ? (~x4 | (x2 ? ~x3 : (x3 | x5))) : (~x2 | x3 | (x4 & x5)))) & (~x1 | x2 | ((x4 | x5 | ~x0 | x3) & (x0 | ~x3 | (x4 & x5))));
  assign n2410 = ~n662 & ~n2411;
  assign n2411 = (x1 | (x0 ? ((x2 | ~x3 | ~x4) & (x4 | x5 | ~x2 | x3)) : (~x4 | (x2 ? (~x3 | ~x5) : x3)))) & (x0 | ((x4 | ~x5 | x2 | x3) & (~x1 | (x2 ? (x3 ? x4 : (~x4 | ~x5)) : (x3 | x4)))));
  assign n2412 = x0 & ((~x1 & ~x2 & x3 & ~x4 & ~x6) | (~x3 & ((x1 & ~x2 & x4 & ~x6) | (~x1 & x6 & (~x2 ^ x4)))));
  assign n2413 = ~n2414 & ~n2415 & ~n2416 & (~n541 | n1115 | n1117);
  assign n2414 = ~x0 & ((~x1 & ~x2 & x3 & ~x4 & x6) | (x2 & ((x1 & (x3 ? (x4 & x6) : (~x4 & ~x6))) | (~x4 & ~x6 & ~x1 & x3))));
  assign n2415 = n2392 & (x2 ? (~x3 & n672) : (x7 & ~n571));
  assign n2416 = n545 & ((~n1116 & n2417) | (x3 & n1121 & n539));
  assign n2417 = ~x5 & (~x1 ^ ~x3);
  assign z170 = ~n2421 | (~x0 & (n2420 | (x1 & ~n2419)));
  assign n2419 = (x6 | ((~x2 | x3 | ~x4 | x5 | x7) & (x2 | ~x7 | (x3 ? (~x4 | x5) : (x4 | ~x5))))) & (~x2 | ~x4 | x5 | ~x6 | (x3 ^ ~x7));
  assign n2420 = x5 & n648 & ((x3 & (x2 ? (~x6 & ~x7) : (x6 & x7))) | (x2 & ~x3 & (x6 ^ x7)));
  assign n2421 = ~n2422 & n2424 & ~n2425 & (x0 ? n2423 : n2426);
  assign n2422 = n2392 & ((x6 & ((x2 & ~x3 & ~x4 & ~x7) | (~x2 & (x3 ? (~x4 & x7) : (x4 & ~x7))))) | (x2 & ~x4 & ~x6 & (x3 ^ x7)));
  assign n2423 = (x1 | x2 | x3 | ~x4 | x5 | ~x7) & (x4 | (x5 ? ((x1 | ~x2 | ~x3 | ~x7) & (x3 | x7 | ~x1 | x2)) : ((x1 ^ ~x2) | (~x3 ^ x7))));
  assign n2424 = (x3 | ~x4 | x7 | ~x0 | ~x1 | x2) & (((~x3 | ~x7) & (~x2 | x3 | x7)) | (x0 ? (x1 | ~x4) : (~x1 | x4)));
  assign n2425 = ~x1 & ((~x4 & ~x7 & x0 & ~x2) | (~x0 & (~x2 | ~x4) & (x3 ^ x7)));
  assign n2426 = x1 ? ((~x5 | x7 | ~x3 | ~x4) & (x3 | ((~x4 | ~x5 | ~x7) & (x2 | x5 | (~x4 ^ x7))))) : (~x2 | ~x4 | (x3 ? (x5 ^ x7) : (x5 | ~x7)));
  assign z171 = n2431 | n2432 | ~n2433 | (~x0 & (~n2428 | ~n2430));
  assign n2428 = (x4 | n2429) & (~x7 | n1116 | n1243 | ~x3 | ~x4);
  assign n2429 = (x1 | x2 | x3 | x5 | x6 | ~x7) & (x7 | ((~x1 | ~x2 | x3 | x5 | ~x6) & (x1 | ~x3 | ~x5 | (~x2 ^ x6))));
  assign n2430 = (~x2 | (x1 ? (x5 | (x4 ^ x6)) : (~x5 | ((~x4 | ~x6) & (x3 | x4 | x6))))) & (x1 | x2 | x4 | (x3 ? (~x5 | x6) : (x5 | ~x6)));
  assign n2431 = ~x2 & ((~x1 & ((~x0 & ~x4 & (x3 ^ x5)) | (x4 & x5 & x0 & ~x3))) | (x0 & x1 & ~x3 & (x4 ^ x5)));
  assign n2432 = n738 & ((n1902 & n1956) | (n985 & ~n592 & ~n1116));
  assign n2433 = n2434 & (~n2392 | ((~x4 | x6 | x2 | ~x3) & (~x2 | ((x4 | ~x6) & (x3 | ~x4 | x6)))));
  assign n2434 = (x0 | ((x4 | x5 | x1 | ~x2) & (~x1 | ((~x4 | ~x5) & (x2 | x4 | x5))))) & (~x4 | x5 | ~x0 | x1);
  assign z172 = n2436 | ~n2440 | (~x5 & ~n2439) | (~x1 & ~n2438);
  assign n2436 = ~x0 & (x1 ? ~n2437 : (n665 & n686));
  assign n2437 = (~x2 | x3 | x4 | x5 | ~x6 | ~x7) & (~x3 | (~x2 ^ x6) | ((~x5 | x7) & (~x4 | x5 | ~x7)));
  assign n2438 = (x5 | ((x2 | x3 | x4 | x6 | ~x7) & (x7 | ((x2 | ~x3 | ~x4 | ~x6) & (~x2 | (x3 ? (~x4 | x6) : (x4 | ~x6))))))) & (~x3 | ~x5 | ~x7 | (~x2 ^ x6));
  assign n2439 = (~x2 | ((x0 | ~x1 | x3 | ~x4 | ~x6) & (x4 | x6 | x1 | ~x3))) & (x1 | x2 | ((x3 | ~x4 | x6) & (x4 | ~x6 | ~x0 | ~x3)));
  assign n2440 = n2441 & (~n664 | ((~x5 | x6 | x2 | ~x3) & (~x2 | (x3 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n2441 = (x2 | ((x5 | x6 | x1 | ~x3) & (x3 | (x1 ? (~x5 & ~n559) : (x5 | ~x6))))) & (x1 | ~x2 | ((~x5 | ~x6) & (x3 | x5 | x6)));
  assign z173 = n2444 | n2446 | n2447 | ~n2448 | (~n620 & ~n2443);
  assign n2443 = x2 ? (~x3 | (~x4 & ~x5) | (x0 & x1)) : (x3 | x4 | x5 | (~x0 & x1));
  assign n2444 = ~x4 & ((n1558 & ~n2445) | (n708 & n540 & n1176));
  assign n2445 = (~x6 | x7 | ~x2 | ~x3) & (x2 | ~x7 | (x1 ? (x3 | x6) : (~x3 | ~x6)));
  assign n2446 = ~n662 & ~n1799 & ((x2 & ~x3 & ~x4 & ~x5) | (~x2 & x3 & (x4 | x5)));
  assign n2447 = x2 & x6 & n738 & (~x3 ^ (~x4 & ~x5));
  assign n2448 = (x2 | ~x3 | x4 | x5 | x6) & (x3 | (~x4 & ~x5) | ((x2 | x6) & (x0 | ~x2 | ~x6)));
  assign z174 = n2452 | (~x4 & (n2451 | ~n2453 | (~x1 & ~n2450)));
  assign n2450 = x6 ? ((x5 | ~x7 | x0 | ~x3) & (~x0 | ~x2 | x3 | ~x5 | x7)) : (x0 ? (x2 | (x3 ? (~x5 | x7) : (x5 | ~x7))) : (~x2 | x5 | (~x3 ^ x7)));
  assign n2451 = n1843 & (x2 ? (x3 & n537) : (~x3 & ~n620));
  assign n2452 = x4 & ((~x2 & ~x3 & ~x7) | ((~x0 | ~x1) & (~x3 ^ x7)));
  assign n2453 = (~x5 & ((~x0 & (x1 ? (~x2 & x7) : x2)) | (~x3 & ~x7) | (x7 & (x3 | (x0 & ~x1 & ~x2))))) | (x5 & (x3 ^ x7)) | (x0 & ((x2 & x5 & ~x7) | (x1 & (x2 | (x5 & x7)))));
  assign z175 = n2455 | n2457 | ~n2458 | ~n2459 | (n605 & ~n2456);
  assign n2455 = ~x1 & ((x0 & x4 & ~x5 & (x2 ^ x3)) | (~x4 & x5 & (~x0 | (~x2 & ~x3))));
  assign n2456 = (~x5 | x6 | ~x7 | ~x0 | x2 | ~x4) & (x0 | x5 | ~x6 | (x2 ? (x4 | ~x7) : (~x4 | x7)));
  assign n2457 = (x4 ^ x5) & ((x0 & ~x1 & x2 & x3) | (x1 & ((~x2 & ~x3) | (~x0 & (~x2 | ~x3)))));
  assign n2458 = ~n1449 | ((x0 | ~x1 | ~x2 | ~x3) & (~x0 | x1 | ~x6 | (~x2 ^ x3)));
  assign n2459 = (x5 | n2460) & (n592 | n2461);
  assign n2460 = (x1 | x2 | x3 | ~x4 | x6) & (x0 | ((~x4 | x6 | ~x2 | ~x3) & (~x1 | x2 | x3 | x4 | ~x6) & (x1 | ((~x4 | x6) & (x4 | ~x6 | ~x2 | ~x3)))));
  assign n2461 = (~x3 | ((~x0 | x1 | x2 | ~x5 | x6) & (x0 | x5 | ~x6 | (~x1 ^ ~x2)))) & (~x0 | x1 | x3 | (x2 ? (~x5 | x6) : (x5 | ~x6)));
  assign z176 = n2464 | ~n2466 | ~n2469 | (n708 & ~n2463);
  assign n2463 = (x4 | ~x6 | ~x7 | x0 | ~x1 | ~x2) & (x2 | ((x0 | ~x1 | ~x4 | ~x6 | x7) & (~x0 | x1 | ~x7 | (~x4 ^ ~x6))));
  assign n2464 = ~n2465 & ((~x1 & ((x0 & (x5 ? x6 : (~x6 & ~x7))) | (x7 & ((x5 & ~x6) | (~x0 & ~x5 & x6))))) | (~x0 & x5 & (~x6 | (x1 & ~x7))));
  assign n2465 = x2 ^ ~x3;
  assign n2466 = ~n2468 & (~n708 | ~n534 | ~n540) & (~n2467 | ~n1546);
  assign n2467 = x6 & x3 & ~x5;
  assign n2468 = x5 & (x0 ? (x1 ? (~x2 & ~x3) : (x2 & x3)) : (~x6 & (x2 ^ ~x3)));
  assign n2469 = (~x6 | n2470) & (x5 | (~n2471 & ~n2472));
  assign n2470 = (x0 | ((x1 | x2 | ~x5 | x7) & (~x1 | (x2 ? (~x3 | (~x5 ^ x7)) : (~x5 | ~x7))))) & (x1 | x2 | x3 | ((~x5 | x7) & (~x0 | x5 | ~x7)));
  assign n2471 = ~x1 & ~n607 & ((n669 & n642) | (n732 & n641));
  assign n2472 = n2473 & (n2237 | n838);
  assign n2473 = ~x3 & ~x2 & ~x0 & x1;
  assign z177 = n2475 | ~n2480 | n2482 | n2483 | (~x1 & ~n2479);
  assign n2475 = x7 & ((n2476 & n2477) | (n1148 & ~n2478));
  assign n2476 = x4 & (x5 ^ ~x6);
  assign n2477 = ~x3 & x2 & ~x0 & x1;
  assign n2478 = (x0 | x1 | x3 | x5 | x6) & ((~x1 ^ x5) | (x0 ? (~x3 | x6) : (x3 | ~x6)));
  assign n2479 = (x0 | ~x2 | x3 | x4 | x6 | x7) & (~x4 | (((x2 ^ ~x7) | (x0 ? (~x3 | x6) : (x3 | ~x6))) & (x0 | x2 | x3 | x6 | x7)));
  assign n2480 = n2481 & (~n2328 | ((x6 | ~x7 | ~x2 | x4) & (x2 | (x4 ? (x6 | ~x7) : (~x6 | x7)))));
  assign n2481 = (~x3 | ((~x0 | x1 | x2 | ~x6 | x7) & (x0 | (x6 ? ((x1 | (~x2 & ~x7)) & (~x2 | ~x7)) : ((x2 | x7) & (~x1 | (x2 & x7))))))) & (~x0 | x2 | x3 | ((x1 | ~x6 | ~x7) & (x6 | (~x1 & x7))));
  assign n2482 = x2 & ((~x0 & x1 & ~x3 & ~x6 & ~x7) | (~x1 & ((x6 & x7 & ~x0 & ~x3) | (x0 & ((~x6 & x7) | (~x3 & x6 & ~x7))))));
  assign n2483 = ~x7 & (~n2484 | (~x2 & (n2117 | (n983 & n958))));
  assign n2484 = (~n1546 | ~n1179) & (n912 | n2485);
  assign n2485 = (x0 | ~x1 | x2 | x3 | ~x4) & (~x0 | x1 | ~x2 | ~x3 | x4);
  assign z178 = n2487 | n2491 | ~n2492 | (~x1 & ~n2490);
  assign n2487 = ~x2 & ((~x3 & ~n2489) | (x3 & ~x4 & n738 & n2488));
  assign n2488 = ~x5 & (x6 ^ ~x7);
  assign n2489 = (~x0 | x1 | ~x4 | ~x5 | ~x6 | x7) & (x0 | (x1 ? (~x7 | (x4 ? (x5 | x6) : (~x5 | ~x6))) : (x4 | x7 | (~x5 ^ x6))));
  assign n2490 = (~x4 | x5 | ~x7 | ~x0 | x2 | x3) & (x4 | ((x0 | ~x2 | x3 | x5 | ~x7) & (~x5 | ((x3 | ~x7 | x0 | x2) & (~x0 | ~x3 | (x2 ^ ~x7))))));
  assign n2491 = ~x3 & ((~x4 & ~x7 & ~x0 & x1) | (~x1 & ((~x0 & x4 & (x2 ^ x7)) | (~x4 & x7 & x0 & ~x2))));
  assign n2492 = n2495 & (~x1 | n2494) & (x1 | ~x2 | x4 | n2493);
  assign n2493 = (~x0 | ~x3 | x5 | x6 | ~x7) & (x0 | x3 | ~x5 | (~x6 ^ x7));
  assign n2494 = (x0 | x3 | ~x4 | (x2 ? (x5 ^ x7) : (~x5 | x7))) & (~x0 | x2 | ~x3 | x4 | x5 | x7);
  assign n2495 = (~x0 | x3 | (x1 ? (x2 | x7) : (~x2 | ~x7))) & (~x3 | ((x1 | ~x4 | (~x2 ^ x7)) & (x0 | (x1 ? (~x2 ^ ~x7) : (~x2 ^ x7)))));
  assign z179 = n2499 | ~n2501 | n2505 | (x4 ? ~n2504 : ~n2497);
  assign n2497 = (x2 | ~n598 | ~n618) & (~x6 | ~n2127 | n2498);
  assign n2498 = (~x1 | x2 | x3 | x7) & (x1 | ~x2 | ~x3 | ~x7);
  assign n2499 = ~n910 & (x0 ? (~x3 & n965) : (~n2500 | n635));
  assign n2500 = x3 ? (x4 | x5) : (~x4 | ~x5);
  assign n2501 = ~n2502 & (~n650 | (x0 ? (x1 | ~x5) : (x1 ? ~x2 : (x2 | x5))));
  assign n2502 = x4 & n664 & ((n871 & n2155) | (n563 & n2503));
  assign n2503 = x7 & ~x5 & x6;
  assign n2504 = x0 ? (x1 | ~x3) : (x1 ? ((~x3 | x5) & (~x2 | x3 | ~x5)) : (x3 | (x2 & x5)));
  assign n2505 = n2237 & ((x0 & ~x1 & ~x2 & x3 & ~x5) | (~x0 & x5 & (x1 ? (~x2 & x3) : ~x3)));
  assign z180 = ~n2515 | n2513 | n2511 | ~n2510 | n2507 | n2509;
  assign n2507 = ~x0 & ((x4 & ~n2508) | (~x1 & n665 & n1231));
  assign n2508 = (x1 | ~x2 | ~x3 | ~x5 | ~x6 | x7) & (~x1 | ~x7 | ((x2 | x3 | x5 | ~x6) & (~x5 | x6 | ~x2 | ~x3)));
  assign n2509 = x1 & ((x0 & ~x2 & ~x3 & ~x4 & x5) | (~x0 & ((~x2 & x3 & ~x4 & ~x5) | (x4 & x5 & x2 & ~x3))));
  assign n2510 = x2 | x4 | ~n738 | (x5 ? (~x3 & ~n540) : x3);
  assign n2511 = x6 & n2512 & (x0 ? (~x5 & ~n2465) : (x5 & (~n2465 | ~n1809)));
  assign n2512 = ~x1 & ~x4;
  assign n2513 = ~n592 & ((n2514 & n677) | (x6 & n2127 & ~n2156));
  assign n2514 = ~x6 & ~x3 & x5;
  assign n2515 = n2516 & (~x4 | n2517);
  assign n2516 = (~x0 | x1 | ~x2 | x4 | ~x5) & (x0 | (x1 ? (x2 ? (x4 | x5) : (~x4 | ~x5)) : (~x4 | x5)));
  assign n2517 = x1 ? ((x3 | x5 | x6 | ~x0 | x2) & (~x3 | ~x5 | ~x6 | x0 | ~x2)) : (x6 | (~x2 & ~x3) | (~x0 ^ x5));
  assign z181 = ~n2521 | (~x2 & (n2520 | (~x0 & ~n2519)));
  assign n2519 = (x6 | ((x3 | ((x5 | x7 | x1 | ~x4) & (~x1 | (~x4 ^ ~x5)))) & (x1 | ~x3 | ~x7 | (~x4 ^ x5)))) & (~x1 | x3 | (x4 ? (x5 ? x7 : (~x6 | ~x7)) : (x5 | x7)));
  assign n2520 = ~x3 & ~x4 & x5 & n738 & (x6 | n543);
  assign n2521 = ~n2523 & n2524 & ~n2526 & (x0 ? n2525 : n2522);
  assign n2522 = (x1 | x2 | x3 | ~x5 | x6 | ~x7) & (~x3 | ((x1 | ((x6 | x7 | x2 | x5) & (~x6 | ~x7 | ~x2 | ~x5))) & (~x5 | x6 | ~x7 | ~x1 | ~x2)));
  assign n2523 = (~x0 | (~x1 & (~x5 | ~x6))) & (x0 | (x5 & (x1 | x6))) & (x5 | x6) & (x2 | x3) & (~x2 | ~x3);
  assign n2524 = (x0 | x1 | ~x2 | x5 | x6) & (~x5 | (x0 ? (x6 | (x1 ? (x2 | x3) : (~x2 | ~x3))) : (~x6 | (x1 ? (~x2 | ~x3) : (x2 | x3)))));
  assign n2525 = (x1 | x2 | x3 | x5 | x6 | x7) & (~x6 | (x1 ? (x2 | x3) : (~x2 | ~x3)) | (~x5 ^ x7));
  assign n2526 = n616 & n2527 & ((~x1 & ~x4 & x5 & x6) | (x1 & ~x6 & (~x4 ^ ~x5)));
  assign n2527 = x3 & ~x7;
  assign z182 = n2529 | n2531 | ~n2532 | n2535 | (~n662 & ~n2534);
  assign n2529 = x3 & ((~x4 & ~n2530) | (x2 & n2135 & n598));
  assign n2530 = x0 ? (x5 | ((~x6 | ~x7 | x1 | ~x2) & (~x1 | x2 | x6 | x7))) : (~x1 | ~x5 | (x2 ? (~x6 | x7) : (x6 | ~x7)));
  assign n2531 = ~x1 & x6 & ((x2 & ~x3) | (x0 & ~x2 & x3));
  assign n2532 = n2533 & (~n587 | ~n1476) & (n1446 | ~n1317 | n599);
  assign n2533 = x0 | ~x1 | (x2 ? ~n1136 : ~n2288);
  assign n2534 = x1 ? (x2 | x3) : (~x2 | ~x3 | ((~x4 | ~x5) & (~x0 | (~x4 & ~x5))));
  assign n2535 = ~n620 & ((~x1 & ~x2 & ~x3) | (~x0 & ((x1 & x2 & x3 & x4) | (~x1 & ~x2 & ~x4))));
  assign z183 = n2537 | ~n2540 | (n1317 & (~n2539 | ~n2543 | ~n2544));
  assign n2537 = x0 & ((~x6 & ~n2538) | (n1386 & n943));
  assign n2538 = (~x1 | x2 | ~x3 | x4 | x5 | ~x7) & (x1 | ((x2 | x3 | ~x4 | ~x5 | ~x7) & (~x2 | ~x3 | x4 | x5 | x7)));
  assign n2539 = (x1 | x4 | (~x2 ^ x7)) & (~x4 | ((~x1 | ~x2 | ~x7) & (x2 | x7)));
  assign n2540 = (x1 | ((~x2 | x3 | x7) & (~x0 | ~x3 | (x2 ^ x7)))) & n2541 & (x3 | ((~x1 | x2 | ~x7) & (x0 | (~x2 ^ x7))));
  assign n2541 = ~n534 | (~n2542 & ~n1979);
  assign n2542 = x7 & ~x3 & ~x4;
  assign n2543 = (~x4 | ~x5 | ~x7 | x1 | ~x2) & (x7 | ((~x4 | x5 | x1 | ~x2) & (~x1 | x4 | (~x2 ^ x5))));
  assign n2544 = (x5 | ~x6 | ~x7 | x1 | ~x2 | ~x4) & (~x1 | x4 | ((x6 | ~x7 | x2 | x5) & (~x2 | ~x5 | (x6 ^ x7))));
  assign z184 = n2546 | n2549 | ~n2551 | ~n2555 | (n1122 & ~n2548);
  assign n2546 = ~x7 & ((~x2 & n1543 & n1838) | (~x4 & ~n2547));
  assign n2547 = (~x1 | x2 | ~x3 | x5 | ~x6) & (~x2 | ((x0 | ~x5 | ~x6 | (~x1 ^ x3)) & (~x0 | x1 | ~x3 | x5 | x6)));
  assign n2548 = (x1 | x2 | x4 | ~x5 | ~x6) & (x0 | ((~x5 | ~x6 | x2 | x4) & (~x4 | x5 | ~x1 | ~x2)));
  assign n2549 = ~n2550 & (x1 ? ~x3 : (x3 & x6));
  assign n2550 = (x0 | ~x2 | (x4 ? (x5 | x7) : (~x5 | ~x7))) & (~x4 | ~x5 | ~x7 | ~x0 | x2);
  assign n2551 = ~n2552 & ~n2553 & n2554 & (x3 | ~n2095 | ~n651);
  assign n2552 = ~x0 & ((~x3 & x4 & (~x2 | x5)) | (~x4 & ~x5 & x2 & x3));
  assign n2553 = ~x0 & x3 & ~x4 & ~x6 & (~x2 ^ x5);
  assign n2554 = ~x0 | x1 | ~n923 | (~x2 & ~n1121);
  assign n2555 = ~n2557 & (x5 | ((~n1590 | ~n677) & (n1323 | n2556)));
  assign n2556 = (~x0 | ~x1 | x2 | x4) & (x0 | x1 | ~x2 | ~x4);
  assign n2557 = ~x4 & ((~x0 & ~x1 & ~x2 & x3 & x5) | (x0 & ~x3 & (x1 ? (~x2 & x5) : x2)));
  assign z185 = n2562 | ~n2563 | (x2 ? ~n2567 : (~n2559 | ~n2568));
  assign n2559 = x3 ? (~x6 | n2561) : n2560;
  assign n2560 = x4 ? (~x7 | ((~x1 | x5 | ~x6) & (~x5 | x6 | ~x0 | x1))) : ((x1 | ~x5 | ~x6 | x7) & (x0 | ((~x5 | ~x6 | x7) & (x6 | ~x7 | x1 | x5))));
  assign n2561 = (~x1 | x4 | x5 | x7) & (~x0 | x1 | ~x5 | (~x4 ^ x7));
  assign n2562 = ~x1 & ((x0 & x2 & ~x3 & x4 & ~x5) | (~x2 & (x0 ? (~x5 & (x3 ^ ~x4)) : (x3 & ~x4))));
  assign n2563 = n2566 & (~x2 | (x6 ? (~n1317 | n2565) : n2564));
  assign n2564 = (x0 | x1 | x3 | x4 | x5 | ~x7) & ((x4 ^ x7) | ((~x0 | x1 | ~x3 | x5) & (x0 | ~x1 | x3 | ~x5)));
  assign n2565 = (~x1 | ~x4 | ~x5 | ~x7) & (x1 | x5 | (~x4 ^ x7));
  assign n2566 = (x0 | ~x1 | ~x2 | x4 | x5) & (~x5 | ((x0 | (x1 ? (x2 | ~x4) : (~x2 | x4))) & (~x4 | ((~x0 | x1 | ~x2) & (~x1 | x2 | x3)))));
  assign n2567 = (~x4 | x5 | ~x6 | ~x0 | x1 | ~x3) & (x0 | (x1 ? (~x5 | (x3 ? (x4 | x6) : (~x4 | ~x6))) : (x5 | ((x3 | x4 | ~x6) & (~x4 | x6)))));
  assign n2568 = (x0 | x1 | x3 | x4 | x5 | ~x6) & (x6 | ((~x0 | ((~x1 | x4 | x5) & (x1 | ~x3 | ~x4 | ~x5))) & (x4 | ((~x1 | ~x3 | x5) & (x3 | ~x5 | (x0 & x1))))));
  assign z186 = n2570 | n2572 | ~n2578 | (x2 ? ~n2577 : ~n2576);
  assign n2570 = x1 & ((n2314 & n686) | (~x0 & ~n2571));
  assign n2571 = (~x6 | ((x2 | x4 | (x3 ? (x5 | x7) : (~x5 | ~x7))) & (~x4 | ~x5 | x7 | ~x2 | ~x3))) & (~x2 | x3 | x6 | ((~x5 | x7) & (~x4 | x5 | ~x7)));
  assign n2572 = ~x1 & ((n2573 & ~n2575) | (~x5 & ~n2574));
  assign n2573 = ~x2 & x5;
  assign n2574 = x3 ? (~x4 | ((~x6 | x7 | x0 | ~x2) & (~x0 | (x2 ? (x6 | x7) : (~x6 | ~x7))))) : ((~x6 | ~x7 | x2 | x4) & (x0 | ((x2 | ~x6 | ~x7) & (x6 | x7 | ~x2 | x4))));
  assign n2575 = (x3 | x4 | ~x6 | x7) & (~x3 | ((~x0 | ~x6 | x7) & (x6 | ~x7 | x0 | ~x4)));
  assign n2576 = x1 ? (x5 | ((x3 | (x4 ? x6 : x0)) & (x0 | (x6 & (~x3 | ~x4))))) : ((~x0 | ((~x5 | x6) & (x5 | ~x6 | ~x3 | x4))) & (~x5 | ((x6 | (x3 & x4)) & (x0 | ~x6 | (~x3 & ~x4)))));
  assign n2577 = (x1 | ((x0 | ~x3 | x4 | x5 | x6) & (~x5 | ((x3 | x4 | ~x6) & (~x0 | (x3 & ~x6)))))) & (x0 | ~x1 | ((~x3 | ~x5 | x6) & (x5 | (~x6 & (x3 | x4)))));
  assign n2578 = (n824 | n2579) & (n2556 | (~n730 & (x3 | ~n1365)));
  assign n2579 = (~x1 | x2 | x3 | ~x4 | ~x6) & (x1 | ~x2 | ~x3 | x4 | (x0 ^ ~x6));
  assign z187 = (~x0 & (x1 ? ~n2583 : ~n2582)) | ~n2584 | (x0 & ~x1 & ~n2581);
  assign n2581 = (~x5 | ((~x3 | x4 | x6 | x7) & (x3 | ~x4 | ~x7 | (x2 ^ x6)))) & (~x2 | ~x3 | ((x5 | x6 | x7) & (x4 | ~x6 | ~x7)));
  assign n2582 = (~x2 | x4 | x5 | ((x6 | x7) & (x3 | ~x6 | ~x7))) & (~x3 | ~x4 | ((~x5 | ~x6 | ~x7) & (x2 | ((~x6 | ~x7) & (~x5 | x6 | x7)))));
  assign n2583 = (~x5 | ((x3 | ((~x6 | x7 | x2 | x4) & (~x2 | (x6 ^ x7)))) & (x2 | ~x3 | x4 | ~x6 | ~x7))) & (x3 | ~x4 | ((x5 | x6 | x7) & (~x2 | ~x6 | ~x7)));
  assign n2584 = ~n2586 & n2589 & (n620 | n2585) & (x5 | n2588);
  assign n2585 = (x2 | ((x1 | ((x3 | x4) & (~x0 | (x4 ? ~x3 : ~x5)))) & (x0 | ((x3 | ~x4 | x5) & (~x1 | ~x3 | x4))) & (~x1 | (x3 ? (x4 | x5) : ~x4)))) & (x0 | ~x2 | ~x3 | (x1 & (~x4 | ~x5)));
  assign n2586 = n1421 & ((x0 & x2 & x3 & n2238) | (~x0 & ~x3 & ~n2587));
  assign n2587 = x2 ? (x4 | x6) : (~x4 | ~x6);
  assign n2588 = x0 ? (x1 | ((x3 | ~x4 | ~x6) & (x2 | ~x3 | x4 | x6))) : (~x1 | ((~x4 | x6 | ~x2 | ~x3) & (x3 | x4 | ~x6)));
  assign n2589 = (x4 | (x0 ? (x3 | (x1 ? (x2 | x6) : (~x2 | ~x6))) : (~x3 | (x1 ? (~x2 | x6) : (x2 | ~x6))))) & (x0 | ~x4 | ((~x3 | ~x6 | ~x1 | x2) & (x1 | ~x2 | x3 | x6)));
  assign z188 = ~n2593 | (~x4 & ~n2591) | (~x1 & (~n2599 | (x4 & ~n2600)));
  assign n2591 = (x2 | ~x3 | ~x5 | ~x6 | n2292) & (x3 | (n2592 & (x6 | n2292 | ~x2 | x5)));
  assign n2592 = (~x5 | x6 | ~x7 | ~x0 | ~x1 | x2) & (x0 | x1 | x7 | (x2 ? (~x5 | x6) : (x5 | ~x6)));
  assign n2593 = ~n2594 & ~n2595 & n2596 & ~n2597 & (n620 | n2598);
  assign n2594 = n664 & ((~x2 & ~x3 & x4 & n2205) | (x2 & (x3 ? (x4 & ~n800) : (~x4 & n2205))));
  assign n2595 = ~n906 & ((~x2 & ~x4 & ~x5 & x0 & x1) | (~x0 & ~x1 & x5 & (x2 ^ x4)));
  assign n2596 = ((~x3 ^ x7) | ((x0 | ~x1 | x2 | x4) & (~x0 | x1 | (~x2 ^ x4)))) & (x2 | (x1 ^ x4) | (x0 ? (x3 | x7) : (~x3 | ~x7)));
  assign n2597 = ~x0 & x2 & ((x4 & x7 & ~x1 & ~x3) | (x1 & (x3 ? (~x4 & x7) : (x4 & ~x7))));
  assign n2598 = (x3 | ~x4 | ~x5 | ~x0 | x1 | ~x2) & (x0 | x5 | ((~x3 | x4 | x1 | ~x2) & (~x1 | x2 | x3 | ~x4)));
  assign n2599 = x5 ? ((~x0 | ~x2 | ~x3 | ~x4 | ~x7) & (x0 | x2 | x3 | x4 | x7)) : (x0 ? (~x7 | (x2 ? (x3 | ~x4) : (~x3 | x4))) : (x7 | (x2 ? (~x3 ^ ~x4) : (x3 | ~x4))));
  assign n2600 = (x5 | ((x0 | x2 | ~x3 | ~x6 | x7) & (~x0 | ((x2 | x3 | x6 | x7) & (~x2 | ~x3 | (x6 ^ x7)))))) & (x0 | ~x2 | ~x3 | ~x5 | (x6 ^ x7));
  assign z189 = n2603 | n2605 | n2606 | ~n2607 | (~n2189 & ~n2602);
  assign n2602 = (x2 | ((~x1 | ((~x6 | ~x7 | x4 | ~x5) & (x5 | x6 | x7))) & (~x4 | x5 | (~x6 & ~x7)) & (x6 | ((x7 | (~x4 ^ ~x5)) & (x1 | ~x7 | (~x4 & x5)))))) & (x1 | ((~x2 | x4 | ~x5) & (~x6 | ((x7 | (~x4 ^ ~x5)) & (~x2 | (x4 & ~x5))))));
  assign n2603 = ~x4 & ((n537 & n916 & n750) | (~x6 & ~n2604));
  assign n2604 = (x0 | ~x1 | x2 | x3 | ~x5 | x7) & (x1 | ~x7 | (x0 ? (x2 ? (x3 | x5) : (~x3 | ~x5)) : (x3 | (x2 ^ x5))));
  assign n2605 = x2 & ((x3 & n2135 & x0 & ~x1) | (~x0 & (x1 ? n983 : (~x3 & n2135))));
  assign n2606 = n947 & (x1 ? (x4 & n1120) : (~x4 & ~n912));
  assign n2607 = n2608 & (n868 | ((~x0 | x1 | ~x2 | ~x3) & (x0 | ~x1 | (~x2 ^ ~x3))));
  assign n2608 = (n1716 | (~n1263 & ~n2609)) & (~n1838 | ~n677) & (~n762 | ~n2609);
  assign n2609 = x3 & ~x2 & x0 & ~x1;
  assign z190 = ~n2613 | (~x3 & (x1 ? ~n2612 : ~n2611));
  assign n2611 = (~x0 | ~x2 | ~x4 | x5 | ~x6 | x7) & (x4 | ((~x6 | x7 | x0 | x2) & (~x7 | ((~x5 | x6 | x0 | ~x2) & (~x0 | x5 | (~x2 ^ x6))))));
  assign n2612 = (~x5 | x6 | ~x7 | ~x0 | x2 | ~x4) & (x0 | ((x6 | x7 | ~x4 | ~x5) & (x4 | (x2 ? (~x6 | (~x5 ^ x7)) : (x6 | ~x7)))));
  assign n2613 = ~n2615 & (n846 | n2614) & (x0 ? n2619 : n2618);
  assign n2614 = (x1 & ((~x3 & (x2 | (~x0 & (x4 | x7)))) | (x2 & x4 & x7) | (x3 & (x0 | (~x2 & ~x4 & ~x7))))) | (~x0 & ((~x3 & x4 & x7) | (~x1 & x3 & ~x4))) | (~x1 & ((x0 & ((~x3 & ~x4) | (~x2 & x4 & ~x7))) | (~x4 & x7 & x2 & x3) | (~x2 & ~x7 & (x3 ^ ~x4)))) | (x0 & (x3 ? x4 : (~x4 & ~x7)));
  assign n2615 = x3 & ((n664 & ~n2617) | (~x1 & ~n2616));
  assign n2616 = (x0 | x2 | x4 | x5 | ~x6 | ~x7) & ((x4 ? (x5 | ~x6) : (~x5 | x6)) | (x0 ? (x2 | ~x7) : (~x2 | x7)));
  assign n2617 = (~x2 | ~x6 | (x4 ? (~x5 | ~x7) : (x5 | x7))) & (x2 | ~x4 | ~x5 | x6 | ~x7);
  assign n2618 = x1 ? ((~x2 | ~x5 | x6 | (~x3 ^ ~x4)) & (x5 | ~x6 | ((x3 | ~x4) & (x2 | ~x3 | x4)))) : ((x3 | ~x4 | ~x5 | x6) & (~x3 | ((x5 | ~x6 | ~x2 | x4) & (x2 | (x4 ? (x5 | ~x6) : (~x5 | x6))))));
  assign n2619 = (~x1 | x2 | x3 | x4 | x5 | ~x6) & (x1 | (x3 ? ((~x4 | ~x5 | x6) & (~x2 | ((~x5 | x6) & (~x4 | x5 | ~x6)))) : ((x5 | ~x6 | ~x2 | x4) & (x2 | (x4 ? (x5 | ~x6) : (~x5 | x6))))));
  assign z191 = n1521 | n2621 | n2623 | ~n2627 | (~n927 & ~n2626);
  assign n2621 = ~x5 & ~n2622;
  assign n2622 = x1 ? ((x0 | ((x2 | ~x4 | ~x6) & (x4 | x6 | ~x2 | x3))) & (x2 | ((x3 | ~x4 | ~x6) & (x4 | x6 | ~x0 | ~x3)))) : ((x4 | ~x6 | x0 | ~x2) & (~x3 | ~x4 | (x0 ? (~x2 ^ ~x6) : (~x2 | x6))));
  assign n2623 = ~x0 & ((x2 & ~n2624) | (n563 & ~n2625));
  assign n2624 = (x5 | ~x6 | ~x7 | x1 | ~x3 | ~x4) & (x4 | ~x5 | ((~x6 | x7 | x1 | ~x3) & (~x1 | (x3 ? (x6 | x7) : (~x6 | ~x7)))));
  assign n2625 = (~x1 | x4 | ~x5 | x6 | ~x7) & (x5 | ((~x1 | x7 | (~x4 ^ x6)) & (x6 | ~x7 | x1 | ~x4)));
  assign n2626 = ((~x3 ^ x5) | ((x0 | ~x1 | ~x2 | x6) & (x2 | ~x6 | ~x0 | x1))) & (x2 | ((x6 | (~x0 ^ x3) | (x1 ^ x5)) & (~x3 | ~x5 | ~x6 | x0 | x1))) & (x1 | ~x2 | x3 | (x0 ? (x5 | ~x6) : (x5 ^ x6)));
  assign n2627 = (n2500 | n2629) & (~n568 | ~n1476) & (~x5 | n2628);
  assign n2628 = (x0 | ~x1 | ~x2 | ~x3 | (~x4 ^ x6)) & (x1 | (x0 ? ((~x4 | ~x6 | x2 | ~x3) & (~x2 | x4 | x6)) : ((~x4 | ~x6 | ~x2 | ~x3) & (x2 | ((~x4 | x6) & (x3 | x4 | ~x6))))));
  assign n2629 = (~x0 | x1 | ~x2 | ~x6 | x7) & (x0 | x2 | ~x7 | (~x1 ^ x6));
  assign z192 = ~n2634 | (x2 & ~n2638) | (~x2 & ~n2631) | (~n912 & ~n2637);
  assign n2631 = x0 ? n2633 : n2632;
  assign n2632 = ((~x5 ^ ~x6) | ((x1 | ~x3 | ~x7) & (x4 | x7 | ~x1 | x3))) & (~x5 | ~x6 | ~x7 | x1 | ~x4) & (~x1 | (x3 ? ((~x6 | x7 | x4 | x5) & (x6 | ~x7 | ~x4 | ~x5)) : (x5 | ~x7 | (~x4 ^ x6))));
  assign n2633 = (x5 | ~x6 | x7 | ~x1 | x3 | ~x4) & (x1 | (x3 ? (x5 ? (~x6 | x7) : ((x6 | x7) & (~x4 | ~x6 | ~x7))) : ((~x6 | ~x7 | x4 | ~x5) & (~x4 | x6 | (~x5 & ~x7)))));
  assign n2634 = x4 ? n2636 : n2635;
  assign n2635 = x1 ? ((x2 | ((x3 | ~x5 | ~x7) & (x5 | x7 | ~x0 | ~x3))) & (x0 | (x2 ? (x5 | (x3 ^ x7)) : (~x5 | ~x7)))) : ((~x0 | ((x3 | x5 | ~x7) & (~x2 | ~x5 | x7))) & (x2 | x3 | (~x5 ^ x7)) & (x0 | (x2 ? (x3 ? (x5 | x7) : (~x5 | ~x7)) : (~x5 | x7))));
  assign n2636 = ((~x5 ^ x7) | ((~x2 | x3 | ~x0 | x1) & (x0 | (x1 ? (~x2 | ~x3) : (x2 | x3))))) & (~x1 | x2 | ((x3 | ~x5 | ~x7) & (x5 | x7 | x0 | ~x3))) & (x0 | x1 | ~x2 | (x3 ? (x5 | x7) : (~x5 | ~x7)));
  assign n2637 = x1 ? (x3 | ((x4 | x7 | ~x0 | x2) & (x0 | (x2 ? ~x7 : (~x4 | x7))))) : ((x0 | ~x2 | x3 | x4 | x7) & (~x3 | (x0 ? (x2 ? (~x4 | x7) : (x4 | ~x7)) : (~x4 | (~x2 ^ ~x7)))));
  assign n2638 = (n846 | n2640) & (~n1743 | ~n1621) & (x1 | n2639);
  assign n2639 = (x0 | ~x3 | ~x5 | (x4 ? (~x6 | x7) : (x6 | ~x7))) & (x3 | ((x5 | ~x6 | x7 | x0 | ~x4) & (~x0 | ((x6 | x7 | x4 | x5) & (~x6 | ~x7 | ~x4 | ~x5)))));
  assign n2640 = (~x0 | x1 | ~x3 | ~x7) & (x0 | ~x1 | x7 | (~x3 ^ x4));
  assign z193 = n2643 | ~n2645 | (~n662 & ~n2642);
  assign n2642 = (x0 | (x1 ? ((~x2 | x3 | x4) & (~x4 | ~x5 | x2 | ~x3)) : (~x3 | (x2 ? (~x4 | x5) : x4)))) & (x1 | (((~x0 & ~x5) | (x2 ? (~x3 | x4) : (x3 | ~x4))) & (~x0 | x3 | ~x5 | (x2 & ~x4))));
  assign n2643 = x4 & ((n985 & n540 & n1546) | (~x5 & ~n2644));
  assign n2644 = (x2 | ((x3 | ~x6 | x7 | x0 | ~x1) & (~x0 | ((x6 | ~x7 | ~x1 | x3) & (x1 | ~x3 | ~x6 | x7))))) & (x0 | ~x2 | x6 | ~x7 | (x1 ^ x3));
  assign n2645 = x6 ? ((x7 | n2646) & n2648) : (n2647 & (~x7 | n2646));
  assign n2646 = (x2 | ((x0 | ~x1 | x3 | ~x4 | ~x5) & (~x0 | ((~x4 | ~x5 | x1 | ~x3) & (~x1 | x3 | x4))))) & (x4 | ((x1 | ~x2 | x3 | x5) & (x0 | (~x2 & x5) | (x1 ^ x3))));
  assign n2647 = ((x3 ? (x4 | x5) : (~x4 | ~x5)) | (x0 ? (~x1 | x2) : (x1 | ~x2))) & ((~x4 ^ x5) | ((x0 | x2 | (x1 ^ x3)) & (~x2 | x3 | ~x0 | x1))) & (~x0 | x1 | x2 | x3 | x4 | x5) & (~x3 | ~x4 | ~x5 | x0 | ~x1 | ~x2);
  assign n2648 = ((x2 ^ x4) | (x0 ? (x1 | ~x3) : (~x1 | x3))) & (x1 | ~x3 | ~x4 | (x2 ? ~x5 : x0));
  assign z194 = n2651 | n2657 | n2658 | ~n2659 | (~x0 & ~n2650);
  assign n2650 = (x2 | x3 | x4 | ~x5 | x7) & (~x1 | (x2 ? ((x3 | ~x4 | ~x5 | x7) & (x5 | ~x7 | ~x3 | x4)) : ((~x4 | ~x5 | ~x7) & (x3 | x4 | x7))));
  assign n2651 = ~x6 & (n2652 | n2654 | (n723 & n650 & n677));
  assign n2652 = x4 & ((~x3 & n2205 & n677) | (n1156 & ~n2653));
  assign n2653 = (~x0 | ~x1 | x2 | x3) & (x0 | ~x2 | (x1 ^ x3));
  assign n2654 = ~n2655 & ~n2656;
  assign n2655 = x2 ? (x3 | ~x5) : (~x3 | x5);
  assign n2656 = (~x4 | x7 | ~x0 | x1) & (x4 | ~x7 | x0 | ~x1);
  assign n2657 = ~n906 & ((~x2 & ~x4 & ~x5 & x0 & x1) | (~x1 & ((~x4 & ~x5 & ~x0 & x2) | (x5 & (x0 ? (x2 ^ ~x4) : (~x2 & x4))))));
  assign n2658 = ~n592 & (x0 ? ((x3 & ~x5 & ~x1 & x2) | (x1 & ~x2 & ~x3 & x5)) : ((~x1 & ~x2 & ~x5) | (x2 & (x1 ? (x3 ^ ~x5) : (~x3 & x5)))));
  assign n2659 = n2662 & (n2354 | n2661) & (~x6 | ~n2095 | n2660);
  assign n2660 = (x0 | ~x1 | ~x2 | ~x3 | x7) & (x2 | ((~x0 | (x1 ? (x3 | x7) : (~x3 | ~x7))) & (x3 | ~x7 | x0 | ~x1)));
  assign n2661 = (~x0 | x1 | ~x2 | x4 | x6 | ~x7) & (x0 | ~x4 | x7 | (x1 ? (x2 | x6) : (~x2 | ~x6)));
  assign n2662 = x4 ? ((x5 | n2663) & (~x7 | ~n1887 | (x3 & ~x5))) : (x5 ? n2663 : (x7 | ~n1887));
  assign n2663 = (~x2 | x3 | x7 | ~x0 | x1) & (x0 | ~x3 | (x1 ? (x2 | x7) : (~x2 | ~x7)));
  assign z195 = ~n2667 | (x6 & (x2 ? ~n2665 : ~n2666));
  assign n2665 = ((x3 ? (~x4 | x7) : (x4 | ~x7)) | (x0 ? (x1 | x5) : (~x1 | ~x5))) & (x1 | ~x5 | ((~x4 | x7 | x0 | x3) & (x4 | ~x7 | ~x0 | ~x3)));
  assign n2666 = (~x1 | x3 | ~x4 | ~x5 | x7) & (~x3 | ((~x0 | x1 | ~x4 | ~x5 | x7) & (x0 | x4 | ~x7 | (~x1 ^ x5))));
  assign n2667 = n2670 & n2673 & (x5 ? (x6 | n2669) : n2668);
  assign n2668 = x1 ? (x4 | ((x3 | ~x6 | ~x0 | x2) & (x0 | ~x2 | (x3 ^ x6)))) : ((x0 | ~x2 | x3 | x4 | ~x6) & (~x3 | ((~x0 | (x2 ? x6 : (x4 | ~x6))) & (x4 | x6 | x0 | x2))));
  assign n2669 = x1 ? ((x3 | x4 | x7 | ~x0 | x2) & (x0 | ~x3 | (x2 ? (x4 | x7) : (~x4 | ~x7)))) : (x0 ? ((x2 | ~x3 | x4 | x7) & (~x4 | ~x7 | ~x2 | x3)) : ((~x4 | ~x7 | x2 | x3) & (~x2 | (x3 ? (~x4 | ~x7) : (x4 | x7)))));
  assign n2670 = ~n2672 & (n2671 | (~n965 & (~x4 | n912)));
  assign n2671 = (x0 | ~x2 | (x1 ^ x3)) & (x2 | ((~x1 | x3) & (~x0 | x1 | ~x3)));
  assign n2672 = ~x0 & x1 & ((x4 & ~x5 & x2 & ~x3) | (~x2 & x3 & ~x4 & x5));
  assign n2673 = ~n2674 & (~x6 | ~n1701 | n2675);
  assign n2674 = ~x1 & ((~x0 & x3 & (x2 ? (~x4 & x5) : (x4 & ~x5))) | (~x3 & ~x4 & x5 & (x0 | ~x2)));
  assign n2675 = (x2 | ~x3 | x0 | ~x1) & (x1 | (x0 ? (~x2 | x3) : (~x2 ^ ~x3)));
  assign z196 = ~n2682 | (x0 ? (n2681 | (x5 & ~n2680)) : ~n2677);
  assign n2677 = (n1446 | n2679) & (~n2285 | ~n1621) & (~x3 | n2678);
  assign n2678 = (~x1 | x2 | x4 | x5 | x6 | x7) & (~x6 | (x1 ? ((~x5 | ~x7 | ~x2 | ~x4) & (x2 | (x4 ? (~x5 | x7) : (x5 | ~x7)))) : ((x2 | x4 | ~x5 | ~x7) & (~x2 | ~x4 | x5 | x7))));
  assign n2679 = (~x1 | ~x3 | x5 | ~x6 | x7) & (x1 | x3 | ~x5 | x6 | ~x7);
  assign n2680 = x1 ? (x2 | x3 | (x4 ? (~x6 | ~x7) : (~x6 ^ x7))) : (x6 ? (x2 ? (x3 ? (x4 | ~x7) : (~x4 | x7)) : (~x3 | (x4 ^ x7))) : (~x7 | ((x3 | ~x4) & (x2 | ~x3 | x4))));
  assign n2681 = n709 & ((~x3 & ~x4 & ~x6 & ~x7) | (x6 & (x2 ? (x7 & (x3 ^ ~x4)) : (~x7 & (~x3 ^ ~x4)))));
  assign n2682 = ~n2685 & (x6 ? n2683 : n2684) & (n1323 | n2686);
  assign n2683 = (~x3 | x4 | x5 | ~x0 | x1 | ~x2) & (x0 | ((~x1 | x2 | x3 | x5) & (x4 | (x1 ? ((x3 | x5) & (~x2 | ~x3 | ~x5)) : (x2 ? (x3 | ~x5) : (~x3 | x5))))));
  assign n2684 = ((~x4 ^ x5) | ((~x0 | x1 | x3) & (x2 | ~x3 | x0 | ~x1))) & (~x4 | ((x0 | ~x1 | ~x2 | x3 | ~x5) & (x1 | ((x2 | x3 | x5) & (~x3 | (x0 ? (~x2 | ~x5) : (~x2 ^ x5)))))));
  assign n2685 = ~n783 & ((~x0 & ~x1 & x5 & (x2 ^ ~x3)) | (~x5 & (x0 ? (~x2 & (x1 ^ x3)) : (x2 & (~x1 ^ x3)))));
  assign n2686 = (x5 | x7 | (x0 ? (x1 ? (x2 | x4) : (~x2 | ~x4)) : (x1 | (~x2 ^ x4)))) & (x0 | ~x5 | ~x7 | (x1 ? (~x2 ^ x4) : (~x2 | ~x4)));
  assign z197 = n2688 | ~n2691 | ~n2695 | (~n662 & ~n2690);
  assign n2688 = ~x1 & ((n1415 & n943) | (n543 & ~n2689));
  assign n2689 = (x2 | x3 | x5 | (~x0 & ~x4)) & (x0 | ((~x2 | x3 | x4 | ~x5) & (~x3 | ((~x4 | x5) & (x2 | x4 | ~x5)))));
  assign n2690 = x5 ? (x1 ? ((x0 | ((x3 | x4) & (~x2 | ~x3 | ~x4))) & (x2 | x3 | ~x4)) : ((x3 | ~x4 | x0 | ~x2) & (~x3 | (x0 ? (~x2 ^ x4) : (x2 | x4))))) : (x1 ? ((x3 | x4 | ~x0 | x2) & (x0 | ~x3 | (~x2 ^ x4))) : ((~x0 | ((x3 | ~x4) & (x2 | ~x3 | x4))) & (x2 | x3 | ~x4) & (x0 | ~x2 | (~x3 ^ ~x4))));
  assign n2691 = (n1350 | n2694) & (n868 | n2693) & (~n694 | ~n2692);
  assign n2692 = x7 & x5 & ~x3 & ~x4;
  assign n2693 = (x1 | (x0 ? (~x2 | (~x3 ^ x7)) : ((x3 | x6 | ~x7) & (x2 | ~x3 | x7)))) & (x0 | ((x6 | ~x7 | ~x2 | ~x3) & (~x1 | (x2 ? (x3 | x7) : (~x3 | ~x7)))));
  assign n2694 = (~x0 | x1 | ~x3 | ~x7) & (x0 | x7 | (~x1 ^ ~x3));
  assign n2695 = (x7 | n2696) & (~x1 | x6 | ~x7 | n2697);
  assign n2696 = x1 ? (x2 | x3 | x5 | (x0 & ~x4)) : ((~x3 | x4 | ~x5 | x0 | ~x2) & (~x0 | ((x2 | ~x3 | ~x4 | x5) & (x3 | x4 | ~x5))));
  assign n2697 = (~x3 | x4 | x5 | ~x0 | x2) & (x0 | ((~x2 | (x3 ? (x4 | ~x5) : (~x4 | x5))) & (x2 | x3 | x4 | ~x5)));
  assign z198 = ~n2706 | (~x2 & ~n2699);
  assign n2699 = ~n2701 & n2702 & ~n2704 & ~n2705 & (x3 | n2700);
  assign n2700 = x0 ? (x1 | ((x6 | x7 | x4 | x5) & (~x6 | ~x7 | ~x4 | ~x5))) : (~x1 | ((~x6 | ~x7 | ~x4 | x5) & (x4 | x7 | (~x5 ^ x6))));
  assign n2701 = (x4 ^ ~x5) & ((x0 & ~x6 & (~x1 ^ ~x3)) | (~x0 & ~x1 & x3 & x6));
  assign n2702 = ~n2703 & (~n587 | ~n1743) & (~n586 | (~n872 & ~n838));
  assign n2703 = ~x0 & ((~x1 & ~x3 & x4 & ~x6 & ~x7) | (x6 & x7 & x1 & ~x4));
  assign n2704 = ~x0 & ((~x1 & ~x3 & ~x4 & x5 & x6) | (x1 & x4 & ~x6 & (x3 ^ x5)));
  assign n2705 = ~n627 & ((x3 & ~x6 & ~x7 & ~x0 & ~x1) | (x0 & x6 & x7 & (~x1 ^ ~x3)));
  assign n2706 = (n620 | n2707) & (~x2 | (~n2709 & (x1 | n2708)));
  assign n2707 = x1 ? ((x0 | ((~x4 | ~x5 | x2 | ~x3) & (~x2 | (x3 ? (x4 | ~x5) : (~x4 | x5))))) & (x2 | x4 | ((~x3 | x5) & (~x0 | x3 | ~x5)))) : (((~x3 ^ x5) | (x0 ? (~x2 | ~x4) : (~x2 ^ x4))) & (~x3 | ~x4 | ~x5 | x0 | ~x2) & (x4 | ((x2 | x3 | x5) & (~x0 | ((x3 | x5) & (x2 | ~x3 | ~x5))))));
  assign n2708 = x0 ? ((~x3 | ((x5 | ~x6 | ~x7) & (x4 | ~x5 | x6))) & (x3 | ((~x5 | ~x6 | ~x7) & (~x4 | x5 | x6))) & (~x6 | ~x7 | (~x4 ^ ~x5))) : ((~x3 | ((x5 | x6 | x7) & (x4 | ~x5 | ~x6))) & (x6 | x7 | (~x4 ^ ~x5)) & (x3 | ((~x5 | x6 | x7) & (~x4 | x5 | ~x6))));
  assign n2709 = n664 & (x6 ? (x3 ? (x4 & ~x5) : (x4 ? x5 : (~x5 & x7))) : (x3 ? (~x7 & (~x4 | x5)) : (~x4 & x5)));
  assign z199 = ~n2715 | (x0 ? ~n2711 : (x2 ? ~n2714 : ~n2713));
  assign n2711 = x1 ? (~n563 | ~n568) : n2712;
  assign n2712 = x5 ? ((x2 | x3 | ~x4 | ~x6 | x7) & (x4 | ((~x3 | x6 | x7) & (x2 | ~x7 | (x3 ^ x6))))) : ((~x6 | ((x2 | x3 | ~x4 | ~x7) & ((~x3 ^ ~x4) | (x2 ^ x7)))) & (x2 | x6 | (x3 ? (x4 | ~x7) : (~x4 | x7))));
  assign n2713 = x1 ? ((~x3 | x4 | x5 | ~x6 | ~x7) & (x3 | ~x4 | ~x5 | x6 | x7)) : (((~x3 ^ ~x4) | (x5 ? (x6 | ~x7) : (~x6 | x7))) & (~x3 | x4 | x5 | x6 | ~x7) & (x3 | ~x4 | ~x5 | ~x6 | x7) & ((x6 ^ x7) | (x3 ? (x4 | ~x5) : (~x4 | x5))));
  assign n2714 = ((~x4 ^ ~x7) | (((~x1 ^ ~x3) | (~x5 ^ ~x6)) & (~x5 | x6 | ~x1 | x3) & (x5 | ~x6 | x1 | ~x3))) & ((~x1 ^ ~x3) | ((~x6 | ~x7 | x4 | x5) & (x6 | x7 | ~x4 | ~x5)));
  assign n2715 = ~n2719 & (n620 | n2716) & (x2 ? n2718 : n2717);
  assign n2716 = (~x2 | ((x0 | ~x1 | x3 | x4 | x5) & (x1 | ((~x3 | ~x4 | ~x5) & (~x0 | x4 | (~x3 ^ x5)))))) & (~x1 | x2 | ((x3 | ~x4 | x5) & (x4 | ~x5 | x0 | ~x3)));
  assign n2717 = (~x4 | ~x5 | ~x7 | ~x0 | x1 | ~x3) & (~x1 | ((~x5 | ~x7 | x3 | ~x4) & (x5 | x7 | ~x3 | x4) & (((x3 | x4) & (x0 | ~x3 | ~x4)) | (~x5 ^ x7))));
  assign n2718 = ((x4 ? (x5 | x7) : (~x5 | ~x7)) | ((x0 | ~x1 | x3) & (x1 | ~x3))) & (~x0 | x1 | x3 | (x4 ? (~x5 ^ x7) : (x5 | x7)));
  assign n2719 = ~n1429 & ((x0 & ~x1 & x2 & ~x3 & x4) | (x1 & ~x2 & ((~x3 & ~x4) | (~x0 & x3 & x4))));
  assign z200 = n2721 | ~n2725 | ~n2732 | (~x2 & ~n2724);
  assign n2721 = ~x1 & ((n2205 & ~n2723) | (~x5 & ~n2722));
  assign n2722 = x6 ? (~x7 | ((x3 | ~x4 | x0 | ~x2) & (~x0 | (x2 ? (~x3 ^ ~x4) : (~x3 | x4))))) : (((x4 ^ x7) | (x0 ? (~x2 | x3) : (x2 | ~x3))) & (x3 | x4 | ~x7 | ~x0 | x2));
  assign n2723 = (x0 | x2 | ~x3 | x4 | ~x6) & (~x0 | ~x2 | ((~x4 | x6) & (x3 | x4 | ~x6)));
  assign n2724 = (x0 | ((~x7 | (~x4 ^ ~x5) | (x3 ^ x6)) & (x3 | x7 | (x4 ? (x5 | ~x6) : (~x5 | x6))))) & (x3 | ((~x6 | ~x7 | x4 | ~x5) & (~x0 | ~x4 | x5 | x6 | x7)));
  assign n2725 = ~n2727 & n2729 & ((x6 & (x7 | n2728)) | (n2726 & (n2728 | (~x6 & ~x7))));
  assign n2726 = x0 ? ((x4 | ~x5 | x2 | x3) & (x1 | ~x2 | ~x3 | ~x4 | x5)) : (x2 | ~x3 | (x1 ? (x4 | x5) : (~x4 | ~x5)));
  assign n2727 = ~n1041 & ((~x2 & n985 & x0 & ~x1) | (~x0 & ((x2 & n916) | (x1 & ~x2 & n985))));
  assign n2728 = (x2 | ((~x4 | ~x5 | ~x0 | x3) & (x5 | ((~x0 | (x1 ? (x3 | x4) : (~x3 | ~x4))) & (~x3 | ~x4 | x0 | ~x1))))) & (x0 | ~x2 | x4 | ((x3 | ~x5) & (x1 | ~x3 | x5)));
  assign n2729 = (n2730 | n2731) & (~n1365 | ~n814 | ~n1176);
  assign n2730 = x3 ? (x4 | x6) : (~x4 | ~x6);
  assign n2731 = (x0 | x1 | ~x2 | ~x5) & (~x0 | x2 | x5);
  assign n2732 = (n857 | n2734) & (~n616 | n2733);
  assign n2733 = (~x3 | ~x4 | x5 | ~x6 | ~x7) & (x7 | ((x3 | x4 | x5 | x6) & (~x4 | (x3 ? (~x5 ^ ~x6) : (~x5 | x6)))));
  assign n2734 = (x2 | ~x3 | x4 | ~x5 | x6 | x7) & (~x2 | ((~x5 | ~x6 | ~x7 | x3 | ~x4) & (~x3 | x4 | (x5 ? (x6 | ~x7) : (~x6 | x7)))));
  assign z201 = ~n2740 | (x0 ? ~n2736 : (x5 ? ~n2739 : ~n2738));
  assign n2736 = x1 ? (~n563 | ~n568) : n2737;
  assign n2737 = ((~x2 & x4) | ((~x6 | ~x7 | ~x3 | x5) & (x6 | x7 | x3 | ~x5))) & (x2 | ~x3 | ~x4 | x5 | x6 | x7) & (x3 | ((~x6 | x7 | ~x4 | x5) & (x2 | ((x5 | ~x6 | x7) & (x6 | ~x7 | ~x4 | ~x5)))));
  assign n2738 = x3 ? (x1 ? ((x4 | ~x6 | ~x7) & (x6 | x7 | ~x2 | ~x4)) : (x7 | ((x4 | x6) & (x2 | ~x4 | ~x6)))) : (~x6 | (x1 & x2) | (x4 ^ x7));
  assign n2739 = (~x7 | (x1 ? (~x2 | ~x4 | (x3 ^ x6)) : (x4 | ((x3 | x6) & (x2 | ~x3 | ~x6))))) & (x6 | x7 | (x1 ? (x3 | x4) : (~x3 | ~x4)));
  assign n2740 = n2742 & ~n2746 & (n846 | n2741) & (n620 | n2748);
  assign n2741 = (x1 | (x0 ? ((~x4 | x7 | ~x2 | ~x3) & (x3 | x4 | ~x7)) : (~x4 | ((~x3 | ~x7) & (x2 | x3 | x7))))) & (~x0 | x2 | x3 | x4 | ~x7) & (x0 | ~x3 | ((~x1 | x4 | x7) & (x2 | ~x4 | ~x7)));
  assign n2742 = (~x3 | n2745) & (n910 | (x0 ? n2744 : (x3 | ~n2743)));
  assign n2743 = ~x7 & x4 & ~x5;
  assign n2744 = (~x3 | x4 | x5 | x7) & (x3 | ~x4 | ~x5 | ~x7);
  assign n2745 = x0 ? (x1 | x2 | (x4 ? (~x5 ^ x7) : (x5 | x7))) : (x1 ? (~x4 | ((~x5 | x7) & (~x2 | x5 | ~x7))) : (x4 | (~x5 ^ x7)));
  assign n2746 = n2747 & ((x0 & ~x2 & ~x4 & x5 & ~x7) | (~x0 & ((~x4 & x5 & x7) | (~x5 & ~x7 & x2 & x4))));
  assign n2747 = x1 & ~x3;
  assign n2748 = x0 ? ((x4 | ~x5 | x1 | ~x3) & (~x1 | x2 | x3 | ~x4 | x5)) : (x3 | ((~x4 | ~x5 | x1 | ~x2) & (~x1 | (x2 ? (x4 | x5) : (~x4 | ~x5)))));
  assign z202 = ~n2752 | (x4 ? (x7 ? ~n2750 : ~n2751) : (x7 ? ~n2751 : ~n2750));
  assign n2750 = x0 ? ((~x1 | x2 | x3 | ~x5 | x6) & (x1 | ((x2 | ((x5 | x6) & (x3 | ~x5 | ~x6))) & (x6 | ((x3 | x5) & (~x2 | ~x3 | ~x5)))))) : ((x1 | x2 | x3 | ~x5 | x6) & (~x6 | (x1 ? (x2 ^ x5) : (~x2 | x5))));
  assign n2751 = (~x1 | ((x0 | ~x5 | x6) & (x3 | ~x6 | ~x0 | x2))) & (x0 | x2 | x3 | x5 | x6) & (x1 | ((~x5 | ~x6 | x0 | x2) & (x5 | (x0 ? (~x6 | (~x2 & ~x3)) : x6))));
  assign n2752 = n2757 & ((x2 & (x3 ? n2755 : n2754)) | (n2753 & (x3 ? n2755 : ~x2)));
  assign n2753 = (~x0 | x1 | x3 | x4 | x5 | ~x6) & (x0 | ((x4 | ~x5 | x6 | x1 | ~x3) & (~x1 | ~x4 | (x3 ? (x5 | x6) : (~x5 | ~x6)))));
  assign n2754 = (~x5 | x6 | ~x7 | ~x0 | x1 | ~x4) & (x0 | x4 | ~x6 | (x1 ? (x5 | x7) : (~x5 | ~x7)));
  assign n2755 = (~n568 | ~n1546) & (n1545 | (~n2756 & (~n738 | ~n1835)));
  assign n2756 = x7 & x4 & ~x0 & x1;
  assign n2757 = ~n2759 & ~n2760 & (x5 | n571 | ~n2758);
  assign n2758 = x2 & ~x0 & x1;
  assign n2759 = ~x2 & ((x0 & ~x6 & (x1 ? (~x4 & ~x5) : (x4 & x5))) | (x4 & ~x5 & x6 & ~x0 & ~x1));
  assign n2760 = ~x1 & x2 & x5 & (x0 ? (~x4 & x6) : (~x4 ^ x6));
  assign z203 = n2762 | n2766 | ~n2768 | (~n912 & ~n2765);
  assign n2762 = ~x0 & (x4 ? ~n2764 : ~n2763);
  assign n2763 = x5 ? (x1 ? (x7 | (x2 ? (~x3 | x6) : ~x6)) : (~x6 | ~x7 | (x2 ^ ~x3))) : (x1 ? ((x2 | x6 | x7) & (~x2 | x3 | ~x6 | ~x7)) : (x3 | (x2 ? (x6 | ~x7) : (~x6 | x7))));
  assign n2764 = x1 ? (x2 | x3 | (x5 ? (~x6 ^ x7) : (x6 | x7))) : (x2 ? ((x6 | ~x7 | x3 | x5) & (~x6 | x7 | ~x3 | ~x5)) : (~x3 | ~x7 | (~x5 ^ ~x6)));
  assign n2765 = (~x3 | ((x0 | (x1 ? (x2 ? (~x4 | x7) : ~x7) : (x2 | x7))) & (~x2 | ~x4 | ~x7 | ~x0 | x1))) & (x2 | x3 | ((x1 | ~x4 | x7) & (~x0 | (x1 ^ x7))));
  assign n2766 = x0 & ((~x1 & ~n2767) | (n1082 & n559));
  assign n2767 = x2 ? (x7 | ((~x4 | ~x5 | ~x6) & (~x3 | (~x5 ^ ~x6)))) : (~x7 | (x5 ? (~x6 | (x3 & x4)) : x6));
  assign n2768 = (x1 | n2771) & (n1099 | n2770) & (x0 | ~x1 | n2769);
  assign n2769 = (x5 | ((x2 | (x3 ? (~x4 | x7) : ~x7)) & (~x2 | x3 | x4 | x7))) & (~x2 | ~x5 | ~x7 | (~x3 ^ ~x4));
  assign n2770 = (x0 | ~x2 | ~x5 | (x1 ^ x7)) & (x5 | ((x0 | ~x1 | ~x2 | x7) & (~x0 | (x1 ? (x2 | x7) : (~x2 | ~x7)))));
  assign n2771 = (~x0 | ((~x2 | x3 | x4 | x5 | ~x7) & (~x5 | x7 | x2 | ~x3))) & (~x2 | x3 | x4 | ~x5 | x7) & (x0 | ~x7 | (x2 ? (~x3 | x5) : (x3 | ~x5)));
  assign z204 = ~n2777 | (x7 ? ~n2775 : (x3 ? ~n2774 : ~n2773));
  assign n2773 = (x4 | ((x0 | ~x5 | (x1 ? (~x2 | x6) : x2)) & (~x0 | ~x1 | x2 | x5 | ~x6))) & (x1 | ~x2 | ~x4 | (x0 ? (x5 ^ x6) : (~x5 | x6)));
  assign n2774 = (x4 | ~x5 | ~x6 | x0 | ~x1 | ~x2) & (x6 | (x0 ? (x2 | (x1 ? (x4 | x5) : (~x4 | ~x5))) : (~x2 | x5 | (~x1 ^ x4))));
  assign n2775 = (x0 | x6 | n2776) & (~x6 | ~n650 | ~n670 | ~x0 | x5);
  assign n2776 = (~x3 | x4 | x5 | x1 | x2) & (x3 | ((~x4 | ~x5 | x1 | ~x2) & (~x1 | (x2 ? (x4 | ~x5) : (~x4 | x5)))));
  assign n2777 = n2779 & (x6 ? (x7 ? (n2778 & n2781) : n2780) : (x7 ? (n2780 & n2781) : n2778));
  assign n2778 = (x2 | ((~x3 | x4 | ~x5 | ~x0 | x1) & (~x4 | (x0 ? (x1 ? x3 : (~x3 | x5)) : (~x1 | ~x3))))) & (x0 | ~x2 | x3 | ((x4 | x5) & (x1 | (x4 & x5))));
  assign n2779 = x0 ? (x1 | (x2 ? (x3 ? (~x4 | ~x6) : (x4 | x6)) : (x3 | ~x6))) : ((~x1 | x3 | ~x4 | (~x2 ^ x6)) & (~x3 | ((x2 | x4 | ~x6) & (x1 | (x2 ? (x4 | x6) : ~x6)))));
  assign n2780 = (x1 | ((~x0 | ~x2 | ~x3 | x4) & (x3 | ~x4 | x0 | x2))) & (x0 | ((~x2 | ~x3 | ~x4) & (~x1 | x2 | x3 | x4)));
  assign n2781 = (x0 | ~x1 | ~x2 | ~x3 | x4 | x6) & (x3 | ((x0 | x1 | x2 | x4 | x6) & (~x0 | ((~x4 | x6 | x1 | ~x2) & (~x1 | x2 | x4 | ~x6)))));
  assign z205 = ~n2784 | (x4 & (n2783 | (n543 & n916 & n924)));
  assign n2783 = n904 & (x0 ? ((x2 & ~x5 & x6 & ~x7) | (~x6 & x7 & ~x2 & x5)) : ((~x2 & x5 & x6 & x7) | (x2 & ~x5 & (x6 ^ ~x7))));
  assign n2784 = n2789 & (x4 | n2785) & (x5 ? n2787 : n2788);
  assign n2785 = (x2 | n2786) & (n1107 | ((~x0 | ~x1 | x2 | x6) & (x0 | (x1 ? (~x2 | ~x6) : (x2 | x6)))));
  assign n2786 = (x5 | ~x6 | x7 | x0 | x1) & (~x0 | ((x1 | ~x3 | x5 | x6 | x7) & (~x1 | x3 | ~x5 | ~x6 | ~x7)));
  assign n2787 = (x1 | ((x0 | ~x2 | ~x4 | (x3 ^ x7)) & ((~x3 ^ x7) | (x0 ? (~x2 | ~x4) : (x2 | x4))))) & (x0 | ~x1 | ((~x4 | x7 | x2 | x3) & (x4 | ~x7 | ~x2 | ~x3)));
  assign n2788 = x0 ? ((~x1 | x2 | x3 | x4 | x7) & (x1 | ~x4 | (x2 ? (x3 | x7) : (~x3 | ~x7)))) : (~x2 | ((~x4 | ~x7 | x1 | x3) & (~x1 | x4 | (~x3 ^ x7))));
  assign n2789 = x0 ? ((x4 | ~x7 | x1 | ~x3) & (x3 | ((~x1 | x2 | ~x4 | ~x7) & (x1 | x7 | (x2 & x4))))) : (((~x3 ^ x7) | (x1 ? (x2 | x4) : (~x2 ^ x4))) & (~x1 | ~x4 | ((~x3 | ~x7) & (~x2 | x3 | x7))));
  assign z206 = n2791 | n2795 | ~n2798 | (~x0 & ~n2794);
  assign n2791 = ~x1 & (x6 ? ~n2793 : ~n2792);
  assign n2792 = x0 ? ((x2 | ~x3 | x4 | x5 | x7) & (~x2 | ((~x5 | ~x7 | x3 | x4) & (x5 | x7 | ~x3 | ~x4)))) : (x2 | ((x3 | x4 | (~x5 ^ x7)) & (x5 | ~x7 | ~x3 | ~x4)));
  assign n2793 = (x2 | ~x3 | ~x4 | ~x5 | x7) & (~x7 | ((~x0 | x2 | x3 | x4 | ~x5) & (x0 | x5 | (x2 ? (~x3 | x4) : (x3 | ~x4)))));
  assign n2794 = (x1 | ~x2 | ((~x5 | ~x6 | x3 | x4) & (x5 | x6 | ~x3 | ~x4))) & (x2 | ((x1 | ~x3 | ~x4 | ~x5 | x6) & (x5 | ((x4 | ~x6 | x1 | x3) & (~x1 | (x3 ? (x4 | ~x6) : (~x4 | x6)))))));
  assign n2795 = x1 & ((n616 & ~n2797) | (~x2 & ~n2796));
  assign n2796 = x0 ? ((~x3 | x4 | x5 | ~x6 | x7) & (~x5 | x6 | ~x7 | x3 | ~x4)) : (~x4 | ~x6 | (x3 ? (~x5 | ~x7) : (x5 | x7)));
  assign n2797 = (~x5 | x6 | x7 | x3 | x4) & (~x3 | x5 | (x4 ? (x6 | ~x7) : (~x6 | x7)));
  assign n2798 = ~n2800 & ~n2802 & (n783 | n2801) & (~x0 | n2799);
  assign n2799 = (~x1 | x2 | ~x3 | x4 | x5 | x6) & (x1 | ((x2 | ~x3 | ~x4 | ~x5 | x6) & (~x2 | x4 | ~x6 | (~x3 ^ x5))));
  assign n2800 = x1 & ((x4 & x5 & ~x0 & x2) | (~x4 & ((~x2 & ~x3 & ~x5) | (~x0 & (x5 ? ~x2 : ~x3)))));
  assign n2801 = (~x0 | ~x1 | x2 | x3 | ~x5) & (x0 | ~x3 | x5 | (~x1 ^ ~x2));
  assign n2802 = ~x1 & (x2 ? (x3 ? (~x4 & x5) : (x4 & ~x5)) : (x4 & (x5 ? ~x3 : x0)));
  assign z207 = (~x2 & ~n2804) | (~x3 & ~n2807) | ~n2810 | (x2 & ~n2808);
  assign n2804 = (x1 | n2806) & (n2805 | ((~x6 | x7 | ~x1 | x4) & (x1 | (x4 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n2805 = x0 ? (~x3 | x5) : (x3 | ~x5);
  assign n2806 = (x6 | ((x0 | x5 | (x3 ? (~x4 | x7) : (x4 | ~x7))) & (~x0 | ~x3 | x4 | ~x5 | ~x7))) & (~x0 | ~x5 | ~x6 | x7 | (~x3 ^ ~x4));
  assign n2807 = (x2 | (x4 ? ((x0 | x5 | x6) & (~x6 | (~x0 ^ (x1 & x5)))) : (~x5 | x6 | (~x0 & ~x1)))) & (x5 | ~x6 | x1 | ~x2) & (x0 | ((~x2 | x5 | ~x6) & (x1 | x4 | ((x5 | ~x6) & (~x2 | ~x5 | x6)))));
  assign n2808 = (~n586 | ~n1166) & (n857 | n2809);
  assign n2809 = (x5 | x6 | x7 | ~x3 | ~x4) & (x3 | ~x5 | (x4 ? (~x6 | ~x7) : (x6 | x7)));
  assign n2810 = (~n616 | n2813) & (~x3 | n2811) & (x2 | n2812);
  assign n2811 = (x2 & (x0 ? x1 : (x5 & ~x6))) | (x1 & (x5 ? x0 : x4)) | (~x5 & (x6 | (~x2 & x4) | (x0 & (x4 | (~x1 & ~x2))))) | (~x4 & x5 & ~x6) | (~x2 & x4 & x6);
  assign n2812 = (x0 | ~x3 | ~x5 | (x4 ? (~x6 | x7) : (x6 | ~x7))) & (x3 | ((x5 | ~x6 | x7 | x0 | ~x4) & (~x0 | ((~x6 | ~x7 | x4 | x5) & (x6 | x7 | ~x4 | ~x5)))));
  assign n2813 = (x3 | ~x4 | x5 | x6 | ~x7) & (~x3 | ((x4 | x5 | ~x6 | x7) & (x6 | ~x7 | ~x4 | ~x5)));
  assign z208 = n2815 | ~n2820 | (~n662 & ~n2819) | (n539 & ~n2818);
  assign n2815 = ~x1 & (x0 ? ~n2817 : ~n2816);
  assign n2816 = (x2 | x3 | x4 | x5 | ~x6 | ~x7) & ((x4 ? (x6 | ~x7) : (~x6 | x7)) | (x2 ? (~x3 | x5) : (x3 | ~x5)));
  assign n2817 = (~x4 | ((x2 | x3 | ~x5 | x6 | x7) & (~x6 | (x2 ? (x3 ? (~x5 | ~x7) : (x5 | x7)) : (~x3 | x7))))) & (x3 | x4 | ((x6 | x7 | ~x2 | x5) & (x2 | (x5 ? (x6 | ~x7) : (~x6 | x7)))));
  assign n2818 = (x0 | ~x3 | ~x4 | ~x6 | (~x5 ^ x7)) & (x3 | x6 | ~x7 | (x5 ? x4 : ~x0));
  assign n2819 = (x2 | ((~x0 | (x1 ? (x3 | ~x4) : (~x3 | x4))) & (~x3 | x4 | (x1 ? x0 : ~x5)))) & (x0 | ((x1 | (x3 ? (~x4 | x5) : (x4 | ~x5))) & (~x2 | ((x3 | x4 | ~x5) & (~x4 | (~x3 & x5)))))) & (x1 | ((x4 | ~x5 | ~x0 | ~x3) & (~x2 | ((~x4 | x5) & (x3 | x4 | ~x5)))));
  assign n2820 = ~n2822 & ~n2823 & ~n2824 & n2826 & (x0 | n2821);
  assign n2821 = (x1 | ~x2 | x3 | ~x4 | ~x5 | ~x6) & (x4 | ((x1 | x2 | ~x3 | x5 | x6) & (~x1 | ((x2 | x3 | ~x6) & (~x5 | x6 | ~x2 | ~x3)))));
  assign n2822 = ~n1099 & ((n1843 & ~n2008) | (n1176 & n768));
  assign n2823 = ~n857 & ((n2326 & n768) | (x2 & ~n856));
  assign n2824 = ~x7 & n2825 & ((~n1130 & ~n1243) | (n2095 & n598));
  assign n2825 = ~x2 & x6;
  assign n2826 = x1 | (x0 ? (x2 | ~n2112) : (~x2 | ~n1810));
  assign z209 = ~n2830 | ~n2834 | (~x1 & (x3 | ~n2829) & (~x3 | ~n2828));
  assign n2828 = (x5 | ((~x0 | ~x2 | x4 | x6 | x7) & (~x6 | ((x0 | x2 | ~x4 | ~x7) & (x7 | (x0 ? (~x2 ^ ~x4) : (~x2 | x4))))))) & (~x0 | x4 | ~x5 | x6 | (x2 ^ x7));
  assign n2829 = x2 ? ((x0 | x4 | x6 | (x5 ^ x7)) & (~x4 | ~x6 | (x0 ? (~x5 ^ x7) : (x5 | x7)))) : ((x0 | x5 | (x4 ? (x6 | ~x7) : (~x6 | x7))) & (~x5 | ((x4 | x6 | x7) & (~x0 | ~x4 | ~x6 | ~x7))));
  assign n2830 = (x0 | n2833) & (n620 | n2832) & (x2 | n2831);
  assign n2831 = (x0 | ~x3 | ~x5 | x7 | (x1 ^ x4)) & (x5 | ((x3 | ((x4 | ~x7 | x0 | ~x1) & (~x0 | (x1 ? (x4 | x7) : (~x4 | ~x7))))) & (x0 | ~x3 | ~x7 | (x1 ^ x4))));
  assign n2832 = (~x3 | ~x4 | x5 | x0 | x1 | ~x2) & (x2 | ((~x3 | ((x0 | (x1 ? (x4 | x5) : (~x4 | ~x5))) & (~x4 | x5 | ~x0 | x1))) & (~x0 | x3 | x5 | (x1 ^ x4))));
  assign n2833 = (x3 | ((~x1 | ~x2 | x4 | x5 | x6) & (~x4 | ~x5 | ~x6 | x1 | x2))) & (~x4 | x5 | x6 | x1 | x2 | ~x3) & (~x5 | (x1 ? ((x2 | x4 | ~x6) & (~x4 | x6 | ~x2 | ~x3)) : (~x2 | ~x3 | (x4 ^ x6))));
  assign n2834 = ~n2835 & ~n2839 & (~x2 | n2837) & (~x0 | n2838);
  assign n2835 = x1 & ((n2314 & n698) | (~x0 & ~n2836));
  assign n2836 = (~x4 | ((~x5 | x6 | ~x7 | ~x2 | x3) & (~x6 | ((x5 | ~x7 | ~x2 | x3) & ((x5 ^ x7) | (~x2 ^ ~x3)))))) & (~x5 | x7 | ((~x2 | x3 | x4 | ~x6) & (x2 | x6 | (x3 & x4))));
  assign n2837 = (x4 | (x0 ? (x1 | x3 | (~x5 ^ x7)) : (~x1 | ~x3 | (x5 ^ x7)))) & (x1 | ~x4 | ~x5 | ~x7 | (x0 ^ x3));
  assign n2838 = (x1 | ~x2 | x3 | ~x4 | x5 | x6) & (x2 | ~x5 | ((~x4 | ~x6 | x1 | ~x3) & (x3 | (x1 ? (x4 ^ x6) : (~x4 ^ x6)))));
  assign n2839 = ~n1862 & (x2 ? ((x3 & ~x5 & x0 & ~x1) | (~x0 & ((~x3 & ~x5) | (~x1 & x3 & x5)))) : (x5 & (x0 ? (x1 ^ x3) : (~x1 & ~x3))));
  assign z210 = n2846 | ~n2847 | (~x5 & ~n2841) | (~n620 & ~n2845);
  assign n2841 = (n2842 | n2844) & (~x0 | ~n670 | ~n2288) & (x0 | n2843);
  assign n2842 = x0 ? (x1 | ~x4) : (~x1 | x4);
  assign n2843 = (x1 | ~x2 | ~x3 | x4 | x6 | x7) & (~x4 | ((x1 | ((x2 | x6 | x7) & (~x2 | x3 | ~x6 | ~x7))) & (x6 | x7 | ((x2 | x3) & (~x1 | ~x2 | ~x3)))));
  assign n2844 = (x2 | x3 | ~x6 | ~x7) & (~x2 | (x3 ? (~x6 | ~x7) : (x6 | x7)));
  assign n2845 = ((~x0 ^ x2) | (x1 ? (x3 ? (x4 | x5) : (~x4 | ~x5)) : (~x5 | (~x3 ^ ~x4)))) & (x1 | ((~x0 | ~x2 | ~x3 | (~x4 ^ x5)) & (x3 | ~x4 | ((x2 | x5) & (x0 | (x2 & x5)))))) & (x0 | ~x1 | x2 | x4 | (x3 ^ x5));
  assign n2846 = ~n1215 & (x1 ? ((~x3 & ~x4 & x0 & ~x2) | (~x0 & (x2 ? (x3 ^ ~x4) : (~x3 & x4)))) : (x0 ? (x2 ? (~x3 & x4) : (x3 & ~x4)) : (x2 ? (x3 & ~x4) : (x3 ^ ~x4))));
  assign n2847 = (x0 | n2849) & (x6 | ~n2573 | n2850) & (~x0 | n2848);
  assign n2848 = (~x1 | x2 | x3 | ~x4 | x5 | x6) & (x1 | (((~x2 ^ ~x3) | (x4 ? (~x5 | ~x6) : (x5 | x6))) & (x4 | ~x6 | ~x2 | x3) & (x2 | ~x3 | ~x4 | x5 | x6)));
  assign n2849 = x1 ? (x2 ? ((x3 | ~x4 | x5 | x6) & (~x5 | ~x6 | ~x3 | x4)) : ((~x5 | ~x6 | x3 | x4) & (~x3 | (x4 ? ~x6 : (x5 | x6))))) : ((~x2 | x3 | (x4 ? (~x5 | ~x6) : (x5 | x6))) & (~x3 | ((x2 | x4 | ~x6) & (x5 | x6 | ~x2 | ~x4))));
  assign n2850 = (x1 | ~x3 | ~x7 | (~x0 ^ x4)) & (x3 | (~x0 ^ x7) | (x1 ^ x4));
  assign z211 = (x2 | ~n2852 | ~n2859) & (~n2857 | ~n2860 | ~x2 | n2856);
  assign n2852 = (x3 | (n2853 & (~x6 | n2854))) & (x6 | ((~n1317 | n2855) & (~x3 | n2854)));
  assign n2853 = (~x4 | (x0 ? (~x5 | (x1 ? (~x6 | x7) : (x6 | ~x7))) : (x1 | x5 | (~x6 ^ x7)))) & (~x1 | x4 | ((x6 | ~x7 | x0 | ~x5) & (~x0 | ~x6 | (x5 ^ x7))));
  assign n2854 = (x0 | ~x1 | x4 | x5 | ~x7) & (x1 | ((x5 | x7 | x0 | x4) & (~x0 | (x4 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n2855 = (x1 | x4 | ~x5 | ~x7) & (~x4 | (x1 ? (~x5 ^ ~x7) : (~x5 | x7)));
  assign n2856 = ~n662 & (((x3 ^ x5) & (x0 ? (~x1 & x4) : (x1 & ~x4))) | (~x0 & ~x1 & (x3 ? (~x4 & x5) : (x4 & ~x5))));
  assign n2857 = (~n559 | ~n586) & (x0 | ~x7 | n2858);
  assign n2858 = (x1 | x3 | x4 | x5 | x6) & (~x4 | ~x5 | ~x6 | ~x1 | ~x3);
  assign n2859 = ((~x0 ^ x3) | (x1 ? (x4 ? (x5 | ~x7) : (~x5 | x7)) : (x5 | (~x4 ^ x7)))) & (x0 | ((~x4 | ~x5 | ~x7 | x1 | ~x3) & (x3 | (x1 ? ((~x4 | ~x5 | ~x7) & (x5 | x7)) : (~x5 | (~x4 ^ x7)))))) & (~x0 | ~x3 | ((x4 | x5 | x7) & (x1 | ~x5 | (~x4 ^ x7))));
  assign n2860 = ((x4 ^ x7) | ((x0 | ~x1 | x3 | x5) & (x1 | (x0 ? (~x3 | ~x5) : (~x3 ^ x5))))) & (~x0 | x1 | ((x4 | x5 | ~x7) & (x3 | (x4 ? (x5 | x7) : ~x7)))) & (x0 | ((~x5 | x7 | ~x3 | ~x4) & (~x1 | ((~x4 | ~x5 | x7) & (~x3 | (x4 ? x7 : (~x5 | ~x7)))))));
  assign z212 = ~n2866 | (x0 ? ~n2864 : (x1 ? ~n2862 : ~n2863));
  assign n2862 = x2 ? (~x3 | x7 | (x4 ? x5 : (~x5 | x6))) : (~x6 | ~x7 | (x5 ? x3 : x4));
  assign n2863 = (~x5 | ((x2 | ((x3 | x4 | ~x6 | x7) & (x6 | ~x7 | ~x3 | ~x4))) & (~x4 | ((x3 | x6 | x7) & (~x6 | ~x7 | ~x2 | ~x3))))) & (~x2 | x4 | x5 | ~x6 | (x3 ^ ~x7));
  assign n2864 = x1 ? (~n563 | ~n1163) : n2865;
  assign n2865 = (x3 | ((~x4 | ((~x6 | x7 | ~x2 | x5) & (x2 | ((~x6 | ~x7) & (~x5 | x6 | x7))))) & (~x2 | x4 | x6 | (~x5 ^ x7)))) & (x2 | ~x7 | (x4 ? (x5 | ~x6) : (~x5 | x6)));
  assign n2866 = (x2 | n2869) & (n846 | n2868) & (~x2 | n2867);
  assign n2867 = (x0 | (x1 ? ((x3 | ~x4 | ~x5 | x6) & (x5 | ~x6 | ~x3 | x4)) : (x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))))) & (x1 | ((~x0 | x3 | x4 | x5 | ~x6) & (~x3 | ((~x4 | ~x5 | x6) & (~x0 | ((~x5 | x6) & (~x4 | x5 | ~x6)))))));
  assign n2868 = (x1 | ((~x0 | (x2 ? (x3 | ~x4) : x4)) & (~x3 | ((~x2 | x4 | x7) & (x0 | (~x4 ^ x7)))))) & (x0 | ((x3 | x4 | ~x1 | ~x2) & (~x4 | ((~x1 | (x3 ^ x7)) & (x2 | ~x3 | ~x7))))) & (~x1 | x2 | x3 | (x7 ? ~x0 : ~x4));
  assign n2869 = x0 ? ((~x1 | x3 | x4 | x5 | ~x6) & (x1 | ~x3 | ~x4 | ~x5 | x6)) : (x5 ? (x6 | ((x3 | x4) & (~x1 | (x3 & x4)))) : (~x6 | (x1 ? (~x3 | ~x4) : (~x3 ^ x4))));
  assign z213 = n2873 | ~n2876 | (x2 ? ~n2872 : ~n2871);
  assign n2871 = x0 ? ((~x4 | ~x5 | ~x6 | x1 | ~x3) & (x5 | (x1 ? (x3 ? (x4 | x6) : (~x4 | ~x6)) : (~x4 | x6)))) : ((x5 | ~x6 | x1 | ~x4) & (~x5 | ((x1 | x3 | x4 | x6) & (~x1 | ((x3 | x4 | ~x6) & (~x4 | x6))))));
  assign n2872 = (x1 | ((~x3 | ((~x5 | x6 | x0 | ~x4) & (~x0 | (x4 ? (x5 | ~x6) : (~x5 | x6))))) & (x0 | x4 | ((~x5 | ~x6) & (x3 | x5 | x6))))) & (x0 | ~x1 | x5 | ((x4 | ~x6) & (~x3 | ~x4 | x6)));
  assign n2873 = x2 & ((n738 & ~n2875) | (~x0 & ~n2874));
  assign n2874 = (x1 | ~x3 | x4 | ~x5 | x6 | x7) & (~x1 | ~x4 | ((~x6 | ~x7 | ~x3 | x5) & (x6 | x7 | x3 | ~x5)));
  assign n2875 = (~x3 | x4 | x5 | ~x6 | x7) & (x3 | ~x5 | (x4 ? (~x6 | x7) : (x6 | ~x7)));
  assign n2876 = (~x4 | (x7 ? n2877 : n2878)) & (~x7 | ~n670 | n2879) & (x4 | (x7 ? n2878 : n2877));
  assign n2877 = x5 ? ((~x0 | ~x1 | x2 | x3 | x6) & (x0 | (x1 ? (~x6 | (~x2 & ~x3)) : (x6 | (~x2 ^ x3))))) : ((~x2 | ~x3 | x6 | x0 | x1) & ((x2 & x3) | (x0 ? (x1 | ~x6) : (~x1 | x6))));
  assign n2878 = x5 ? (x0 ? ((x3 | ~x6 | ~x1 | x2) & (x1 | (x2 ? (~x3 | ~x6) : x6))) : ((x1 | x2 | ~x6) & (~x3 | x6 | ~x1 | ~x2))) : ((x6 | ((x0 | x1 | x2 | x3) & (~x0 | (x1 ? (x2 | x3) : ~x2)))) & (x0 | ~x6 | (x1 ^ ~x2)));
  assign n2879 = (~x4 | ~x5 | ~x6 | ~x0 | x3) & (x0 | x6 | (x3 ? (x4 | x5) : (~x4 | ~x5)));
  assign z214 = n2882 | n2885 | ~n2886 | ~n2887 | (n539 & ~n2881);
  assign n2881 = (x5 | ~x6 | x7 | ~x0 | x3 | ~x4) & (x0 | (x3 ? (~x5 | (x4 ? (x6 | x7) : (~x6 | ~x7))) : (x5 | x6 | (~x4 ^ x7))));
  assign n2882 = ~x1 & (x6 ? ~n2883 : (n2326 & ~n2884));
  assign n2883 = (x4 | ~x5 | x7 | ~x0 | x2 | ~x3) & ((x2 ? (x3 | ~x5) : (~x3 | x5)) | (x0 ? (~x4 | ~x7) : (x4 | x7)));
  assign n2884 = (~x0 | x3 | x5 | x7) & (x0 | ~x7 | (~x3 ^ ~x5));
  assign n2885 = ~n1099 & ((x0 & ~x1 & x2 & x5 & ~x7) | (~x0 & x7 & (x1 ? (x2 ^ ~x5) : (~x2 & x5))));
  assign n2886 = (x3 | ((x0 | ~x1 | x2 | ~x5 | x7) & (~x0 | ~x7 | (x1 ? (x2 | ~x5) : (~x2 | x5))))) & (x0 | ~x2 | ~x3 | x5 | (x1 ^ ~x7));
  assign n2887 = (~x5 | (x6 ? n2888 : n2890)) & (x7 | n2889) & (x5 | (x6 ? n2890 : n2888));
  assign n2888 = x0 ? (x1 | (x3 ? (x2 ? ~x7 : (~x4 | x7)) : (x4 | x7))) : ((~x7 | ((x1 | x2 | x3 | x4) & (~x1 | (x2 ? (x3 | x4) : (~x3 | ~x4))))) & (x1 | ~x2 | x7 | (~x3 ^ x4)));
  assign n2889 = (~x3 | x4 | x5 | ~x0 | x2) & (x0 | ((~x1 | x2 | ~x3 | x4 | ~x5) & (x1 | ((x2 | ~x3 | ~x4 | x5) & (~x2 | (x3 ? (~x4 | ~x5) : (x4 | x5)))))));
  assign n2890 = x2 ? ((~x0 | x1 | ~x3 | ~x4 | x7) & (x0 | (x1 ? (x3 ? (~x4 | ~x7) : x7) : (x3 | ~x7)))) : ((x0 | x1 | x3 | x7) & (~x0 | ((x4 | x7 | ~x1 | x3) & (x1 | ~x7 | (x3 & x4)))));
  assign z216 = ~n2896 | (~x0 & ~n2892) | (~x3 & (n2893 | n2894));
  assign n2892 = (x2 | ((x1 | x3 | ~x4 | x5 | x7) & (~x1 | ~x3 | x4 | ~x5 | ~x7))) & (~x1 | ((x5 | ~x7 | ~x3 | ~x4) & (~x2 | (x4 ^ x7) | (~x3 & x5))));
  assign n2893 = ~n927 & (x1 ? (~x6 & ((~x2 & ~x5) | (~x0 & x2 & x5))) : (x6 & (x2 ^ ~x5)));
  assign n2894 = n543 & n2512 & (x0 ? n2895 : n1184);
  assign n2895 = x2 & x5;
  assign n2896 = n594 & ~n2898 & (n989 | n2897) & (~n568 | ~n2609);
  assign n2897 = (~x0 | x2 | x3 | ~x4 | x5 | x7) & (x0 | ~x5 | ((x4 | ~x7 | ~x2 | x3) & (~x4 | x7 | x2 | ~x3)));
  assign n2898 = (x4 ^ x7) & ((x1 & ~x2 & ~x3 & x5) | (~x1 & ((x3 & ~x5) | (x2 & (x3 | ~x5)))));
  assign z217 = n2900 | ~n2904 | (~n607 & ~n2903);
  assign n2900 = ~x1 & (x0 ? ~n2902 : ~n2901);
  assign n2901 = x3 ? ((~x5 | x6 | ~x7 | x2 | ~x4) & (x5 | ~x6 | x7 | ~x2 | x4)) : (x2 ? ((x6 | x7 | x4 | x5) & (~x6 | ~x7 | ~x4 | ~x5)) : (~x4 | ~x6 | (~x5 ^ x7)));
  assign n2902 = (x2 | ~x3 | ~x4 | x5 | x6 | x7) & (x3 | ((x2 | x4 | x5 | x6 | ~x7) & (~x2 | ~x4 | ~x6 | (x5 ^ x7))));
  assign n2903 = (x0 | ~x1 | x3 | x4 | x5 | x6) & (~x4 | ((x0 | ~x1 | (x3 ? (~x5 | x6) : (x5 | ~x6))) & (~x0 | x1 | ~x3 | ~x5 | x6)));
  assign n2904 = (~n2747 | n2907) & (x2 | n2905) & (~x2 | n2906);
  assign n2905 = (x4 & ((x3 & ~x6) | (~x0 & ~x5))) | (~x3 & ((~x0 & ((x5 & x6) | (x1 & ~x4 & ~x6))) | (x5 & x6 & (x1 | ~x4)))) | (~x5 & ~x6) | (x3 & (~x5 | (x0 & x1)));
  assign n2906 = (x5 & (x3 | x4 | ~x6)) | (x0 & x1) | (~x3 & ~x5 & x6) | (~x0 & ~x4 & ((~x3 & ~x6) | (~x1 & ~x5 & x6)));
  assign n2907 = (~x0 | x2 | x4 | x5 | x6 | ~x7) & (~x5 | ((~x6 | x7 | x2 | ~x4) & (x0 | ((~x6 | ~x7 | ~x2 | ~x4) & (x2 | x4 | x6 | x7)))));
  assign z218 = n2909 | n2912 | ~n2914 | (x1 ? ~n2913 : ~n2911);
  assign n2909 = ~x0 & (x1 ? ~n2910 : (~n633 | (n563 & n1382)));
  assign n2910 = (x5 | x7 | ((~x3 | (x2 ? (x4 | x6) : (~x4 | ~x6))) & (x2 | x3 | (~x4 ^ x6)))) & (x3 | ~x7 | ((~x4 | ~x6) & (~x5 | x6 | x2 | x4)));
  assign n2911 = (~x6 | ((~x3 | ~x4 | ~x5 | ~x0 | x2) & (x3 | ((~x0 | (x2 ? x4 : (~x4 | x5))) & (x4 | ~x5) & (x0 | (x2 ? (~x4 | x5) : x4)))))) & (~x3 | x6 | ((x0 | (x5 ? ~x2 : ~x4)) & (x4 | (~x0 & ~x5)) & (~x2 | ~x4 | x5)));
  assign n2912 = ~n622 & ((x1 & ~x2 & ~x3 & ~x6) | (~x0 & ((x1 & ~x3 & ~x6) | (~x1 & x2 & x3 & x6))));
  assign n2913 = (x4 | ((x2 | x3 | ~x5 | ~x6) & (x0 | ((~x2 | x3 | ~x6) & (~x3 | ~x5 | x6))))) & (x5 | ((x3 | ~x6 | ~x0 | x2) & (x0 | ~x3 | x6 | (x2 & ~x4))));
  assign n2914 = (n620 | n2915) & (~x0 | (~n2917 & (x2 | n2916)));
  assign n2915 = (x1 | ((~x2 | ((~x4 | ~x5 | ~x0 | ~x3) & (x4 | x5 | x0 | x3))) & (~x0 | x2 | x5 | (~x3 ^ ~x4)))) & (x0 | ~x3 | ~x4 | ~x5 | (~x1 & x2));
  assign n2916 = (~x1 | ((~x3 | x4 | x5 | x6 | x7) & (~x5 | ~x6 | ~x7 | x3 | ~x4))) & (~x5 | x6 | ~x7 | x1 | ~x3 | ~x4);
  assign n2917 = x4 & n538 & ((n544 & n1343) | (~x3 & ~n662));
  assign z219 = ~n2921 | ~n2925 | (~n1041 & ~n2919) | (~x2 & ~n2920);
  assign n2919 = (x0 | ~x1 | ~x2 | x3 | x5 | x7) & (x1 | ((x0 | x2 | x3 | x5 | x7) & (~x3 | ((~x5 | x7 | x0 | ~x2) & (~x0 | (x2 ? (x5 | x7) : (~x5 | ~x7)))))));
  assign n2920 = (x4 | ~x5 | x7 | ~x0 | x1) & (x3 | (x0 ? (x1 | (x4 ? x7 : (x5 | ~x7))) : (~x1 | ~x7 | (~x4 & x5))));
  assign n2921 = ~n2924 & ((x4 & ~x7 & (x5 | n2923)) | (~x4 & (x7 | (~x5 & n2922))) | (n2922 & (n2923 | (~x5 & x7))));
  assign n2922 = x0 ? (x1 | (~x2 ^ (x3 & ~x5))) : ((x1 | x2 | x3 | ~x5) & (~x1 | (x2 ? (x3 | ~x5) : ~x3)));
  assign n2923 = (x0 | x1 | (~x2 ^ x3)) & (~x1 | (x0 ? (x2 | x3) : (~x2 | ~x3)));
  assign n2924 = ~x5 & n538 & ((x0 & x3 & x4 & x7) | (~x0 & ((~x4 & x7) | (x3 & x4 & ~x7))));
  assign n2925 = x0 ? (x2 | n2928) : (~n2927 & (~x4 | n2926));
  assign n2926 = (x5 | ((~x6 | ~x7 | x1 | x2) & (~x1 | ((~x2 | x3 | ~x6 | ~x7) & (x6 | x7 | x2 | ~x3))))) & (x1 | ~x2 | ~x5 | (x3 ? (~x6 | ~x7) : (x6 | x7)));
  assign n2927 = x7 & n642 & ((x3 & ~x5 & ~x1 & ~x2) | (x1 & (x2 ? ~x5 : (~x3 & x5))));
  assign n2928 = (~x1 | x4 | x5 | x6 | ~x7) & (x3 | ((~x5 | x6 | ~x7 | x1 | ~x4) & (~x1 | x5 | ~x6 | (~x4 ^ ~x7))));
  assign z220 = ~n2932 | (~x2 & ((x4 & ~n2930) | (x3 & ~x4 & ~n2931)));
  assign n2930 = x0 ? ((~x1 | x3 | ~x5 | ~x6 | ~x7) & (x1 | ((x6 | ~x7 | x3 | x5) & (~x3 | ~x6 | (~x5 ^ x7))))) : (~x3 | ((~x1 | x6 | (x5 ^ x7)) & (~x6 | x7 | x1 | x5)));
  assign n2931 = (~x0 | x1 | ~x5 | ~x6 | x7) & (x0 | ((x6 | ~x7 | ~x1 | ~x5) & (x1 | ~x6 | (x5 ^ x7))));
  assign n2932 = n2934 & ~n2939 & (~n871 | n2933) & (x0 | n2938);
  assign n2933 = (x0 | ~x1 | x4 | x5 | ~x6 | x7) & (x1 | x6 | ((x5 | ~x7 | x0 | x4) & (~x0 | ((x5 | x7) & (x4 | ~x5 | ~x7)))));
  assign n2934 = ~n2935 & ~n2936 & (n1099 | n2937);
  assign n2935 = ~x1 & (((~x0 ^ x5) & (x2 ^ (x3 & ~x6))) | (~x2 & ~x3 & x6 & (x0 ^ x5)));
  assign n2936 = x1 & ((~x5 & ~x6 & ~x0 & x2) | (~x2 & ((~x5 & ~x6 & x0 & ~x3) | (~x0 & x5 & (~x3 | x6)))));
  assign n2937 = (x5 | ~x6 | x7 | ~x0 | ~x1 | x2) & (x0 | ~x2 | ~x5 | (x1 ? (~x6 | ~x7) : (x6 | x7)));
  assign n2938 = (~x4 | ((x1 | x6 | (x2 ? (~x3 | ~x5) : (x3 | x5))) & (~x1 | ~x2 | ~x3 | x5 | ~x6))) & (~x1 | x3 | x4 | ~x6 | (x2 ^ x5));
  assign n2939 = n651 & ((~x1 & ~x3 & x4 & x5 & ~x6) | (~x4 & (x1 ? (x3 ? (~x5 & ~x6) : (x5 & x6)) : (~x5 & (~x3 ^ x6)))));
  assign z221 = ~n2942 | ~n2946 | (~n620 & ~n2941);
  assign n2941 = x1 ? ((x2 | ((x4 | ~x5 | x0 | x3) & (~x0 | (x3 ? (x4 | x5) : ~x4)))) & (x0 | ~x2 | (x3 ? x4 : (~x4 | ~x5)))) : (x2 | ~x3 | (x5 ? (~x0 & x4) : (x0 & ~x4)));
  assign n2942 = (~n975 | n2945) & (~x1 | n2944) & (n662 | n2943);
  assign n2943 = (x1 | ((~x0 | ((~x2 | ~x3 | x4) & (~x4 | x5 | x2 | x3))) & (~x2 | ((~x3 | x4 | x5) & (~x4 | ~x5 | x0 | x3))))) & (x0 | ~x1 | x2 | ~x3 | (~x4 ^ x5));
  assign n2944 = (x0 | ((~x4 | ~x6 | (~x2 ^ ~x3)) & (~x2 | x3 | x6 | (x4 & x5)))) & (x2 | x3 | x4 | x6 | (~x0 & x5));
  assign n2945 = (x3 | x4 | ~x5 | ~x6 | ~x7) & (~x3 | ((x4 | x5 | ~x6 | ~x7) & (x6 | x7 | ~x4 | ~x5)));
  assign n2946 = x1 | ((~n1415 | ~n565) & n2947 & (~x2 | n2948));
  assign n2947 = x3 ? ((~x0 | x2 | x4 | x5 | x6) & (~x4 | ((~x2 | ~x5 | x6) & (x0 | (x2 ? x6 : (~x5 | ~x6)))))) : ((~x6 | ((~x2 | x4) & (~x0 | x5 | (~x2 & x4)))) & (x2 | x6 | ((~x4 | ~x5) & (x0 | (~x4 & ~x5)))));
  assign n2948 = (x0 | ~x3 | x4 | ~x5 | x6 | x7) & (~x4 | ((x0 | x3 | x5 | ~x6 | ~x7) & (~x0 | ((~x6 | ~x7 | x3 | ~x5) & (x6 | x7 | ~x3 | x5)))));
  assign z222 = ~n2950 | (x1 & ~n2956) | (~x3 & (~n2958 | (~x1 & ~n2957)));
  assign n2950 = ~n2951 & n2955 & (~x3 | (~n2953 & (~n2014 | n2954)));
  assign n2951 = ~x1 & ~n2952;
  assign n2952 = x4 ? (x7 ? ((~x0 | x2 | x3 | ~x5) & ((~x0 ^ ~x2) | (x3 ^ x5))) : ((~x0 | x2 | x3 | x5) & (x0 | (x2 ? (x3 | ~x5) : (~x3 | x5))))) : ((x0 | ~x2 | ~x3 | x5 | x7) & (x2 | ((~x5 | ~x7 | x0 | x3) & (~x0 | (x3 ? (~x5 | x7) : (x5 | ~x7))))));
  assign n2953 = ~n662 & ((x0 & ~x1 & x2 & x4 & ~x5) | (~x0 & x5 & (x1 ? (~x2 & x4) : (x2 & ~x4))));
  assign n2954 = (~x6 | x7 | x0 | ~x1) & (x6 | ~x7 | ~x0 | x1);
  assign n2955 = x3 ? ((~x4 | ~x7 | x0 | ~x2) & (x7 | ((x0 | ~x1 | ~x2 | x4) & (x1 | (x0 ? (~x2 ^ x4) : (x2 | x4)))))) : ((~x0 | ~x1 | x2 | ~x4 | x7) & (~x7 | ((x1 | ~x2 | x4) & (x0 | ((~x2 | x4) & (~x1 | x2 | ~x4))))));
  assign n2956 = (x0 | ~x2 | x3 | ~x4 | ~x5 | x7) & (x2 | ((x0 | ~x3 | ~x4 | x5 | x7) & (x4 | (x0 ? (x5 | (~x3 ^ x7)) : (~x5 | x7)))));
  assign n2957 = (x0 | x2 | x4 | x5 | ~x6 | ~x7) & (~x4 | ~x5 | ((x6 | ~x7 | x0 | x2) & (~x0 | x7 | (x2 ^ x6))));
  assign n2958 = (~x1 | x6 | ~x7 | n2959) & (~x6 | ((~x7 | ~n1449 | ~n924) & (x1 | x7 | n2959)));
  assign n2959 = (x4 | ~x5 | ~x0 | x2) & (x0 | x5 | (~x2 ^ ~x4));
  assign z223 = x2 ? ~n1864 : (~n1859 | ~n1861 | (~x5 & ~n2961));
  assign n2961 = (~x4 | (x0 ? (x1 | (x3 ? (x6 | ~x7) : (~x6 | x7))) : (~x1 | x3 | (~x6 ^ x7)))) & (x0 | ~x1 | ~x3 | x4 | x6 | ~x7);
  assign z224 = n1877 | ~n2963 | (~x2 & ~n2967) | (~x1 & ~n2968);
  assign n2963 = ~n2966 & ~n2964 & (~n738 | n2354 | x6 | ~n2327);
  assign n2964 = ~n824 & ~n2965;
  assign n2965 = ((~x4 ^ x6) | (x0 ? (x3 | (x1 ^ ~x2)) : (x1 | ~x3))) & (~x0 | x1 | x2 | x3 | x4 | x6) & (x0 | ((~x4 | ~x6 | x1 | x3) & (~x1 | ((~x3 | ~x4 | ~x6) & (x4 | x6 | ~x2 | x3)))));
  assign n2966 = ~n1115 & ((x4 & x6 & x0 & ~x1) | (~x0 & (x1 ? ((x4 & ~x6) | (x2 & ~x4 & x6)) : (~x4 & ~x6))));
  assign n2967 = (x4 | ((~x0 | x1 | ~x5 | (~x3 ^ x6)) & (~x1 | ((x5 | x6 | ~x0 | x3) & (x0 | (x3 ? (x5 | ~x6) : (~x5 | x6))))))) & (~x0 | x3 | ~x4 | ~x5 | (x1 ^ x6));
  assign n2968 = (~x0 | n1876) & (n1875 | ((~x2 | ~x4 | x6) & (x0 | (~x4 & ~x6))));
  assign z225 = n1883 | ~n2971 | (~n592 & ~n2970) | (~x2 & n1881);
  assign n2970 = ((~x2 & ~x3) | (x0 ? (x1 | ~x6) : (~x1 | x6))) & (x5 | ~x6 | x0 | x1) & (~x0 | x2 | x3 | (x1 ? ~x6 : (x5 | x6)));
  assign n2971 = ~n1889 & (~n664 | ~n957) & (~n1886 | ~n1887);
  assign z226 = n1896 | n2974 | n2976 | ~n2977 | (x0 & ~n2973);
  assign n2973 = (~x7 | n933 | x5 | ~x6) & (x6 | ((~x4 | ~n1386 | (x5 ^ x7)) & (~x5 | ~x7 | n933)));
  assign n2974 = ~n846 & ~n2975;
  assign n2975 = (x1 | ((x3 | x4 | x7 | ~x0 | x2) & (x0 | ~x7))) & (x0 | ~x1 | x7 | (~x2 & ~x3 & ~x4));
  assign n2976 = ~x2 & ~x5 & ((x0 & ~x1 & (x3 ^ x7)) | (x1 & (x0 ? (~x3 & ~x7) : (x3 & x7))));
  assign n2977 = ~n2978 & (~x2 | ~n738 | ~n691) & (~n698 | ~n2473);
  assign n2978 = ~x0 & ((~x5 & x7 & x1 & x2) | (~x1 & x5 & ~x7));
  assign z227 = ~n2980 | (~x2 & (n1900 | (~x4 & n732 & ~n1351)));
  assign n2980 = x6 ? (x7 ? n2981 : n1906) : (x7 ? n1906 : n2981);
  assign n2981 = x1 ? (x2 | x3 | (~x0 & (x4 | x5))) : (~x2 & ~x3 & (x0 | (~x4 & ~x5)));
  assign z228 = x7 & (~n1799 | n720 | (n694 & n1112));
  assign z229 = ~n2986 | (n1977 & (x0 ? (~x2 & n2984) : (x2 & n2985)));
  assign n2984 = ~x6 & x3 & ~x4;
  assign n2985 = x6 & ~x3 & x4;
  assign n2986 = (~x0 & (~x1 | ~x2)) | (x1 & (x2 ? (x0 | (~x3 & ~n1701)) : (x3 & ~n686)));
  assign z230 = ~n2988 | (x3 & ((n872 & n1546) | (n651 & ~n1000)));
  assign n2988 = n2989 & (~n650 | ((~n768 | ~n1546) & (~n767 | ~n694)));
  assign n2989 = x1 ? ((x2 | (x0 & x3)) & (x0 | x3 | (x4 & ~n730))) : (~x2 | (~x0 & (~x3 | ~x4)));
  assign z231 = ~n2994 | ~n2991 | n2992;
  assign n2991 = x2 ? ((~x3 | ~x4 | ~x5 | ~x0 | x1) & (x0 | ((x3 | x4) & (x1 | (x3 & (x4 | x5)))))) : ((~x3 | (x0 ? (x1 | x5) : (~x1 & (~x4 | ~x5)))) & (~x0 | ((x1 | x4 | ~x5) & (x3 | (~x1 & ~x4)))));
  assign n2992 = x3 & ((~x5 & ~n2993) | (n1546 & n1846));
  assign n2993 = (~x4 | ~x6 | ~x7 | x0 | x1 | x2) & (~x0 | ((~x1 | x2 | x4 | ~x6 | x7) & (~x4 | x6 | ~x7 | x1 | ~x2)));
  assign n2994 = (x5 | n2995) & (~n587 | ~n2473) & (~n534 | ~n1478);
  assign n2995 = (x3 | ~x4 | x6 | x0 | ~x1 | ~x2) & (~x0 | ~x3 | ((~x4 | ~x6 | x1 | ~x2) & (~x1 | x2 | x4 | x6)));
  assign z232 = x2 ? (~n2997 | (x3 & ~n3002)) : (~n2998 | ~n2999);
  assign n2997 = (x0 | ((~x1 | (~x3 ^ ~x4)) & (x3 | ~x4 | (x1 & (x5 | x6))))) & (x1 | (x3 ? (x4 | (~x0 & x5)) : (~x4 | ~x5)));
  assign n2998 = x1 ? ((~x0 | ((x3 | ~x5 | ~x6) & (x5 | x6 | ~x3 | x4))) & (~x4 | ~x5 | ~x6 | x0 | ~x3) & (x3 | ((x0 | (~x5 ^ x6)) & (x4 | ~x5 | ~x6) & (~x4 | (x5 & x6))))) : ((x0 | ((~x5 | ~x6 | x3 | ~x4) & (~x3 | x5 | x6))) & (x4 | x5 | ~x0 | x3) & (~x3 | ((~x0 | (~x5 ^ x6)) & (~x4 | x5 | x6) & (x4 | (~x5 & ~x6)))));
  assign n2999 = (x4 | x5 | n3000 | ~x0 | ~x3) & (x0 | ~x4 | (x3 ? n3001 : (~x5 | n3000)));
  assign n3000 = x1 ? (~x6 | x7) : (x6 | ~x7);
  assign n3001 = (~x6 | x7 | x1 | x5) & (x6 | ~x7 | ~x1 | ~x5);
  assign n3002 = (~x0 | x1 | ~x4 | x5 | x6 | x7) & (x0 | x4 | ~x5 | (x1 ? (~x6 | ~x7) : (x6 | x7)));
  assign z233 = ~n3014 | n3013 | n3012 | n3009 | n3004 | n3006;
  assign n3004 = ~x1 & ~n3005;
  assign n3005 = (~x0 | ~x4 | x5 | (x2 ? (x3 | ~x6) : (~x3 | x6))) & (x4 | ((~x0 | x5 | (x2 ? (~x3 | ~x6) : x3)) & (~x2 | x3 | ~x5 | ~x6) & (x0 | ((~x2 | x3 | ~x6) & (~x5 | x6 | x2 | ~x3)))));
  assign n3006 = x2 & ((n664 & n3008) | (~x1 & ~n3007));
  assign n3007 = (~x5 | ~x6 | ~x7 | x0 | x3 | ~x4) & (x6 | (x0 ? ((x3 | x4 | ~x5 | ~x7) & (~x3 | ~x4 | x5 | x7)) : (x4 | (x3 ? (~x5 | x7) : (x5 | ~x7)))));
  assign n3008 = ~x4 & x6 & (x3 ? (x5 & ~x7) : (~x5 & x7));
  assign n3009 = ~x2 & ((n1122 & ~n3011) | (~x7 & ~n3010));
  assign n3010 = ((x1 ^ x6) | ((x0 | x3 | ~x4 | ~x5) & (~x0 | ~x3 | x4 | x5))) & (x0 | ~x3 | ~x4 | (x1 ? (~x5 | x6) : (x5 | ~x6)));
  assign n3011 = (x0 | x1 | x4 | ~x5 | ~x6) & (~x4 | ((x5 | x6 | x0 | ~x1) & (~x0 | (x1 ? (~x5 | x6) : (x5 | ~x6)))));
  assign n3012 = (n2327 | n2403) & ((x0 & ~x1 & x3 & x5) | (~x0 & ((x3 & ~x5) | (x1 & ~x3 & x5))));
  assign n3013 = n808 & ((~x0 & x3 & x5 & x6) | (x0 & ~x5 & (~x3 | ~x6)));
  assign n3014 = (n2322 | n3016) & (n3015 | (~n648 & (~x1 | n783)));
  assign n3015 = (x3 | ~x5 | ~x0 | x2) & (x0 | (x2 ? (~x3 | ~x5) : (x3 | x5)));
  assign n3016 = (x0 | (x1 ? (~x4 | x5) : (x4 | ~x5))) & (~x4 | x5 | ~x0 | x1);
  assign z234 = ~n3021 | (~x2 & ~n3024) | (~x3 & ~n3023) | (x2 & ~n3018);
  assign n3018 = (x1 | n3019) & (x0 | ~x1 | n3020);
  assign n3019 = ((x4 ? (~x6 | ~x7) : (x6 | x7)) | (x0 ? (x3 | ~x5) : (x3 ^ x5))) & (~x0 | ~x3 | ~x4 | x5 | x6 | x7) & (x0 | x3 | ~x5 | (x4 ? (~x6 | x7) : (x6 | ~x7)));
  assign n3020 = (~x3 | x4 | ~x5 | ~x6 | x7) & (x3 | ((x6 | ~x7 | ~x4 | ~x5) & (x4 | ~x6 | (x5 ^ x7))));
  assign n3021 = (~x3 | n3022) & (n850 | ((~x0 | ~x1 | x2 | x3) & (x0 | (x1 ? ~x3 : (x2 | x3)))));
  assign n3022 = (x6 | ((~x0 | x4 | x5 | (x1 ^ ~x2)) & (~x4 | (x0 ? (x1 | ~x5) : (x1 ? (~x2 | ~x5) : x5))))) & (x1 | ~x6 | ((x0 | x2 | ~x4 | ~x5) & ((~x2 & x4) | (x0 ^ x5))));
  assign n3023 = ((~x4 ^ x6) | (x0 ? (x1 | x5) : (~x5 | (x1 ^ ~x2)))) & (~x6 | ((~x2 | ~x4 | ~x5 | x0 | ~x1) & (~x0 | x1 | (x2 ? x5 : (~x4 | ~x5))))) & (x0 | ~x1 | x5 | x6 | (~x2 & x4));
  assign n3024 = x0 ? (x5 ? (x6 | n3026) : n3027) : (n3025 & (n3026 | (~x5 ^ ~x6)));
  assign n3025 = ((~x5 ^ x7) | ((~x1 | ~x3 | ~x4 | x6) & (x1 | x3 | x4 | ~x6))) & (x5 | ~x6 | ~x7 | ~x1 | ~x3 | x4) & (x1 | ~x4 | x7 | (x3 ? (x5 | ~x6) : (~x5 | x6)));
  assign n3026 = (~x4 | x7 | ~x1 | x3) & (x4 | ~x7 | x1 | ~x3);
  assign n3027 = (x1 | ~x4 | ~x6 | (x3 ^ x7)) & (x4 | (~x1 ^ ~x6) | (~x3 ^ x7));
  assign z235 = ~n3033 | (x7 ? (x2 ? ~n3029 : ~n3030) : ~n3031);
  assign n3029 = (~x3 | ((x1 | (x4 ^ x6) | (x0 ^ x5)) & (x0 | ~x1 | (x4 ? (~x5 | x6) : (x5 | ~x6))))) & (~x0 | x1 | x3 | ~x4 | (~x5 ^ x6));
  assign n3030 = (~x0 | x1 | x3 | x4 | ~x5 | ~x6) & (x6 | ((x0 | x1 | ~x3 | ~x4 | ~x5) & (x3 | ((x4 | ~x5 | x0 | x1) & (~x0 | (x4 ? x5 : ~x1))))));
  assign n3031 = x0 ? (~n538 | ~n1773) : n3032;
  assign n3032 = x1 ? (x2 | ((x3 | ~x4 | x5 | ~x6) & (~x3 | x4 | (~x5 ^ x6)))) : (x2 ? (x4 | (x3 ? (x5 | x6) : (~x5 | ~x6))) : (~x4 | (x3 ? (~x5 ^ x6) : (x5 | x6))));
  assign n3033 = ~n3036 & n3037 & (n662 | n3034) & (x2 | n3035);
  assign n3034 = x1 ? ((x3 | ~x4 | ~x0 | x2) & (x0 | ((x2 | ((~x4 | x5) & (x3 | x4 | ~x5))) & (~x4 | (x5 ? (~x2 & ~x3) : x3))))) : ((x2 | ((~x3 | x4 | x5) & (~x4 | ~x5 | x0 | x3))) & (~x0 | (x3 ? ((x4 | ~x5) & (~x2 | ~x4 | x5)) : (x4 | x5))) & (~x2 | x4 | (x3 & ~x5)));
  assign n3035 = (x5 | x6 | ~x7 | x0 | x1 | ~x4) & (x4 | ((x0 | ((x6 | ~x7 | ~x1 | ~x5) & (x1 | ~x6 | x7))) & (~x6 | x7 | ((x1 | ~x5) & (~x0 | ~x1 | x5)))));
  assign n3036 = n616 & ((n648 & n1172) | (x1 & ~n1465));
  assign n3037 = (x1 | ((~x4 | n630 | x0 | ~x2) & (~x0 | (x2 ? n856 : (~x4 | n630))))) & (x0 | ~x1 | (x2 ? (x4 | n630) : n856));
  assign z236 = ~n3046 | n3039 | ~n3041;
  assign n3039 = x1 & ((n2314 & n698) | (~x0 & ~n3040));
  assign n3040 = x2 ? (((x4 ? (x5 | ~x7) : (~x5 | x7)) | (x3 ^ x6)) & (~x3 | x6 | ~x7 | (~x4 ^ ~x5))) : ((x6 | x7 | x4 | x5) & (~x7 | ((~x3 | ~x4 | ~x5 | ~x6) & (x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))))));
  assign n3041 = ~n3044 & (~x2 | n3045) & (x1 | (~n3042 & ~n3043));
  assign n3042 = ~n721 & ((~x3 & x4 & x5 & x6 & ~x7) | (~x4 & ~x6 & (x3 ? (~x5 ^ x7) : (~x5 & x7))));
  assign n3043 = x6 & n1701 & ((n616 & n2527) | (x0 & n549));
  assign n3044 = ~n1862 & (x1 ? ((~x3 & x5 & x0 & ~x2) | (~x0 & ~x5 & (x2 ^ ~x3))) : ((~x3 & x5 & ~x0 & x2) | (x3 & (x0 ? (x2 ^ x5) : (~x2 & ~x5)))));
  assign n3045 = (x0 | ~x1 | x3 | ~x4 | ~x5 | x7) & (x1 | (((x3 ^ x5) | (x0 ? (~x4 | ~x7) : (x4 | x7))) & (x5 | ~x7 | x0 | ~x3) & (x4 | ~x5 | x7 | ~x0 | x3)));
  assign n3046 = n3049 & (n620 | n3047) & (x2 | n3048);
  assign n3047 = (x0 | ~x1 | ~x2 | x3 | x4 | x5) & (~x4 | ((x2 | ((x3 | ~x5 | x0 | ~x1) & (~x0 | x5 | (~x1 ^ x3)))) & (x0 | x1 | ~x2 | x3 | x5)));
  assign n3048 = x0 ? ((x5 | x7 | x3 | x4) & (x1 | ((x4 | x5 | x7) & (x3 | ((x5 | x7) & (x4 | ~x5 | ~x7)))))) : ((x1 | x3 | (x4 ? (x5 | ~x7) : (~x5 | x7))) & (~x3 | ((~x5 | ~x7 | x1 | ~x4) & (~x1 | (x4 ? (x5 | x7) : (~x5 | ~x7))))));
  assign n3049 = (n1361 | n3051) & (~n535 | ~n1176) & (~x5 | n3050);
  assign n3050 = (x3 | x4 | x6 | x0 | x1 | ~x2) & (x2 | ((x0 | ~x1 | ~x3 | ~x4 | x6) & (~x0 | ((~x4 | ~x6 | ~x1 | x3) & (x4 | x6 | x1 | ~x3)))));
  assign n3051 = (~x0 | x2 | x3 | ~x5 | x6) & (x0 | ~x6 | (x2 ? (x3 | ~x5) : (~x3 | x5)));
  assign z237 = ~n3053 | (x1 ? (n3062 | (~x6 & ~n3061)) : ~n3057);
  assign n3053 = (~x1 | n3056) & (n620 | n3054) & (x1 | n3055);
  assign n3054 = (x1 | (x3 ? ((x4 | x5 | x0 | ~x2) & ((~x4 ^ x5) | (x0 ^ x2))) : ((~x4 | ~x5 | x0 | ~x2) & (x4 | x5 | (~x0 & x2))))) & (x3 | ~x4 | ~x5 | ~x0 | x2) & (~x1 | ((x2 | ~x3 | x4 | x5) & (x0 | ((x3 | x4 | ~x5) & (~x2 | ~x4 | (x3 ^ x5))))));
  assign n3055 = (x0 | ((x2 | ~x3 | x4 | x6 | x7) & (~x2 | ((x4 | ~x6 | ~x7) & (x3 | ~x4 | x6 | x7))))) & (x2 | x3 | ~x4 | ~x6 | ~x7) & (~x0 | ((x2 | ((x4 | ~x6 | ~x7) & (~x3 | ~x4 | x6))) & (~x6 | ~x7 | x3 | ~x4) & (~x2 | ~x3 | x4 | x6 | x7)));
  assign n3056 = (x0 | (x3 ? ((~x6 | ~x7 | x2 | ~x4) & (~x2 | (x4 ? (x6 | x7) : (~x6 | ~x7)))) : (x6 | (x4 ? x2 : x7)))) & (x2 | x3 | ((~x4 | x6 | x7) & (~x6 | ~x7 | ~x0 | x4)));
  assign n3057 = x0 ? (x2 ? n3059 : (x7 | n3058)) : (x2 ? n3060 : n3059);
  assign n3058 = (~x5 | x6 | x3 | ~x4) & (x4 | (x3 ? (~x5 ^ x6) : (~x5 | ~x6)));
  assign n3059 = x3 ? ((~x4 | ~x5 | ~x6) & (x4 | x5 | x6 | ~x7)) : (x4 ? (x7 | (~x5 ^ x6)) : (~x5 | ~x6));
  assign n3060 = (~x5 | x6 | x7 | ~x3 | ~x4) & ((~x3 ^ ~x6) | (x4 ? (x5 | ~x7) : (~x5 | x7)));
  assign n3061 = ((x0 ? (x2 | x3) : (~x2 | ~x3)) | (x4 ? (x5 | ~x7) : (~x5 | x7))) & (x0 | ((x5 | ~x7 | x3 | x4) & (x2 | ~x3 | ~x4 | ~x5 | x7)));
  assign n3062 = n1205 & ((x2 & ~x3 & x4 & x5) | (~x2 & ((x3 & (x4 ? (~x5 & ~x7) : x5)) | (~x4 & x5 & x7))));
  assign z238 = n3064 | ~n3071 | (~n620 & ~n3070) | (x1 & ~n3069);
  assign n3064 = ~x6 & ((n1887 & ~n3065) | n3067 | (~n1002 & ~n3066));
  assign n3065 = (~x5 | x7 | x3 | ~x4) & (x5 | ~x7 | ~x3 | x4);
  assign n3066 = (x0 | x2 | (x1 ^ x3)) & (~x2 | x3 | ~x0 | x1);
  assign n3067 = ~n3068 & ((n2327 & n691) | (~x2 & n746));
  assign n3068 = x0 ? (x1 | ~x3) : (~x1 | x3);
  assign n3069 = (x0 | x3 | x4 | x5 | ~x7) & (x2 | ((~x0 | ~x3 | x4 | x5 | x7) & (x0 | ((~x5 | x7 | ~x3 | ~x4) & (x3 | x5 | ~x7)))));
  assign n3070 = ((x4 ^ x5) | ((~x0 | ~x1 | x2 | x3) & (x0 | ~x2 | (x1 ^ x3)))) & (x4 | ~x5 | ((~x0 | x1 | ~x2 | ~x3) & (x0 | (x1 ? (~x2 | x3) : (x2 | ~x3)))));
  assign n3071 = ~n3073 & n3074 & (~x6 | (~n3072 & (~n924 | ~n683)));
  assign n3072 = ~x1 & ((~x4 & ~x5 & ~x7 & n2317) | (~n1606 & (x4 ? (x5 ^ ~x7) : (~x5 & x7))));
  assign n3073 = ~n824 & ((~x0 & x1 & (x2 ? (~x3 & x4) : (x3 & ~x4))) | (~x1 & (x0 ? ((~x3 & ~x4) | (x2 & x3 & x4)) : (x3 & (x2 ^ x4)))));
  assign n3074 = (x1 | n3075) & (n1002 | (x0 ? (x2 | (~x1 ^ x3)) : (~x2 | (x1 ^ x3))));
  assign n3075 = ((~x0 ^ ~x2) | ((x3 | ~x4 | ~x5 | x7) & (x5 | ~x7 | ~x3 | x4))) & (x0 | ~x5 | ((x2 | x3 | x4 | ~x7) & (~x4 | x7 | ~x2 | ~x3)));
  assign z239 = ~n3079 | (~x2 & (x0 ? ~n3077 : ~n3078));
  assign n3077 = (x7 | ((~x1 | x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (x4 | x5 | x6 | (x1 & ~x3)))) & (x1 | ~x7 | (x4 ? ((x5 | x6) & (~x3 | ~x5 | ~x6)) : (x5 | ~x6)));
  assign n3078 = (x5 | ((~x4 | ((x6 | x7 | x1 | ~x3) & (~x7 | (x1 ? (x3 ^ x6) : (x3 | ~x6))))) & (x1 | x4 | (x3 ? (~x6 | x7) : (x6 | ~x7))))) & (~x1 | ~x5 | ((x4 | x6 | ~x7) & (x3 | ~x6 | (~x4 ^ ~x7))));
  assign n3079 = ~n3080 & ~n3085 & ~n3086 & (x0 ? n3084 : n3083);
  assign n3080 = x2 & ((~x1 & ~n3081) | (~x7 & n664 & ~n3082));
  assign n3081 = x0 ? (x5 | ((~x3 | x4 | (~x6 ^ x7)) & (~x4 | (x3 ? (x6 | x7) : (~x6 | ~x7))))) : ((x7 | ((~x3 | x4 | x5 | x6) & (x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))))) & (~x3 | ~x7 | (x4 ? (~x5 ^ ~x6) : (x5 | ~x6))));
  assign n3082 = (~x5 | x6 | ~x3 | x4) & (x3 | (x4 ? (~x5 ^ ~x6) : (x5 | ~x6)));
  assign n3083 = x2 ? (x4 ? ((x5 | ~x6 | x1 | ~x3) & (~x5 | x6 | ~x1 | x3)) : ((~x5 | x6 | x1 | ~x3) & (~x6 | (x1 ? (~x3 ^ x5) : (x3 | x5))))) : ((x3 | ((~x5 | ~x6 | x1 | x4) & (~x1 | x5 | (x4 ^ x6)))) & (~x4 | ~x5 | x6 | (x1 & ~x3)));
  assign n3084 = (~x1 | x2 | x3 | x4 | x5 | ~x6) & (x1 | ((~x5 | (x2 ? ((~x4 | x6) & (~x3 | x4 | ~x6)) : (x4 | x6))) & (x2 | ~x4 | ~x6 | (x3 & x5))));
  assign n3085 = ~n846 & ((~x3 & ((~x0 & ~x1 & x2 & x4) | (x0 & (x1 ? (~x2 & x4) : (x2 & ~x4))))) | (~x0 & x3 & ((~x2 & ~x4) | (x1 & x2 & x4))));
  assign n3086 = ~n3087 & ((n690 & n543) | (n814 & n544));
  assign n3087 = (~x0 | x1 | ~x2 | ~x5) & (x0 | (x1 ? (~x2 | x5) : (x2 | ~x5)));
  assign z240 = ~n3091 | (~x6 & (x1 ? ~n3090 : ~n3089));
  assign n3089 = (~x3 | ~x4 | ~x7) & (~x0 | ((~x2 | x3 | x4 | x5 | x7) & (x2 | ~x4 | ((x5 | ~x7) & (x3 | ~x5 | x7)))));
  assign n3090 = (x4 | x5 | ((x0 | ~x3 | x7) & (x2 | ((x3 | x7) & (~x0 | ~x3 | ~x7))))) & (x0 | x3 | ~x7 | (~x4 & (x2 | ~x5)));
  assign n3091 = ~n3094 & ((~x6 & (x7 | n3095)) | (~n3093 & ((x7 & n3095) | (x6 & ~x7 & n3092))));
  assign n3092 = x3 ? (x4 | ((x1 | ~x5) & (x0 | ~x1 | x5))) : ((x1 | ((~x2 | x4 | x5) & (~x0 | x2 | ~x5))) & (~x1 | x2 | x4 | x5) & (x0 | ((x2 | x4 | x5) & (~x1 | (x2 ? (x4 | ~x5) : x5)))));
  assign n3093 = n733 & ((~x0 & x1 & ~x3 & (x2 ^ x5)) | (~x1 & ~x5 & (x2 ? x3 : x0)));
  assign n3094 = ~n2176 & ((x0 & ~x2 & (x1 ? (~x3 & x5) : ~x5)) | (~x0 & (x1 ? ((x2 & ~x3 & ~x5) | (x3 & x5)) : (~x3 & x5))) | (~x1 & ((x3 & ~x5) | (x2 & ~x3 & x5))));
  assign n3095 = (x2 | ((~x0 | ((~x1 | x3 | ~x4 | x5) & (x1 | x4 | ~x5))) & (~x3 | x4 | x0 | x1))) & (x3 | ((~x4 | x5 | x1 | ~x2) & (x0 | (x1 ? (~x5 | (~x2 & ~x4)) : (~x4 | x5))))) & (~x3 | ((x1 | ~x5) & (~x4 | x5 | x0 | ~x1)));
  assign z241 = ~n3102 | (~x5 & (n3097 | ~n3099));
  assign n3097 = n598 & (x2 ? (~x3 & n3098) : ((x3 & n3098) | (x4 & n543)));
  assign n3098 = ~x7 & ~x4 & x6;
  assign n3099 = ~n3101 & (n1041 | n3100) & (~n650 | ~n544 | ~n694);
  assign n3100 = x0 ? (x1 & (x2 | x3)) : (~x1 & (~x2 | ~x3));
  assign n3101 = ~x0 & ~x1 & ~x3 & (x2 ? (x4 & ~x6) : (~x4 & x6));
  assign n3102 = ((~x6 ^ ~x7) & (~n1449 | (n1799 & ~n720))) | (n3103 & (x6 ^ ~x7));
  assign n3103 = (x2 | ((x3 | ~x4 | ~x5) & (x0 | x1 | ~x3 | x4 | x5))) & (x1 | ~x4 | ~x5) & (x0 | ((~x4 | ~x5) & (x1 | ~x2 | x3 | x4 | x5)));
  assign z242 = ~n3106 | (~x7 & n598 & ~n3105);
  assign n3105 = (x4 | x5 | x6 | ~x2 | x3) & (x2 | (x5 ? ~x6 : ((~x3 & ~x4) | x6)));
  assign n3106 = ~n3107 & (~n698 | ~n754) & (x2 | ~n1156 | ~n598);
  assign n3107 = (~x0 | ~x1 | (~x2 & ~x3)) & (x0 | x1 | x2) & (~x5 | ~x7) & (x5 | x7);
  assign z243 = n3111 | n3112 | (n677 & n3109) | (n1835 & ~n3110);
  assign n3109 = ~x7 & x3 & ~x6;
  assign n3110 = (~x3 | x5 | ~x6 | ~x0 | ~x1 | x2) & (x0 | x1 | x3 | (x2 ? (x5 ^ x6) : (~x5 | x6)));
  assign n3111 = x6 & (x1 ? (~x0 | (~x2 & ~x3)) : (x0 | x7 | (x2 & x3)));
  assign n3112 = ~x3 & x4 & ~x7 & n598 & (x2 ^ ~x6);
  assign z244 = ~n3116 | (~x4 & ((n732 & ~n3114) | (~x2 & ~n3115)));
  assign n3114 = (x5 | ~x7 | ~x1 | x2) & (x1 | (x2 ? (~x5 ^ ~x7) : (~x5 | x7)));
  assign n3115 = (~x0 | ~x1 | ~x3 | x5 | x6 | ~x7) & (x0 | x3 | ((x6 | ~x7 | ~x1 | ~x5) & (~x6 | x7 | x1 | x5)));
  assign n3116 = (~x0 & ((~x2 & ~x3 & ~x4) | (~x1 & ((~x3 & ~x4) | (~x2 & x7))))) | (x2 & (~x7 | (x0 & x1))) | (x1 & ~x7) | (x0 & (~x7 | (x1 & x3)));
  assign z245 = ~n3123 | ~n3122 | n3118 | n3121;
  assign n3118 = ~x2 & ((n735 & ~n3119) | (~x4 & n732 & n3120));
  assign n3119 = (x1 | x3 | ~x4 | ~x5 | x6) & (~x1 | ~x3 | x4 | x5 | ~x6);
  assign n3120 = x7 & (x1 ? (x5 & x6) : (~x5 & ~x6));
  assign n3121 = ~x0 & ((x3 & x4 & x5 & x1 & x2) | (~x1 & ~x3 & ~x4 & (x2 ^ x5)));
  assign n3122 = x1 | x2 | ((x0 | (~x3 & ~x4)) & (x3 | (x4 ? x5 : ~x0)));
  assign n3123 = (x0 | x1 | x3 | ~x6 | ~n2014) & (~x0 | (x1 ? (x3 ? (x6 | ~n2014) : x2) : ~x2));
  assign z246 = n3126 | ~n3127 | (x6 & ~n3125);
  assign n3125 = (x0 | ~x1 | ~x2 | x3 | x4 | x5) & (x1 | ~x4 | ((~x3 | ~x5 | x0 | ~x2) & (~x0 | (x2 ? (~x3 | x5) : (x3 | ~x5)))));
  assign n3126 = x1 & ((~x3 & ((~x0 & x2 & x5) | (~x2 & (x0 | ~x4)))) | (~x0 & x2 & (x5 ? ~x4 : (x3 | x4))));
  assign n3127 = ~n3128 & ~n3129 & (x2 | (~n766 & (~n678 | ~n958)));
  assign n3128 = n694 & n1112;
  assign n3129 = ~x1 & ((~x0 & ((~x2 & x4 & x5) | (~x4 & ~x5 & x2 & ~x3))) | (x3 & (~x2 | (x0 & x4 & x5))));
  assign z247 = ~n3133 | (x7 & (x0 ? ~n3132 : ~n3131));
  assign n3131 = (~x4 | ~x5 | ~x6 | ~x1 | ~x2 | x3) & (x4 | ((x1 | ~x2 | ~x3 | x5 | x6) & (x2 | ((~x1 | ~x5 | (~x3 ^ x6)) & (x5 | x6 | x1 | x3)))));
  assign n3132 = (~x1 | x2 | x3 | x4 | ~x5 | ~x6) & (x1 | ((~x2 | x3 | ~x4 | ~x5 | x6) & (x2 | x5 | (x3 ? (x4 | ~x6) : (~x4 | x6)))));
  assign n3133 = (~n3134 | n3137) & (x1 | n3135) & (~x1 | n3136);
  assign n3134 = ~x2 & ~x7;
  assign n3135 = (~x4 & ((x3 & ((~x2 & ~x5) | (~x0 & (~x2 | (~x5 & ~x6))))) | (~x2 & ~x5 & ~x6) | (~x3 & (x0 | (x2 & x5))))) | (x0 & ~x3 & ~x6) | (x4 & ((x2 & ((x0 & (x5 ^ x6)) | (~x3 & ~x6) | (x3 & x5 & x6))) | (~x3 & ((~x2 & x5) | (~x0 & x6)))));
  assign n3136 = (x2 | (x0 ? ((x3 | ~x4) & (x5 | x6 | ~x3 | x4)) : (~x3 | ~x4))) & (x0 | ((~x3 | ~x4 | x5) & (x4 | ((~x3 | ~x5 | ~x6) & (~x2 | (~x3 & (x5 | x6)))))));
  assign n3137 = (x0 | x1 | x3 | ~x4 | x5 | ~x6) & (~x0 | ((x1 | x3 | ~x4 | ~x5 | x6) & (~x1 | ~x3 | x4 | x5 | ~x6)));
  assign z248 = n3139 | ~n3142 | n3148 | (~x0 & ~n3147);
  assign n3139 = x1 & ((n665 & n1835 & ~n3141) | (~x3 & ~n3140));
  assign n3140 = (x0 | ~x2 | ~x4 | x5 | x6 | ~x7) & (~x5 | ((x0 | ~x2 | ~x4 | ~x6 | x7) & (x2 | (x0 ? (x4 ? (x6 | ~x7) : (~x6 | x7)) : (~x7 | (x4 ^ x6))))));
  assign n3141 = x0 ? (x5 | ~x6) : (~x5 | x6);
  assign n3142 = ~n3144 & ~n3146 & (n783 | n3145) & (~x0 | n3143);
  assign n3143 = (x1 | ~x2 | ~x3 | ~x4 | x5 | x6) & (x4 | ((~x1 | x2 | ~x3 | x5 | x6) & (x1 | x3 | ~x6 | (x2 & ~x5))));
  assign n3144 = ~x1 & ((x5 & (x0 ? (x3 & (x2 ^ x4)) : (~x3 & (~x2 ^ x4)))) | (x2 & ~x5 & (x0 ? (~x3 & x4) : (x3 ^ ~x4))));
  assign n3145 = (~x2 | x3 | x5 | x0 | ~x1) & (x2 | ((x0 | x1 | ~x3 | ~x5) & (~x0 | ((x3 | ~x5) & (x1 | ~x3 | x5)))));
  assign n3146 = x1 & ((~x3 & ~x4 & ~x5 & x0 & ~x2) | (~x0 & x3 & (x2 ? (x4 & ~x5) : (~x4 ^ x5))));
  assign n3147 = (~x5 | ((x3 | x4 | ~x6 | ~x1 | x2) & (~x2 | ((~x4 | x6 | x1 | ~x3) & (~x1 | (x3 ? (x4 | ~x6) : (~x4 | x6))))))) & (x1 | x2 | ((~x3 | x4 | ~x6) & (x3 | ~x4 | x5 | x6)));
  assign n3148 = ~x1 & ((n1120 & ~n1568 & ~n3149) | (~x6 & ~n3150));
  assign n3149 = x0 ? (~x3 | x4) : (x3 | ~x4);
  assign n3150 = (~x0 | x2 | ~x4 | x5 | (~x3 ^ ~x7)) & ((x2 ^ ~x7) | ((~x4 | ~x5 | ~x0 | x3) & (x4 | x5 | x0 | ~x3)));
  assign z249 = n3155 | ~n3158 | (x2 & ~n3153) | (~x0 & ~n3152);
  assign n3152 = x3 ? ((~x6 | (x1 ? (x5 | (x2 & x4)) : (x4 | ~x5))) & (x1 | ~x5 | x6 | (x2 & ~x4))) : (((x5 ^ x6) | (x1 ? (~x2 | x4) : ~x4)) & (~x5 | x6 | ~x1 | ~x4) & (x4 | x5 | ~x6 | (x1 & x2)));
  assign n3153 = (x1 | n3154) & (x0 | ~x1 | (~n2356 & (n692 | ~n2476)));
  assign n3154 = x4 ? ((x3 ^ x7) | (x0 ? (~x5 | x6) : (x5 | ~x6))) : ((~x5 | x6 | ~x7 | x0 | ~x3) & (x5 | (x3 ^ ~x7) | (x0 ^ x6)));
  assign n3155 = ~x2 & (x0 ? ~n3156 : ~n3157);
  assign n3156 = (x3 | ((x6 | x7 | ~x4 | ~x5) & (~x1 | x4 | ~x6 | (~x5 ^ x7)))) & (~x3 | x4 | x5 | ~x6 | x7) & (x1 | ~x4 | x6 | ((x5 | x7) & (~x3 | ~x5 | ~x7)));
  assign n3157 = x5 ? ((x6 | x7 | ~x1 | x4) & (~x6 | ((x3 | x4 | ~x7) & (~x1 | ~x4 | (x3 ^ x7))))) : (x3 ? ((~x1 | ~x4 | x6 | ~x7) & (x1 | (x4 ? (~x6 | ~x7) : (x6 | x7)))) : ((~x6 | x7 | x1 | ~x4) & (x4 | x6 | ~x7)));
  assign n3158 = (~x0 | n3159) & (n850 | ((x0 | ~x1 | ~x2 | ~x3) & (~x0 | x3 | (x1 ^ ~x2))));
  assign n3159 = (x2 | ~x3 | x4 | x5 | x6) & (x1 | ((x2 | x4 | (x5 ^ x6)) & (~x3 | ((~x5 | ~x6) & (~x2 | x5 | x6)))));
  assign z250 = (~x2 & ~n3161) | (~x0 & ~n3164) | ~n3166 | (x0 & ~n3165);
  assign n3161 = (x3 | n3163) & (n671 | n2348) & (n1429 | n3162);
  assign n3162 = (~x3 | x4 | x0 | x1) & (x3 | ~x4 | ~x0 | ~x1);
  assign n3163 = (~x0 | ~x1 | ~x4 | x5 | x6 | ~x7) & (~x5 | ((x0 | x1 | ~x4 | ~x6 | ~x7) & (x7 | ((x0 | ~x1 | x4 | ~x6) & (~x0 | x6 | (~x1 ^ ~x4))))));
  assign n3164 = (x2 | ((~x5 | x6 | x1 | ~x4) & (x5 | ((~x6 | ~x7 | x1 | x4) & (~x1 | (x4 ? ~x6 : (x6 | x7))))))) & (x1 | ~x5 | (x4 ? (x6 | ~x7) : (~x6 | (~x2 & x7))));
  assign n3165 = (~x6 | ((~x1 | x2 | x4 | x5 | x7) & (x1 | ((~x5 | ~x7 | x2 | ~x4) & (~x2 | x4 | x5 | x7))))) & (x1 | ~x2 | x6 | ~x7 | (~x4 ^ x5));
  assign n3166 = ~n3169 & n3170 & (x6 ? (x7 ? n3167 : n3168) : (x7 ? n3168 : n3167));
  assign n3167 = (x0 | ~x1 | ((x4 | ~x5) & (~x2 | ~x4 | x5))) & (x1 | ((x4 | x5 | x0 | ~x2) & (~x0 | ~x4 | (~x2 & x5))));
  assign n3168 = (x2 | ((~x0 | x4 | (x1 ? (x3 | ~x5) : (~x3 | x5))) & (~x4 | ~x5 | x0 | ~x1))) & (x0 | ~x4 | (x1 ? (x3 | ~x5) : x5));
  assign n3169 = ~n2176 & (x2 ? (n664 & n985) : (n738 & n916));
  assign n3170 = (n2176 | n3171) & (n3172 | (~n644 & (~n2205 | ~n538)));
  assign n3171 = (~x2 | x5 | x0 | ~x1) & (x2 | ~x5 | ~x0 | x1);
  assign n3172 = (~x0 | x3 | ~x4 | ~x6) & (x0 | ~x3 | x4 | x6);
  assign z251 = ~n3179 | n3174 | n3176;
  assign n3174 = x7 & ((n750 & n1112) | (~x2 & ~n3175));
  assign n3175 = (~x1 | ((~x0 | ~x3 | x4 | x5 | x6) & (x0 | x3 | (x4 ? x5 : (~x5 | x6))))) & (~x0 | x1 | ~x5 | (x3 ? (x4 | x6) : (~x4 | ~x6)));
  assign n3176 = ~x7 & ((x6 & ~n3177) | (~x0 & ~x6 & ~n3178));
  assign n3177 = (~x0 | x1 | x2 | x3 | x4 | ~x5) & ((x4 ^ x5) | ((~x0 | x1 | ~x2 | ~x3) & (x0 | ~x1 | x2 | x3)));
  assign n3178 = (x1 | ~x2 | x3 | ~x4 | ~x5) & (x2 | ((~x4 | x5 | x1 | x3) & (~x1 | ~x3 | (~x4 ^ x5))));
  assign n3179 = ~n3180 & ~n3182 & ~n3183 & n3184 & (x2 | n3181);
  assign n3180 = ~n824 & ((~x6 & ((x0 & ~x1 & ~x2 & ~x3) | (~x0 & x1 & x2 & x3))) | (~x1 & ((~x0 & x3 & x6) | ((~x0 | x6) & (x2 ^ x3)))));
  assign n3181 = (x0 | ~x1 | x6 | (x3 ? (x5 | ~x7) : (~x5 | x7))) & (x1 | ((~x5 | x6 | ~x7 | x0 | x3) & (~x0 | ((~x6 | ~x7 | x3 | x5) & (x6 | x7 | ~x3 | ~x5)))));
  assign n3182 = ~x3 & ((~x0 & ~x5 & (x1 ? (x2 & ~x6) : (~x2 & x6))) | (x0 & x1 & ~x2 & x5 & x6));
  assign n3183 = ~n800 & (x0 ? (~x6 & (x1 ? (~x2 & ~x3) : x2)) : (x1 & x6 & (x2 | x3)));
  assign n3184 = ~x3 | ~x5 | ~n538 | (x0 ? (~x6 | ~x7) : x6);
  assign z252 = ~n3189 | (~n1115 & ~n3193) | (~x1 & (~n3186 | ~n3194));
  assign n3186 = (~x2 | ~n3187) & (~x0 | ~n3188 | (x2 ^ ~x4));
  assign n3187 = ~x7 & ((~x0 & ~x3 & x4 & ~x5 & x6) | (~x6 & ((~x0 & x3 & x4 & x5) | (x0 & ~x4 & (~x3 ^ x5)))));
  assign n3188 = ~x6 & x7 & (x3 ^ ~x5);
  assign n3189 = ~n3190 & ~n3191 & (~n588 | ~n1231) & (n620 | n3192);
  assign n3190 = ~n2354 & ((x0 & ~x1 & ~x2 & n540) | (~x0 & (x1 ? (x2 ? n540 : n537) : (x2 & n537))));
  assign n3191 = n664 & (x2 ? (x7 & (x3 ? (x4 & ~x6) : x6)) : (~x7 & (x3 ? (x4 ^ x6) : (x4 ^ ~x6))));
  assign n3192 = (x0 | x1 | x2 | x3) & (~x0 | ((x1 | ~x2 | ~x3 | ~x4) & (~x1 | x2 | (x3 & (x4 | x5)))));
  assign n3193 = x0 ? (x1 | (x2 ? (x4 | x6) : ((~x4 | ~x6 | ~x7) & (x6 | x7)))) : ((~x1 | (x2 ? (x6 | x7) : (~x6 | ~x7))) & (~x2 | ((x1 | ~x6 | ~x7) & (~x4 | x6 | x7))));
  assign n3194 = x3 ? ((~x6 | ~x7 | x2 | x4) & (x0 | ((x2 | ~x6) & (x6 | x7 | ~x2 | x4)))) : ((x4 | ~x6 | x7 | x0 | ~x2) & (~x0 | x6 | (x2 ? ~x4 : (x4 | ~x7))));
  assign z253 = ~n3196 | ~n3199 | n3201 | (~x0 & ~n3202);
  assign n3196 = ~n3198 & n3197 & (~x3 | x4 | ~n2488 | ~n2758);
  assign n3197 = (x0 | x1 | ~x3 | (~x2 ^ x7)) & (x3 | ((x0 | ~x1 | ~x2 | x7) & (~x0 | (x1 ? (x2 | x7) : (~x2 | ~x7)))));
  assign n3198 = ~x2 & ((x5 & ~n1323 & ~n2656) | (n686 & n958));
  assign n3199 = ~n3200 & (~n664 | ((x2 | x3 | x4 | x7) & (~x4 | (x2 ? (~x3 | ~x7) : (~x3 ^ x7)))));
  assign n3200 = n651 & ((~x4 & ~x5 & ~x7 & x1 & x3) | (~x1 & x4 & (x3 ? (x5 ^ ~x7) : (~x5 & x7))));
  assign n3201 = ~x1 & ((~x3 & ((~x4 & x7 & x0 & ~x2) | (~x0 & (x2 ? (~x4 & x7) : (x4 & ~x7))))) | (x0 & x3 & (x2 ? (x4 ^ x7) : (~x4 & ~x7))));
  assign n3202 = (x1 | ~x2 | x3 | ~x4 | (~x5 ^ x7)) & (x4 | ((x1 | x2 | x3 | ~x5 | x7) & (~x1 | ~x3 | ~x7 | (x2 ^ x5))));
  assign z255 = ~n3208 | (x1 ? ~n3204 : (x2 ? ~n3206 : ~n3207));
  assign n3204 = x0 ? (~n563 | ~n568) : n3205;
  assign n3205 = (x2 | ~x3 | x4 | ~x5 | ~x6 | ~x7) & (~x4 | ((x2 | ~x3 | ~x5 | x6 | x7) & (x5 | ((x6 | ~x7 | x2 | x3) & (~x2 | x7 | (~x3 ^ x6))))));
  assign n3206 = (x6 | ((~x0 | ~x3 | x4 | x5 | x7) & (x0 | ((x3 | x4 | ~x5 | x7) & (x5 | ~x7 | ~x3 | ~x4))))) & (~x0 | ~x4 | ~x6 | (x3 ? (~x5 | x7) : (x5 | ~x7)));
  assign n3207 = (~x4 | ((x0 | x3 | x5 | x6 | x7) & (~x0 | ~x5 | ~x7 | (~x3 ^ x6)))) & (x0 | x4 | ~x6 | (x3 ? (~x5 | x7) : (x5 | ~x7)));
  assign n3208 = n987 & (x0 ? (~x5 | n3210) : n3209);
  assign n3209 = (x5 | ((~x1 | x2 | x3 | ~x4 | ~x6) & (~x2 | (x1 ? (x3 ? (x4 | ~x6) : (~x4 | x6)) : (~x3 | (x4 ^ x6)))))) & (x1 | x2 | ~x3 | ~x5 | (x4 ^ x6));
  assign n3210 = (~x1 | x2 | x3 | x4 | ~x6) & (x1 | ((~x4 | x6 | ~x2 | ~x3) & (x2 | ((x4 | x6) & (~x3 | ~x4 | ~x6)))));
  assign z256 = ~n3213 | ~n3216 | (x2 ? ~n994 : ~n3212);
  assign n3212 = (x3 | ((~x0 | (x1 ? (~x5 | ~x6) : (x5 | x6))) & (x0 | ((~x4 | x5 | ~x6) & (~x5 | x6 | x1 | x4))) & (x5 | x6 | ~x1 | x4))) & (~x0 | x1 | x4 | ~x5 | ~x6) & (~x3 | ((~x4 | ~x5 | ~x6 | (x0 & x1)) & (x5 | ((x1 | x4 | x6) & (x0 | (x6 & (x1 | x4)))))));
  assign n3213 = x7 ? ((~x5 | n3214) & (x2 | ~x4 | n3215)) : ((x5 | n3214) & (~x2 | x4 | n3215));
  assign n3214 = (x3 | x4 | x6 | x0 | x1 | ~x2) & (x2 | ((~x3 | x4 | ~x6 | x0 | ~x1) & (~x0 | ~x4 | x6 | (~x1 ^ x3))));
  assign n3215 = (~x0 | x1 | x3 | ~x5 | ~x6) & (x0 | ~x1 | x6 | (~x3 ^ ~x5));
  assign n3216 = x0 ? (x1 | n3219) : (~n3218 & (~x4 | n3217));
  assign n3217 = (x1 | ((x2 | x3 | x5 | x6 | ~x7) & (~x5 | x7 | (x2 ? (~x3 ^ x6) : (x3 | x6))))) & (~x2 | x5 | ~x7 | ((~x3 | x6) & (~x1 | x3 | ~x6)));
  assign n3218 = x6 & n1148 & ((x1 & ~x3 & ~x5 & ~x7) | (~x1 & x7 & (x3 ^ ~x5)));
  assign n3219 = (x5 | ~x6 | x7 | x2 | x4) & (~x2 | ((~x3 | x4 | ~x5 | x6 | x7) & (~x7 | ((x5 | ~x6 | x3 | ~x4) & (~x3 | (x4 ? (~x5 | ~x6) : (x5 | x6)))))));
  assign z257 = ~n3223 | (~x5 & (x7 ? ~n3221 : ~n3222));
  assign n3221 = (~x6 | (x0 ? (x1 | (x2 ? (x3 | ~x4) : x4)) : (x3 | ((x2 | x4) & (~x1 | ~x2 | ~x4))))) & (x0 | ~x1 | x6 | (x2 ? (~x3 ^ ~x4) : (x3 | ~x4)));
  assign n3222 = (x1 | ((~x3 | ((x4 | x6 | x0 | ~x2) & ((~x0 ^ x4) | (~x2 ^ ~x6)))) & (~x2 | x3 | (x0 ? (~x4 | x6) : (x4 | ~x6))))) & (x2 | x3 | ((~x4 | ~x6) & (x4 | x6 | ~x0 | ~x1)));
  assign n3223 = ~n3224 & n3229 & (x6 | n3227) & (x2 | n3228);
  assign n3224 = x5 & ((n664 & ~n3226) | (~x1 & ~n3225));
  assign n3225 = ((x6 ^ x7) | ((~x3 | x4 | x0 | x2) & (~x2 | (x0 ? (~x3 ^ ~x4) : (x3 | ~x4))))) & (~x6 | ((x0 | ~x2 | ~x3 | x4 | x7) & (~x0 | x2 | x3 | ~x4 | ~x7)));
  assign n3226 = (x2 | x3 | x4 | x6 | x7) & (~x3 | (~x6 ^ x7) | (~x2 ^ x4));
  assign n3227 = (~x3 | ~x4 | ~x5 | x0 | ~x1 | ~x2) & (x3 | ((~x2 | ((x0 | (x1 ? (x4 | ~x5) : (~x4 | x5))) & (x4 | x5 | ~x0 | x1))) & (x0 | ~x1 | x2 | (x4 ^ x5))));
  assign n3228 = x3 ? (x0 ? (x1 | ~x4 | (~x6 ^ x7)) : (~x1 | x4 | (x6 ^ x7))) : (x6 | ((~x4 | ~x7 | x0 | x1) & (~x0 | (x1 ? (~x4 | ~x7) : (x4 | x7)))));
  assign n3229 = (~x6 | n3230) & (n1007 | n1009) & (~x2 | x6 | n3231);
  assign n3230 = (x2 | (x0 ? (x4 | (x1 ? (x3 | x5) : ~x5)) : (~x3 | ~x4 | (x1 & x5)))) & (x0 | ~x2 | ((~x3 | x4 | x5) & (~x4 | ~x5 | ~x1 | x3)));
  assign n3231 = (x0 | ~x1 | x3 | ~x4 | x7) & (x1 | ~x7 | (x0 ? (~x3 | x4) : (~x3 ^ ~x4)));
  assign z258 = ~n3236 | (x3 ? (n3235 | (~x1 & ~n2220)) : ~n3233);
  assign n3233 = (x2 | n3234) & (~n738 | n1002 | ~x2 | x6);
  assign n3234 = (x1 | (x0 ? (~x6 | (x4 ? (x5 | ~x7) : (~x5 | x7))) : (x5 | x6 | (~x4 ^ x7)))) & (x0 | ~x1 | x5 | ~x7 | (~x4 ^ x6));
  assign n3235 = ~n824 & (x0 ? (~x1 & n2403) : (~x4 & ~n1117));
  assign n3236 = ~n3238 & ~n3239 & ~n3240 & n3241 & (n620 | n3237);
  assign n3237 = x3 ? ((~x0 | x1 | ~x2 | x4 | ~x5) & (x0 | ~x4 | x5 | (~x1 ^ ~x2))) : ((~x1 | (x4 ^ x5) | (~x0 ^ x2)) & (x0 | x1 | ~x5 | (~x2 ^ x4)));
  assign n3238 = ~n824 & (((x0 ? (~x1 & x2) : (x1 & ~x2)) & (x3 ^ ~x4)) | (x0 & ~x1 & ~x2 & ~x3 & x4) | (~x0 & ((x3 & ~x4 & x1 & x2) | (~x1 & (x2 ? (~x3 & x4) : (x3 & ~x4))))));
  assign n3239 = ~x2 & ((n1153 & n1880) | (~x5 & n541 & ~n1150));
  assign n3240 = n616 & ((n1153 & n758) | (~x4 & n1156 & n605));
  assign n3241 = (n1002 | ((x0 | x1 | x2 | x3) & ((~x1 ^ x3) | (~x0 ^ x2)))) & (n3065 | (x0 ? (x1 | ~x2) : (~x1 | x2)));
  assign z259 = ~n3246 | (x3 & ~n3243);
  assign n3243 = (n607 | n3245) & (~x0 | ~n539 | ~n559) & (x0 | n3244);
  assign n3244 = (~x5 | ((~x4 | ((x6 | ~x7 | x1 | ~x2) & (x7 | (x1 ? (~x2 ^ x6) : (x2 | x6))))) & (x1 | x4 | ~x6 | (x2 ^ x7)))) & (x1 | x4 | x5 | x6 | (x2 ^ x7));
  assign n3245 = (~x0 | x1 | x4 | x5 | ~x6) & ((x0 ? (x1 | ~x4) : (~x1 | x4)) | (~x5 ^ ~x6));
  assign n3246 = ~n3247 & (x3 | n3250) & (x5 ? n3248 : n3249);
  assign n3247 = ~n846 & ((x2 & ((~x0 & x4 & (x1 ^ x3)) | (~x1 & ~x4 & (x0 | ~x3)))) | (x0 & ~x3 & (x1 ? (~x2 & x4) : ~x4)));
  assign n3248 = (x1 | x2 | x3 | ~x4 | ~x6) & (x6 | ((x1 | ((x2 | ~x3 | x4) & (~x4 | ((~x2 | x3) & (~x0 | (~x2 & x3)))))) & (x0 | ((x2 | x3 | x4) & (~x1 | (x2 ? (~x3 | x4) : ~x4))))));
  assign n3249 = (x0 | ~x1 | x2 | ~x3 | ~x4 | x6) & (~x6 | ((~x3 | ((x1 | x2 | ~x4) & (x0 | (x1 ? (x2 ^ x4) : (~x2 | x4))))) & (~x1 | x3 | x4 | (~x0 ^ x2))));
  assign n3250 = x0 ? (n850 | (~n1599 & (~x1 | ~n3134))) : n3251;
  assign n3251 = (x5 | ((~x6 | ((~x1 | (x2 ? (~x4 | x7) : ~x7)) & (x2 | x4 | ~x7) & (x1 | x7 | (x2 ^ ~x4)))) & (x1 | ~x4 | x6 | (x2 ^ ~x7)))) & (~x1 | x4 | ((x2 | ~x6 | ~x7) & (x6 | x7 | ~x2 | ~x5)));
  assign z260 = (~x2 & (~n3254 | (~x3 & ~n3253))) | ~n3257;
  assign n3253 = x6 ? ((x1 | x4 | ~x5 | x7) & (x0 | ((x1 | x5 | ~x7) & (x4 | ~x5 | x7)))) : ((x5 | ~x7 | x1 | ~x4) & (~x0 | ((~x1 | x4 | x5 | x7) & (x1 | ~x4 | ~x5))));
  assign n3254 = (x7 | n3255 | x3 | ~x6) & (~x3 | ((x1 | n3256) & (~x7 | n3255 | ~x1 | x6)));
  assign n3255 = x0 ? (x4 | x5) : (~x4 | ~x5);
  assign n3256 = x0 ? ((~x6 | x7 | x4 | ~x5) & (~x4 | x5 | x6 | ~x7)) : (x5 ? (x6 | ~x7) : (x7 | (~x4 ^ x6)));
  assign n3257 = ~n3259 & (n662 | n3258) & (~x2 | (~n3260 & n3261));
  assign n3258 = (x0 | ((~x1 | ((x3 | x5) & (x2 | ~x3 | ~x5))) & (x1 | ~x4 | ((x3 | ~x5) & (~x2 | ~x3 | x5))) & (x4 | ((~x3 | ~x5) & (~x2 | x3 | x5))))) & (x5 | ((~x1 | x2 | x3 | ~x4) & (~x0 | x1 | (x4 ? x3 : x2)))) & (~x0 | x1 | ~x3 | (x4 & ~x5));
  assign n3259 = ~n2176 & (x3 ? ((~x1 & ~x5) | (~x0 & (~x5 | (~x1 & x2)))) : (x5 & (x0 ^ (x1 & x2))));
  assign n3260 = n1416 & ((x1 & ~x3 & x4 & x5 & ~x6) | (~x1 & x6 & (x3 ? (~x4 & ~x5) : x5)));
  assign n3261 = ((~x3 ^ ~x5) | (x0 ? (x1 | ~n3098) : ~n3262)) & (x3 | ~n3098 | x0 | ~x1) & (~x0 | x1 | ~x3 | ~n3262);
  assign n3262 = x7 & x4 & ~x6;
  assign z261 = ~n3269 | (x2 ? ~n3266 : (x0 ? ~n3264 : ~n3265));
  assign n3264 = (x5 | ~x6 | x7 | ~x1 | ~x3 | x4) & (x1 | (x3 ? ((x4 | ~x5 | ~x6 | x7) & (~x4 | x6 | ~x7)) : (~x5 | ~x7 | (~x4 & x6))));
  assign n3265 = (x3 | ((x6 | ~x7 | x4 | x5) & (~x1 | ((x5 | x6 | ~x7) & (x4 | ~x5 | x7))))) & (~x1 | ~x5 | ((~x4 | ~x6 | x7) & (~x3 | x4 | x6 | ~x7)));
  assign n3266 = x0 ? (x1 | n3268) : n3267;
  assign n3267 = (~x1 | ~x3 | ~x4 | ~x5 | ~x6 | x7) & (x1 | ((~x3 | ~x5 | (x4 ? (x6 | ~x7) : (~x6 | x7))) & (x5 | (x4 ? (~x6 | x7) : (x6 | ~x7)))));
  assign n3268 = (~x4 | x5 | x6 | ~x7) & (x4 | ~x6 | x7 | (x3 & x5));
  assign n3269 = n3272 & (x6 ? (x7 ? n3271 : n3270) : (x7 ? n3270 : n3271));
  assign n3270 = (x4 | ((~x1 | ((x3 | ~x5 | ~x0 | x2) & (x0 | x5 | (~x2 & ~x3)))) & (~x0 | x1 | (x2 ? (~x3 | ~x5) : (x3 | x5))))) & (x0 | x1 | ~x4 | ~x5 | (x2 & x3));
  assign n3271 = x1 ? ((x0 | ~x4 | x5) & (x2 | ((x3 | ~x4 | ~x5) & (x0 | (~x4 & (x3 | x5)))))) : ((~x2 | ((x4 | x5) & (~x0 | ~x4 | ~x5))) & (x2 | x3 | ((x4 | ~x5) & (~x0 | ~x4 | x5))) & (x0 | x4 | ~x5) & (~x0 | ~x3 | (x4 ^ x5)));
  assign n3272 = (~x1 | n3273) & (x0 | x1 | ~n1184 | n3274);
  assign n3273 = (x4 | ~x5 | x6 | x0 | ~x2) & (x3 | ((~x0 | x2 | x5 | (~x4 ^ x6)) & (~x4 | ~x5 | ~x6 | x0 | ~x2)));
  assign n3274 = (~x4 | ~x6) & (~x3 | x4 | x6);
  assign z262 = ~n3278 | ~n3283 | (~x0 & (n3277 | (~x3 & ~n3276)));
  assign n3276 = (~x7 | (x1 ? (x2 | ((x5 | x6) & (x4 | ~x5 | ~x6))) : (~x2 | (~x5 ^ ~x6)))) & (x4 | ~x6 | x7 | (x1 ? (~x2 | x5) : (x2 | ~x5)));
  assign n3277 = x7 & n904 & ((n1365 & n2326) | (x2 & ~n846));
  assign n3278 = ~n3279 & ~n3280 & (x1 ? (x0 | n3282) : n3281);
  assign n3279 = x2 & ((x3 & ~x5 & x7 & x0 & ~x1) | (~x0 & ((x5 & ~x7 & ~x1 & ~x3) | (x1 & (x3 ? (~x5 & ~x7) : (x5 & x7))))));
  assign n3280 = ~x2 & (((~x1 ^ x7) & (x0 ? (~x3 & ~x5) : (x3 & x5))) | (~x5 & x7 & ~x0 & ~x1) | (~x3 & x5 & ~x7 & x0 & x1));
  assign n3281 = (x0 | x2 | x3 | ~x4 | ~x5 | x7) & (~x0 | x5 | ((~x4 | ~x7 | ~x2 | x3) & (x2 | ~x3 | x4 | x7)));
  assign n3282 = (x2 | x3 | ~x4 | ~x5 | ~x7) & (~x2 | ((~x3 | x4 | ~x5 | ~x7) & (x5 | x7 | x3 | ~x4)));
  assign n3283 = (n912 | n3284) & (~x0 | (~n3285 & (~n698 | ~n811)));
  assign n3284 = (x1 | ((~x3 | x7 | x0 | ~x2) & (~x0 | ~x7 | (x2 & (x3 | x4))))) & (x0 | ~x1 | ((x2 | x7) & (~x4 | ~x7 | ~x2 | ~x3)));
  assign n3285 = n873 & ((~x2 & x3 & n872) | (~n846 & (x2 | n814)));
  assign z263 = ~n3287 | n3296 | n3297 | (~n662 & ~n3295);
  assign n3287 = ~n3288 & n3292 & (~x3 | (~n3289 & (~n698 | ~n1546)));
  assign n3288 = ~x2 & (x0 ? ((x1 & ~x3 & x6) | (~x1 & x3 & x4 & ~x6)) : ((~x4 & ~x6 & x1 & ~x3) | (~x1 & x6 & (x3 ^ x4))));
  assign n3289 = n735 & ((n3290 & n539) | (n538 & n3291));
  assign n3290 = x6 & ~x4 & ~x5;
  assign n3291 = ~x6 & x4 & x5;
  assign n3292 = (~n2328 | n3294) & (~n685 | ~n837) & (n620 | n3293);
  assign n3293 = (~x2 | ~x3 | ~x4 | x0 | ~x1) & (x1 | ((x0 | ~x2 | x3) & (x2 | ((~x0 | (x3 & (x4 | x5))) & (~x4 | ~x5 | x0 | ~x3)))));
  assign n3294 = (~x2 | x4 | ~x5 | ~x6) & (x2 | ~x4 | x5 | x6);
  assign n3295 = (~x3 | ((x0 | ~x1 | x2) & (~x0 | x1 | ~x2 | x4))) & (x1 | ((x0 | x2 | x3 | x4 | ~x5) & (~x0 | ~x2 | ~x4 | (x3 & x5)))) & (x0 | ~x1 | ((x2 | ~x4 | ~x5) & (x4 | x5 | ~x2 | x3)));
  assign n3296 = x2 & ((x0 & ~x1 & ~x3 & ~x4 & ~x6) | (~x0 & ((~x1 & x3 & x4 & ~x6) | (x1 & x6 & (x3 ^ x4)))));
  assign n3297 = n904 & ((~x0 & ~x2 & x4 & ~x5 & x6) | (x5 & ((~x0 & x2 & ~x4 & ~x6) | (x0 & (x2 ? (x4 & x6) : (~x4 & ~x6))))));
  assign z264 = n3299 | ~n3303 | ~n3304 | (x4 & ~n3302);
  assign n3299 = x6 & ((n2328 & ~n3300) | (~x1 & ~n3301));
  assign n3300 = (~x5 | x7 | x2 | ~x4) & (x5 | ~x7 | ~x2 | x4);
  assign n3301 = (~x2 | ((x0 | ~x3 | x4 | x5 | ~x7) & (~x0 | ~x4 | (x3 ? (~x5 | ~x7) : (x5 | x7))))) & (x0 | x2 | x3 | x4 | (x5 ^ x7));
  assign n3302 = (x0 | ~x1 | x2 | x3 | x5 | ~x7) & (x1 | ((~x3 | x5 | ~x7 | x0 | x2) & (x7 | ((x0 | x2 | ~x3 | ~x5) & (~x0 | ~x2 | (~x3 ^ x5))))));
  assign n3303 = x3 ? ((~x2 | ((x0 | ~x7 | (~x1 ^ x4)) & (x4 | x7 | ~x0 | x1))) & (x0 | ~x1 | x7 | (x2 & ~x4))) : ((~x0 | x2 | (x1 ^ x7)) & (~x2 | ((x4 | ~x7 | ~x0 | x1) & (x0 | (x1 ? (~x4 | ~x7) : x7)))));
  assign n3304 = ~n3306 & (x4 | n3307) & (~x3 | x6 | n3305);
  assign n3305 = (x4 | x5 | x7 | x0 | x1 | ~x2) & (~x0 | ((~x1 | x2 | x4 | x5 | ~x7) & (x1 | ~x2 | ~x4 | ~x5 | x7)));
  assign n3306 = ~x2 & x7 & ((~x3 & ~x4 & ~x0 & x1) | (~x1 & (x0 ? (x3 & x4) : (x3 ^ x4))));
  assign n3307 = ((x5 ^ x7) | ((~x2 | x3 | x0 | ~x1) & (x2 | ~x3 | ~x0 | x1))) & (x0 | x1 | ~x5 | (x2 ? (~x3 | ~x7) : (x3 | x7)));
  assign z265 = ~n3309 | ~n3310 | (x2 ? ~n3314 : ~n3313);
  assign n3309 = ((~x2 ^ x4) | (x0 ? (x1 | x3) : (~x1 | ~x3))) & (x0 | ((x2 | ((~x1 | (x4 ? x5 : x3)) & (~x3 | ((~x4 | x5) & (x1 | x4 | ~x5))))) & (x1 | ~x2 | ~x4 | (x3 & ~x5)))) & (~x0 | ((~x4 | ~x5 | x2 | x3) & (x1 | ((~x2 | ((x4 | ~x5) & (~x3 | ~x4 | x5))) & (x4 | ((x3 | ~x5) & (x2 | ~x3 | x5)))))));
  assign n3310 = x2 ? (x3 | n3312) : ((x3 | n3311) & (~n686 | ~n937));
  assign n3311 = (x0 | x1 | x4 | x5 | x6 | ~x7) & ((x1 ? (~x4 | x6) : (x4 | ~x6)) | (x0 ? (x5 | ~x7) : (~x5 | x7)));
  assign n3312 = (~x0 | x1 | ~x4 | x5 | x6 | x7) & (x0 | ((x1 | x4 | ~x5 | ~x6 | ~x7) & (~x1 | ((~x6 | x7 | x4 | x5) & (x6 | ~x7 | ~x4 | ~x5)))));
  assign n3313 = (x1 | ((x0 | x4 | ((x5 | ~x6) & (x3 | ~x5 | x6))) & (~x0 | ~x3 | ~x4 | ~x5 | ~x6))) & (~x0 | ~x1 | x5 | (x3 ? (x4 | x6) : (~x4 | ~x6)));
  assign n3314 = (~x0 | x1 | ~x3 | ~x4 | ~x5 | x6) & (x0 | ((x1 | ~x3 | x4 | x5 | x6) & (~x1 | x3 | (x4 ? (~x5 | ~x6) : (x5 | x6)))));
  assign z266 = ~n3316 | ~n3323 | (~x2 & (~n3321 | (~x7 & ~n3320)));
  assign n3316 = ~n3318 & (~n738 | n3319) & (~x2 | n692 | n3317);
  assign n3317 = (~x4 | x5 | x6 | ~x0 | x1) & (x0 | ((x1 | x4 | ~x5 | ~x6) & (~x1 | (x4 ? (~x5 | x6) : (x5 | ~x6)))));
  assign n3318 = x1 & ((x5 & x6 & ~x0 & x3) | (~x3 & ((x5 & x6 & x0 & ~x2) | (~x0 & ~x5 & (x2 ^ x6)))));
  assign n3319 = (~x5 | x6 | ~x3 | ~x4) & (x2 | ((x3 | ~x4 | ~x6) & (~x3 | x4 | x5 | x6)));
  assign n3320 = (~x0 | ~x1 | ~x3 | x4 | x5 | ~x6) & (x0 | x3 | ~x5 | (x1 ? (~x4 | x6) : (x4 | ~x6)));
  assign n3321 = x1 ? ((x3 | x7 | n3322) & (~x7 | n1019 | x0 | ~x3)) : ((~x3 | ~x7 | n3322) & (x7 | n1019 | ~x0 | x3));
  assign n3322 = (~x0 | ~x4 | x5 | x6) & (x0 | x4 | ~x5 | ~x6);
  assign n3323 = ~n3325 & (x0 | n3324) & (n1115 | n3326);
  assign n3324 = (x1 | x3 | x4 | x5 | ~x6) & (~x1 | ((~x2 | x3 | ~x4 | x5 | ~x6) & (x6 | ((~x3 | x4 | ~x5) & (x2 | ((x4 | ~x5) & (x3 | ~x4 | x5)))))));
  assign n3325 = ~x1 & ((~x6 & ((~x3 & ~x5 & x0 & ~x2) | (~x0 & (x3 ^ x5)))) | (x0 & x6 & ((x3 & ~x5) | (x2 & ~x3 & x5))));
  assign n3326 = (x0 | x1 | ~x4 | ~x6) & (~x0 | x4 | x6 | (x1 ^ ~x2));
  assign z267 = (~x6 & ~n3328) | (x6 & ~n3330) | ~n3332 | (~x2 & ~n3331);
  assign n3328 = (n592 | n928) & (x2 | n3329);
  assign n3329 = (x0 | ~x1 | x3 | ~x4 | ~x5 | x7) & (x4 | ~x7 | ((x0 | x1 | x3 | x5) & (~x0 | (x1 ? (~x3 | x5) : (x3 | ~x5)))));
  assign n3330 = x4 ? (~x7 | (n925 & (x0 | x3 | ~n2306))) : (x7 | (n925 & (~x0 | ~x3 | ~n2306)));
  assign n3331 = (~x4 | ~x5 | x6 | ~x0 | ~x1 | x3) & (x4 | ((x6 | ((~x0 | x1 | x3 | x5) & (x0 | (x1 ? (x3 | ~x5) : (~x3 | x5))))) & (~x0 | ~x6 | (x1 ? x3 : (~x3 | x5)))));
  assign n3332 = (x4 | ((x1 | (x0 ? (~x6 | (~x2 & ~x5)) : (~x5 | x6))) & (x0 | ((~x2 | x5 | x6) & (~x1 | (x5 ^ x6)))))) & (x1 | ~x4 | (x0 ? (~x5 | x6) : (x5 | ~x6)));
  assign z268 = ~n3338 | (~x2 & (n3335 | ~n3337 | (x1 & ~n3334)));
  assign n3334 = (~x0 | ~x3 | x4 | x5 | x7) & (x0 | x3 | ((~x6 | ~x7 | x4 | x5) & (x7 | (x4 ? (~x5 ^ x6) : (~x5 ^ ~x6)))));
  assign n3335 = n605 & ((n545 & n1902) | (x7 & ~n1041 & n3336));
  assign n3336 = x0 & x5;
  assign n3337 = (~x3 | ((x6 | x7 | x1 | x5) & ((~x5 ^ x6) | (x0 ? (x1 | ~x7) : (~x1 | x7))))) & (~x0 | x3 | ((x6 | (x1 ? (~x5 | ~x7) : (~x5 ^ x7))) & (~x1 | x5 | (~x6 & x7))));
  assign n3338 = (x1 | ((~x0 | ((x5 | ~x6 | x7) & (x6 | ~x7 | ~x2 | ~x5))) & (~x2 | x5 | (x6 ^ x7)) & (x0 | (x5 ? (~x6 | x7) : ~x7)))) & (x0 | ((x5 | x6 | ~x7) & (~x1 | ((~x5 | ~x6 | ~x7) & (~x2 | x7 | (~x5 ^ x6))))));
  assign z269 = n3340 | n3342 | ~n3343 | (n724 & (x2 | ~x7));
  assign n3340 = ~x2 & ((n565 & n1489) | (~x7 & n2127 & ~n3341));
  assign n3341 = (~x1 | ~x3 | x4 | x6) & (x1 | x3 | ~x4 | ~x6);
  assign n3342 = n563 & ((n3098 & n738) | (x7 & n664 & ~n783));
  assign n3343 = (x2 | ((~x3 | ~x6 | ~x7 | x0 | ~x1) & (~x0 | x3 | ((~x6 | ~x7) & (~x1 | x6 | x7))))) & (x1 | (x0 ? (x6 ? ~x7 : (x7 | (~x2 & ~x3))) : (~x6 ^ x7)));
  assign z270 = ~n3347 | (~x2 & ((~x6 & ~n3345) | (~x3 & ~n3346)));
  assign n3345 = (x0 | ~x1 | x3 | x4 | ~x5 | ~x7) & (~x0 | ((x1 | x3 | ~x4 | ~x5 | x7) & (~x1 | ~x3 | x4 | x5 | ~x7)));
  assign n3346 = (x0 | ~x1 | x4 | x5 | ~x7) & (~x0 | x1 | ~x4 | (~x5 ^ ~x7));
  assign n3347 = (~x0 | x2 | x3 | (x1 ? ~x7 : (x4 | x7))) & ((~x2 & ~x3) | ((x1 | ~x7) & (x0 | ~x1 | x7))) & (x0 | (x1 ? (~x4 | x7) : ~x7));
  assign z271 = n3349 | ~n3352 | (n3134 & ~n3350) | (x1 & ~n3351);
  assign n3349 = ~x3 & ((x0 & ~x1 & ~x2 & x4 & ~x5) | (~x0 & ((~x4 & x5 & ~x1 & x2) | (x1 & (x2 ? (x4 & x5) : (~x4 & ~x5))))));
  assign n3350 = (x0 | ~x1 | x3 | x4 | ~x5 | ~x6) & (~x0 | ((x1 | x3 | ~x4 | ~x5 | x6) & (~x1 | ~x3 | x4 | x5 | ~x6)));
  assign n3351 = (~x0 | x2 | ~x3 | x4 | x5 | x6) & (x0 | x3 | ((x5 | ~x6 | ~x2 | ~x4) & (~x5 | x6 | x2 | x4)));
  assign n3352 = (~x0 | x2 | x3 | (~x1 & x4)) & (~x2 | ((~x3 | (x0 & x1)) & (x0 | x1 | (~x4 & ~n837))));
  assign z272 = ~n3354 | ~n3357;
  assign n3354 = (x2 | n3355) & (~x3 | ~x7 | n3356 | x0 | ~x2);
  assign n3355 = (~x1 | ((~x0 | ((x3 | ~x5) & (x5 | x6 | ~x3 | x4))) & (x3 | x4 | (x6 ? x5 : x0)))) & (~x0 | x3 | (x5 ? x4 : (x1 & ~x4))) & (~x3 | ((x0 | x1 | (~x5 & ~x6)) & (~x4 | (x0 & (x1 | ~x5 | ~x6)))));
  assign n3356 = (~x5 | x6 | x1 | x4) & (x5 | ~x6 | ~x1 | ~x4);
  assign n3357 = (~x2 | n3358) & (x7 | ((~n1546 | ~n921) & (x2 | n3350)));
  assign n3358 = (x0 | ((~x1 | x3 | (x4 & (x5 | x6))) & (~x3 | ((~x4 | ~x5) & (x1 | (~x4 & (~x5 | ~x6))))))) & (x1 | x3 | (~x0 & (x4 | x5 | x6)));
  assign z273 = ~n3363 | (~x5 & (~n3362 | (x1 ? ~n3360 : ~n3361)));
  assign n3360 = (x0 | ~x2 | x3 | x4 | x6 | ~x7) & (~x6 | (x0 ? (x2 | (x3 ? (x4 | x7) : (~x4 | ~x7))) : (~x2 | ~x3 | (~x4 ^ x7))));
  assign n3361 = (~x0 | ~x2 | ~x3 | ~x4 | x6 | ~x7) & (x0 | x3 | ((x6 | ~x7 | x2 | ~x4) & (~x2 | x4 | ~x6 | x7)));
  assign n3362 = (x6 | ((~x2 | x3 | x4 | x0 | x1) & (~x3 | ((~x0 | ~x1 | x2 | x4) & (x0 | (x1 ? (~x2 | ~x4) : (x2 | x4))))))) & (x0 | x1 | x2 | ~x4 | ~x6);
  assign n3363 = n3367 & ~n3368 & ~n3369 & (~x5 | (~n3364 & ~n3366));
  assign n3364 = ~x2 & ~n3365;
  assign n3365 = x0 ? (x1 | x6 | (x3 ? (x4 | ~x7) : (~x4 | x7))) : (~x1 | x3 | ~x6 | (x4 ^ x7));
  assign n3366 = ~x4 & n538 & ((n1317 & n540) | (n537 & n610));
  assign n3367 = (x0 | (x1 ? (x4 | (x5 ? (~x2 & ~x3) : x2)) : ((x2 | ~x4 | ~x5) & (x4 | x5 | ~x2 | ~x3)))) & (x3 | ~x4 | ~x5 | ~x0 | ~x1 | x2) & (x1 | ((~x0 | x2 | x3 | x4 | ~x5) & (~x4 | ((~x2 | ~x5 | (~x0 & x3)) & (~x0 | x5 | (x2 & x3))))));
  assign n3368 = ~n1041 & (x2 ? (n664 & n916) : (n985 & n738));
  assign n3369 = ~n2111 & (x3 ? (n538 & n641) : (n539 & n642));
  assign z274 = ~n3374 | n3380 | ~n3381 | (~x2 & (~n3371 | ~n3379));
  assign n3371 = (n800 | n3372) & (~x6 | n3373);
  assign n3372 = (x0 | ~x1 | x3 | ~x4 | ~x6) & (~x0 | x1 | x6 | (~x3 ^ x4));
  assign n3373 = (~x0 | ~x1 | ~x3 | x4 | x5 | x7) & (x0 | ((~x4 | ~x5 | ~x7 | x1 | ~x3) & (~x1 | x4 | (x3 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n3374 = ~n3375 & ~n3376 & ((x3 & ~n641) | n3378 | (~x3 & ~n642));
  assign n3375 = ~n1099 & (x0 ? ((x1 & ~x2 & ~x5 & ~x6) | (~x1 & (x2 ? x5 : (~x5 & x6)))) : ((x1 & ~x2 & x5 & ~x6) | (~x5 & x6 & ~x1 & x2)));
  assign n3376 = ~n846 & ~n3377;
  assign n3377 = (x2 | x3 | x4 | ~x0 | ~x1) & (x0 | ((x1 | x2 | ~x3 | x4) & (x3 | ~x4 | ~x1 | ~x2)));
  assign n3378 = (x2 | ~x5 | x0 | ~x1) & (x1 | (x0 ? (~x2 ^ ~x5) : (~x2 | x5)));
  assign n3379 = (((x5 | ~x6 | x3 | x4) & (~x5 | x6 | ~x3 | ~x4)) | (x0 ^ ~x1)) & (x0 | ((~x3 | ((~x5 | ~x6 | ~x1 | x4) & (x5 | x6 | x1 | ~x4))) & (x1 | x3 | ~x5 | (x4 & ~x6))));
  assign n3380 = n616 & (x1 ? ((~x3 & ~x4 & x5 & x6) | (x3 & ~x5 & ~x6)) : (x4 & ~x6 & (~x3 ^ x5)));
  assign n3381 = (n824 | n3382) & (~x2 | (~n3383 & (~n1743 | ~n762)));
  assign n3382 = (~x4 | ((~x0 | ((x3 | ~x6 | ~x1 | x2) & (~x3 | x6 | x1 | ~x2))) & (x0 | x1 | x2 | x3 | x6))) & (x0 | ~x1 | ~x2 | x4 | (x3 ^ x6));
  assign n3383 = n2512 & ((x0 & ~x3 & x6 & ~n800) | (~x0 & (x3 ? (~x6 & ~n800) : n767)));
  assign z275 = ~n3387 | ~n3394 | (~n662 & ~n3385) | (~x0 & ~n3386);
  assign n3385 = (~x2 | x3 | x4 | x0 | ~x1) & (x1 | ~x3 | x5 | (x0 ? (x2 ^ x4) : (~x2 | x4)));
  assign n3386 = x1 ? ((x2 | x3 | x4 | x5 | x6) & (~x3 | ~x6 | (x2 ? (~x4 | ~x5) : (~x4 ^ x5)))) : ((~x2 | x3 | x4 | ~x5 | ~x6) & (x2 | ~x3 | ~x4 | x5 | x6));
  assign n3387 = ~n3388 & ~n3390 & ~n3392 & n3393 & (x1 | n3389);
  assign n3388 = ~x6 & ((~x0 & x2 & x4 & (x1 ^ x3)) | (~x2 & ((x0 & (x1 ? (~x3 & ~x4) : (x3 & x4))) | (x3 & ~x4 & ~x0 & ~x1))));
  assign n3389 = (~x5 | ~x6 | ~x7 | ~x2 | ~x3 | x4) & (x2 | x3 | ~x4 | ((x6 | x7) & (x5 | ~x6 | ~x7)));
  assign n3390 = n3391 & ((n597 & n563) | (x2 & ~n2500));
  assign n3391 = x6 & x0 & ~x1;
  assign n3392 = (n586 | n1743) & ((n1901 & n2326) | (n2327 & n1902));
  assign n3393 = (~n1082 | ~n1621) & (x3 | ~x6 | ~n598 | n1204);
  assign n3394 = ~n3396 & (n620 | n3395);
  assign n3395 = x2 ? ((x4 | x5 | x1 | x3) & ((x4 & x5) | (x0 ? (x1 | x3) : (~x1 | ~x3)))) : ((~x1 | (x3 ? (x4 | x5) : ~x4)) & (x0 | ~x5 | (x1 ? x3 : (~x3 | ~x4))));
  assign n3396 = ~x1 & ((x5 & ~n3397) | (x0 & n1812 & n678));
  assign n3397 = x0 ? ((~x2 | ~x3 | ~x4 | x6 | x7) & (x2 | x4 | (x3 ? (x6 | x7) : (~x6 | ~x7)))) : ((x2 | x3 | ~x4 | ~x6 | ~x7) & (~x2 | ~x3 | x4 | x6 | x7));
  assign z276 = n3404 | ~n3405 | (x1 ? ~n3399 : (n3401 | ~n3402));
  assign n3399 = x0 ? (~n563 | ~n762) : n3400;
  assign n3400 = (~x3 | (~x6 ^ x7) | (x2 ? (x4 | x5) : (~x4 | ~x5))) & (x2 | x3 | ((~x6 | ~x7 | x4 | ~x5) & (x5 | ((x6 | ~x7) & (~x4 | ~x6 | x7)))));
  assign n3401 = ~n927 & ((x3 & ~x5 & ~x6 & ~x0 & ~x2) | (x2 & ((x5 & ~x6 & ~x0 & ~x3) | (x0 & x6 & (x3 ^ ~x5)))));
  assign n3402 = (x6 | n3403) & (~n651 | n692 | ~x6 | ~n1449);
  assign n3403 = (x2 | x3 | x4 | ~x5 | ~x7) & (x0 | ~x2 | ~x3 | ~x4 | x5 | x7);
  assign n3404 = ~n592 & ((x0 & ((x3 & ~x5 & ~x1 & x2) | (x1 & ~x2 & ~x3 & x5))) | (~x1 & ~x2 & ((~x3 & ~x5) | (~x0 & x3 & x5))));
  assign n3405 = ~n3407 & ~n3408 & ~n3409 & n3410 & (x0 | n3406);
  assign n3406 = x2 ? (x1 ? (~x5 | ((~x4 | ~x7) & (~x3 | x4 | x7))) : (x5 | ((x4 | x7) & (x3 | ~x4 | ~x7)))) : ((x1 | ~x3 | x4 | x5 | ~x7) & (x7 | ((x3 | ~x4 | ~x5) & (~x1 | (x3 ? (x4 | x5) : ~x5)))));
  assign n3407 = ~x1 & x3 & ((x4 & x7 & ~x0 & x2) | (x0 & ~x2 & (~x4 ^ x7)));
  assign n3408 = ~n906 & (x0 ? ((~x1 & x2 & x4 & x5) | (x1 & ~x2 & ~x4 & ~x5)) : (x2 & (x1 ? (x4 & ~x5) : (~x4 & x5))));
  assign n3409 = ~n627 & ((~x7 & n738 & x2 & ~x3) | (~x2 & x3 & x7 & n664));
  assign n3410 = x3 | x7 | (x4 ? (~x5 | ~n534) : ~n750);
  assign z277 = ~n3416 | (x0 ? ~n3414 : (n3413 | (x1 & ~n3412)));
  assign n3412 = (x2 | x3 | x4 | x5 | ~x6 | ~x7) & (x7 | (x2 ? ((~x3 | x4 | ~x5 | ~x6) & (x3 | (x4 ? (~x5 | x6) : (x5 | ~x6)))) : ((x3 | ~x5 | ~x6) & (x5 | x6 | ~x3 | ~x4))));
  assign n3413 = n1599 & (((x2 ^ x6) & (x3 ? (x4 & ~x5) : (~x4 & x5))) | (~x5 & ~x6 & ~x2 & ~x4) | (x4 & x5 & x6 & x2 & ~x3));
  assign n3414 = x1 ? (~n563 | ~n1166) : n3415;
  assign n3415 = ((x4 ^ x6) | ((x2 | x3 | x5 | x7) & (~x2 | ~x7 | (x3 ^ x5)))) & (x2 | ~x5 | ~x7 | (x3 ? (x4 | ~x6) : (~x4 | x6)));
  assign n3416 = ~n3417 & n3419 & (x4 | n1014) & (~x2 | n3418);
  assign n3417 = ~n912 & (x1 ? ((~x2 & ~x3 & x4) | (x3 & ~x4 & ~x0 & x2)) : ((x0 & x2 & ~x3 & ~x4) | (~x0 & x3 & (~x2 ^ x4))));
  assign n3418 = (x0 | ~x1 | x3 | x4 | x5 | x6) & (x1 | (x4 ? (x5 | x6) : (~x5 | ~x6)) | (x0 ^ x3));
  assign n3419 = ~n3420 & (x2 | n3421);
  assign n3420 = x4 & ((~x0 & x1 & x2 & (~x3 ^ x5)) | (~x1 & (x0 ? (x2 ? (~x3 & x5) : (x3 & ~x5)) : (~x2 & (~x3 ^ x5)))));
  assign n3421 = (~x5 | ((x3 | ~x6 | ~x0 | x1) & (x0 | ~x1 | (x3 ? (~x4 | ~x6) : (x4 | x6))))) & (~x0 | x1 | x5 | x6 | (~x3 ^ x4));
  assign z278 = ~n3424 | n3432 | (n545 & ~n3434) | (~x3 & ~n3423);
  assign n3423 = (x1 | ((~x4 | ((x5 | ~x6 | x0 | ~x2) & (~x0 | ~x5 | (x2 & x6)))) & (x0 | x4 | (x2 ? (x5 ^ x6) : (x5 | ~x6))))) & (x0 | ~x1 | (x4 ? (x2 ? (x5 ^ x6) : (x5 | ~x6)) : (~x5 | x6)));
  assign n3424 = n3427 & (n592 | n3426) & (~x3 | n3425);
  assign n3425 = x0 ? (x1 | ((x5 | ~x6 | x2 | x4) & (~x2 | (x4 ? (x5 | ~x6) : (x5 ^ x6))))) : ((x1 | x2 | ~x4 | ~x5 | x6) & (~x1 | ~x2 | x4 | x5 | ~x6));
  assign n3426 = x0 ? (x1 | (x3 ? (~x5 | (~x2 ^ x6)) : (x5 | x6))) : ((~x2 | ((~x1 | ~x6 | (~x3 ^ ~x5)) & (~x5 | x6 | x1 | x3))) & (x1 | x2 | (x3 ? (x5 | x6) : (~x5 | ~x6))));
  assign n3427 = ~n3430 & n3431 & (n1465 | n1957) & (n3428 | n3429);
  assign n3428 = (x3 | x5) & (~x2 | ~x3 | ~x5);
  assign n3429 = (x4 | x6 | x7 | x0 | ~x1) & (~x4 | ~x6 | ~x7 | ~x0 | x1);
  assign n3430 = ~x1 & x2 & ~x4 & (x0 ? (~x3 & x6) : (x3 & ~x6));
  assign n3431 = ((x1 ^ ~x6) | ((x3 | x4 | ~x0 | x2) & (x0 | ~x3 | (x2 ^ x4)))) & (x2 | ~x4 | (x0 ? (x1 ? (x3 | ~x6) : (~x3 | x6)) : (x1 ? (~x3 | ~x6) : (x3 | x6))));
  assign n3432 = ~x4 & ((~x7 & ~n3433) | (~x3 & n537 & n975));
  assign n3433 = (x1 | (~x0 ^ ~x3) | (x2 ? (x5 | ~x6) : (~x5 | x6))) & (~x3 | x5 | x6 | ~x0 | ~x1 | x2);
  assign n3434 = (~x1 | x2 | x3 | ~x5 | x6 | x7) & (~x7 | ((x1 | x2 | ~x3 | x5 | ~x6) & (x3 | ~x5 | (x1 ? (~x2 ^ x6) : (~x2 | ~x6)))));
  assign z279 = ~n3439 | ~n3445 | (x1 ? ~n3436 : ~n3438);
  assign n3436 = x0 ? (~n665 | ~n698) : n3437;
  assign n3437 = x3 ? (x2 ? ((x6 | x7 | x4 | x5) & (~x6 | ~x7 | ~x4 | ~x5)) : (x4 ? (x5 ? (~x6 | x7) : (x6 | ~x7)) : (x7 | (~x5 ^ x6)))) : ((x2 | x4 | x5 | x6 | ~x7) & (~x6 | ((x5 | x7 | x2 | ~x4) & (~x2 | (x4 ? (x5 | ~x7) : (~x5 | x7))))));
  assign n3438 = x3 ? (x0 ? ((x5 | x7 | x2 | x4) & (~x5 | ~x7 | ~x2 | ~x4)) : ((x5 | x7 | ~x2 | x4) & (x2 | (x4 ? (x5 | ~x7) : (~x5 | x7))))) : ((~x4 | ~x5 | ~x7 | x0 | ~x2) & (~x0 | ((~x2 | x4 | ~x5 | x7) & (~x4 | x5 | ~x7))));
  assign n3439 = n3440 & ~n3442 & ~n3443 & (x3 | n3444);
  assign n3440 = (n620 | n3441) & (~x3 | n1019 | ~n2758);
  assign n3441 = (x3 | (x0 ? (x2 | x5) : (~x2 | ~x5)) | (x1 ^ x4)) & (x1 | ~x2 | ~x3 | (x0 ? (x4 | ~x5) : (~x4 | x5)));
  assign n3442 = ~n1862 & (x1 ? (~x2 & (x0 ? (~x3 & x5) : (x3 ^ ~x5))) : ((x3 & x5 & ~x0 & x2) | ((x2 ^ x5) & (x0 ^ ~x3))));
  assign n3443 = ~n783 & (x0 ? ((x3 & ~x5 & ~x1 & x2) | (x1 & ~x2 & ~x3 & x5)) : (~x1 & x2 & (x3 ^ ~x5)));
  assign n3444 = (x0 | ~x1 | ~x2 | ~x4 | x5 | x6) & (~x0 | x1 | x2 | ~x5 | (~x4 ^ x6));
  assign n3445 = x1 ? n3447 : ((n3446 | n856) & (x2 | n3448));
  assign n3446 = x0 ? (~x2 | x3) : (x2 | ~x3);
  assign n3447 = (~x0 | x2 | x3 | x4 | x5 | x7) & (x0 | ((~x2 | ~x3 | (x4 ? (x5 | x7) : (~x5 | ~x7))) & (x3 | ((x5 | ~x7 | ~x2 | x4) & (x2 | ~x5 | (x4 ^ x7))))));
  assign n3448 = (~x6 | ((x0 | x3 | x5 | x7) & (~x4 | ((~x5 | ~x7 | x0 | x3) & (~x0 | ~x3 | (x5 ^ x7)))))) & (x4 | ~x5 | x6 | (x0 ? (x3 ^ x7) : (x3 | ~x7)));
  assign z280 = ~n3454 | ~n3460 | (~n662 & ~n3450) | (~x0 & ~n3451);
  assign n3450 = x1 ? (~x5 | ((x3 | x4 | ~x0 | x2) & (x0 | ~x2 | (~x3 ^ ~x4)))) : ((~x3 | x4 | ~x5 | x0 | ~x2) & (~x4 | ((~x3 | ~x5 | x0 | x2) & (~x0 | (x2 ? (x3 | ~x5) : (~x3 | x5))))));
  assign n3451 = ~n3452 & (~n808 | ((~x3 | x5 | x6 | x7) & (x3 | ~x6 | (~x5 ^ x7))));
  assign n3452 = ~x1 & ((n1902 & n3453) | (x2 & x3 & ~n2351));
  assign n3453 = x4 & ~x2 & ~x3;
  assign n3454 = ~n3457 & ~n3459 & (x3 ? n3455 : (~n651 | n3456));
  assign n3455 = x0 ? (x1 | ((x5 | ~x6 | x2 | x4) & (~x5 | (x2 ? (x4 ^ x6) : (~x4 | x6))))) : ((~x4 | x5 | (x1 ? (~x2 | ~x6) : (~x2 ^ x6))) & (~x1 | x4 | ~x5 | (~x2 ^ ~x6)));
  assign n3456 = (~x5 | x6 | x7 | ~x1 | ~x4) & (x1 | ((~x4 | x5 | ~x6 | ~x7) & (x6 | x7 | x4 | ~x5)));
  assign n3457 = ~n1031 & ~n3458;
  assign n3458 = (~x2 | x5 | x6 | x7) & (x2 | ~x5 | ~x6 | ~x7);
  assign n3459 = ~n1429 & (n1954 | (x3 & n897 & ~n885));
  assign n3460 = (n620 | n3461) & (x3 | n3462);
  assign n3461 = x0 ? ((x1 | ((~x2 | (x3 ? (~x4 | x5) : x4)) & (x3 | (x4 ? x2 : ~x5)))) & (x2 | ((x3 | ~x4 | ~x5) & (x4 | x5 | ~x1 | ~x3)))) : ((x5 | ((x3 | ~x4 | x1 | ~x2) & (~x1 | x4 | (~x2 ^ ~x3)))) & (~x3 | (x1 ? (x2 | ~x4) : (x2 ? (~x4 | ~x5) : x4))));
  assign n3462 = (x5 | ((~x6 | (x0 ? (x1 ? (x2 | x4) : (~x2 | ~x4)) : (x1 ? (~x2 ^ x4) : (x2 | x4)))) & (~x0 | x2 | x6 | (x1 ^ x4)))) & (x0 | ~x5 | ((~x4 | x6 | ~x1 | ~x2) & (x1 | (x2 ? (x4 ^ x6) : (~x4 | x6)))));
  assign z281 = n3464 | n3466 | ~n3470 | (~n620 & ~n3469);
  assign n3464 = x1 & ((n1415 & n698) | (~x0 & ~n3465));
  assign n3465 = x7 ? ((~x4 | ((~x3 | (x2 ? (x5 | x6) : (~x5 | ~x6))) & (~x2 | x3 | (~x5 ^ x6)))) & (x2 | x4 | ((x5 | ~x6) & (x3 | ~x5 | x6)))) : ((~x2 | x6 | (x3 ? (x4 | ~x5) : (~x4 | x5))) & (x2 | ~x3 | ~x4 | x5 | ~x6));
  assign n3466 = ~x1 & (x3 ? ~n3468 : ~n3467);
  assign n3467 = (~x6 | (x2 ? (x4 | (x0 ? (x5 ^ x7) : (x5 | ~x7))) : (~x4 | ((x5 | ~x7) & (~x0 | ~x5 | x7))))) & (x0 | ~x2 | x6 | (x4 ? (~x5 | x7) : (x5 ^ x7)));
  assign n3468 = (~x0 | ~x2 | ~x4 | ~x5 | x6 | x7) & (x4 | ((x5 | ~x6 | x7 | x0 | x2) & ((x6 ^ x7) | (x0 ? (~x2 | x5) : (x2 | ~x5)))));
  assign n3469 = (~x1 | x2 | x3 | ~x4 | ~x5) & (x1 | ((x0 | ~x2 | ~x3 | (x4 ^ x5)) & (x2 | x4 | ~x5 | (~x0 & x3))));
  assign n3470 = ~n3471 & n3472 & (~n897 | n3475) & (~x2 | n3474);
  assign n3471 = ~n592 & ((x3 & x5 & ~x0 & x1) | (~x1 & ~x2 & ~x5 & (x0 | ~x3)));
  assign n3472 = x0 ? (x3 ? n3473 : (n1002 | (x1 ^ ~x2))) : ((~x3 | n1002 | x1 | ~x2) & (x3 | n3473));
  assign n3473 = (x4 | x5 | x7 | ~x1 | x2) & (x1 | ~x4 | ((~x5 | ~x7) & (~x2 | x5 | x7)));
  assign n3474 = (~x5 | ((x0 | ~x1 | x3 | x4 | x7) & (~x0 | x1 | (x3 ? (x4 | ~x7) : (~x4 | x7))))) & (x0 | ~x1 | x4 | x5 | (~x3 ^ x7));
  assign n3475 = (x1 | ~x3 | ~x4 | ~x5 | x7) & (x5 | ((x1 | ~x3 | ~x4 | ~x7) & (~x1 | (x3 ? (x4 | x7) : (~x4 | ~x7)))));
  assign z282 = n3480 | ~n3482 | ~n3483 | (~x1 & (~n3477 | ~n3481));
  assign n3477 = ~n3479 & (x5 | n3478) & (~n1317 | n2587 | ~x5 | x7);
  assign n3478 = (x0 | ~x2 | ~x3 | ~x4 | ~x6 | x7) & (x3 | x6 | ((x4 | ~x7 | x0 | x2) & (~x0 | (x2 ? (x4 | ~x7) : (~x4 | x7)))));
  assign n3479 = ~n1041 & (x3 ? (n651 & n691) : (n723 & n616));
  assign n3480 = ~n846 & (x2 ? ((~x1 & x3 & x4) | (~x0 & (x1 ? (x3 & ~x4) : x4))) : ((x0 & ~x1 & ~x4) | (x1 & ~x3 & x4)));
  assign n3481 = x0 ? (~x2 | x3 | x5 | (~x4 ^ x6)) : (x2 | ~x5 | ((x4 | ~x6) & (~x3 | ~x4 | x6)));
  assign n3482 = (x4 | ~x5 | x6 | ~x1 | x2 | x3) & (x1 | ((x2 | x3 | ~x4 | ~x5 | x6) & (~x2 | ~x3 | x4 | x5 | ~x6)));
  assign n3483 = ~n3484 & ~n3487 & (x4 ? (x7 ? n3486 : n3485) : (x7 ? n3485 : n3486));
  assign n3484 = ~n2465 & ((x0 & ~x1 & x4 & n1121) | (~x0 & (x1 ? (x4 ? n1120 : n1121) : (~x4 & n1120))));
  assign n3485 = (x0 | ~x3 | x6 | (x1 ? (~x2 | ~x5) : (x2 | x5))) & (x3 | ~x6 | ((~x1 | x2 | x5) & (~x0 | x1 | ~x2 | ~x5)));
  assign n3486 = (x0 | ~x1 | ((x2 | ~x3 | x5 | x6) & (~x5 | ~x6 | ~x2 | x3))) & (x1 | ((x5 | ~x6 | x2 | x3) & (~x0 | ~x2 | ~x3 | ~x5 | x6)));
  assign n3487 = x1 & ((n559 & n2314) | (~x0 & ~n3488));
  assign n3488 = ((~x4 ^ ~x5) | ((~x6 | ~x7 | x2 | ~x3) & (x6 | x7 | ~x2 | x3))) & (~x2 | ~x3 | ~x4 | x5 | ~x6 | ~x7);
  assign z283 = ~n3491 | ~n3497 | (~n800 & ~n3490);
  assign n3490 = x3 ? ((~x4 | x6 | x0 | x2) & (~x2 | ~x6 | ((x1 | ~x4) & (x0 | (x1 & ~x4))))) : (x4 | (x0 ? (x1 ? (x2 | ~x6) : (~x2 | x6)) : (x1 ? (~x2 | x6) : (x2 | ~x6))));
  assign n3491 = n3495 & (~n1122 | n3494) & (x2 | (n3492 & n3493));
  assign n3492 = ((x0 ? (x3 | ~x4) : (~x3 | x4)) | ((~x5 | x7) & (~x1 | x5 | ~x7))) & (x0 | ((~x1 | x4 | ~x5 | x7) & (x1 | x3 | ~x4 | x5 | ~x7))) & (x1 | ((x3 | ~x4 | ~x5 | x7) & (~x0 | ~x3 | x4 | x5 | ~x7)));
  assign n3493 = (~x1 | x3 | x5 | x6 | x7) & (~x5 | ~x6 | ~x7 | x0 | ~x3);
  assign n3494 = (~x0 | x1 | x2 | x5) & (x0 | ~x1 | (~x2 ^ ~x5));
  assign n3495 = ~n3496 & (~x2 | n857 | (~n1079 & (~n543 | ~n985)));
  assign n3496 = x0 & ~x1 & x3 & ~x7 & (x2 ^ x5);
  assign n3497 = x2 ? (n3500 & n3501) : (x1 ? n3498 : n3499);
  assign n3498 = (x5 | x6 | ~x7 | ~x0 | ~x3 | x4) & (~x5 | ~x6 | x7 | x0 | x3 | ~x4);
  assign n3499 = (x7 | (x0 ? (x4 | ((x5 | x6) & (x3 | ~x5 | ~x6))) : (~x4 | x5 | (x3 ^ x6)))) & (~x3 | ~x7 | ((x5 | x6 | x0 | x4) & (~x0 | ~x4 | (~x5 ^ ~x6))));
  assign n3500 = (x0 | ~x3 | x4 | x5 | x7) & (x1 | x3 | ((~x5 | ~x7 | ~x0 | ~x4) & (x0 | (x4 ? (x5 | x7) : (~x5 | ~x7)))));
  assign n3501 = (~x0 | x1 | x3 | ~x5 | n1862) & (x0 | ((x1 | n3502) & (x5 | n1862 | ~x1 | ~x3)));
  assign n3502 = (x3 | x4 | x5 | ~x6 | x7) & (x6 | (x3 ? (x4 ? (x5 | x7) : (~x5 | ~x7)) : (~x5 | (x4 ^ x7))));
  assign z284 = (~n662 & ~n3504) | (~x3 & ~n3505) | ~n3507 | (x3 & ~n3506);
  assign n3504 = (~x3 | ~x4 | ~x5 | x0 | x1 | ~x2) & (x3 | ((x1 | ((~x0 | (x2 ^ x4)) & (x4 | (x2 ? x0 : ~x5)))) & (~x1 | x5 | ((x2 | ~x4) & (x0 | (x2 & ~x4)))) & (x4 | ~x5 | (~x0 ^ x2))));
  assign n3505 = (x4 | x6 | ((x0 | ~x1 | ~x2 | x5) & (~x0 | (x1 ? (x2 | x5) : ~x2)))) & (~x6 | ((x0 | ~x1 | x2 | ~x5) & (~x4 | ((x0 | x2 | ~x5) & ((x0 & x2) | (x1 ^ x5))))));
  assign n3506 = (x1 | ((x5 | x6 | x0 | ~x4) & (~x0 | x4 | ~x6 | (x2 & x5)))) & (x0 | ((x2 | ~x4 | ~x5 | x6) & (~x1 | ((x5 | ~x6 | x2 | x4) & (~x4 | ~x5 | x6)))));
  assign n3507 = (x0 & (x6 ? n3509 : ~n3512)) | (x6 & n3508 & n3509) | (~x6 & n3511 & ~n3512);
  assign n3508 = (x1 | ~x2 | x3 | ~x4 | ~x5 | x7) & (x4 | ((~x1 | ((~x3 | ~x5 | x7) & (~x2 | x3 | x5 | ~x7))) & (~x5 | x7 | x2 | ~x3) & (x1 | x5 | ((~x3 | x7) & (x2 | x3 | ~x7)))));
  assign n3509 = (x2 | ((~x4 | n3510) & (~n669 | ~n691 | ~x1 | x4))) & (~x2 | x4 | n3510) & (~n669 | ~n691 | x1 | ~x4);
  assign n3510 = (~x3 | x5 | x7 | x0 | ~x1) & (~x0 | x1 | ~x5 | (~x3 ^ x7));
  assign n3511 = x4 ? ((~x1 | ((~x3 | x5 | ~x7) & (x2 | x3 | ~x5 | x7))) & (x1 | x2 | x3 | x5 | x7)) : (~x7 | ((~x3 | ~x5) & (x1 | (~x3 & (x2 | x5)))));
  assign n3512 = n1021 & ((x4 & x7) | (n691 & n1148));
  assign z285 = ~n3516 | (x4 & (x2 ? ~n3514 : (~x7 & ~n3515)));
  assign n3514 = (x1 | ~x5 | (x0 ? (x3 ? (x6 | x7) : (~x6 | ~x7)) : ((~x6 | x7) & (x3 | x6 | ~x7)))) & (x0 | ~x1 | x5 | ((~x6 | ~x7) & (~x3 | x6 | x7)));
  assign n3515 = (x0 | ~x1 | x3 | ~x5 | x6) & (x1 | ((x5 | x6 | x0 | x3) & (~x0 | ~x6 | (~x3 ^ x5))));
  assign n3516 = x4 ? n3519 : (n3520 & (x2 ? n3518 : n3517));
  assign n3517 = x1 ? (x0 ? ((x3 | ~x5 | ~x6 | x7) & (x6 | ~x7 | ~x3 | x5)) : (~x5 | (x3 ? (~x6 | x7) : (x6 | ~x7)))) : (x5 | ((x0 | ((~x6 | x7) & (x3 | x6 | ~x7))) & (x7 | ((x3 | ~x6) & (~x0 | ~x3 | x6)))));
  assign n3518 = (((x6 | ~x7) & (~x3 | ~x6 | x7)) | (x0 ? (x1 | ~x5) : (~x1 | x5))) & (x0 | x1 | ~x5 | ((~x6 | ~x7) & (~x3 | x6 | x7)));
  assign n3519 = (x1 | ((x2 | ((x3 | x5 | ~x7) & (~x5 | x7 | ~x0 | ~x3))) & (x5 | (x0 ? (~x2 | x7) : ~x7)) & (~x0 | ~x2 | (x3 ? (~x5 | ~x7) : x7)))) & (~x5 | ~x7 | x0 | x2) & (~x1 | (x5 ? (~x7 | (x0 & (x2 | x3))) : (x7 | ((x2 | x3) & (x0 | (x2 & x3))))));
  assign n3520 = x2 ? ((x1 | x5 | (x0 ^ x7)) & (x0 | ~x5 | x7 | (~x1 & x3))) : (x7 ? ((~x3 | x5 | x0 | ~x1) & (~x0 | (x1 ? (x3 | x5) : ~x3))) : ((x1 | x3 | ~x5) & (x0 | (x1 ? (x3 | x5) : ~x5))));
  assign z286 = (x4 & ~n3522) | (~x2 & ~n3524) | ~n3528 | (~x4 & ~n3525);
  assign n3522 = (x6 | n3523) & (x3 | x5 | ~x6 | ~n616 | n1100);
  assign n3523 = (x0 | ~x1 | ~x5 | (x2 ? (~x3 | ~x7) : (x3 | x7))) & (x1 | ((x0 | x2 | x3 | ~x5 | ~x7) & (x7 | ((~x0 | ~x3 | (x2 ^ x5)) & (x3 | x5 | x0 | x2)))));
  assign n3524 = (~x6 & ((~x0 & (~x3 | (~x4 & ~x5))) | (~x4 & (~x3 | (x0 & x5))))) | (x1 & x5) | (~x5 & (~x1 | (x0 & x3 & (x4 | x6))));
  assign n3525 = ~n3527 & (x7 | n3526) & (x3 | ~n897 | ~n836);
  assign n3526 = (x0 | x1 | x2 | ~x3 | x5 | x6) & (~x0 | ~x6 | ((~x1 | x2 | ~x3 | x5) & (x3 | ~x5 | x1 | ~x2)));
  assign n3527 = ~n824 & ((x0 & ~x1 & ~x2 & ~x6) | (~x0 & x1 & x2 & ~x3 & x6));
  assign n3528 = (n800 | n3530) & (~x2 | n3529);
  assign n3529 = x6 ? ((x1 | ~x3 | x5) & (x0 | ~x1 | ~x5 | (~x3 & ~x4))) : ((x0 | ~x1 | x5) & (x1 | ~x5 | (x3 & x4)));
  assign n3530 = (x0 | ~x3 | x6 | (x1 ? (x2 | x4) : (~x2 | ~x4))) & (x3 | ((~x0 | ((~x4 | ~x6 | x1 | ~x2) & (~x1 | x2 | x4 | x6))) & (x0 | x1 | ~x2 | x4 | ~x6)));
  assign z287 = ~n3536 | (x1 ? ~n3532 : (n3535 | (x2 & ~n3534)));
  assign n3532 = x0 ? (~n665 | ~n686) : n3533;
  assign n3533 = x4 ? (x5 | ((x6 | ~x7 | x2 | x3) & (~x2 | (x3 ? (x6 | ~x7) : (~x6 | x7))))) : ((~x5 | ((x2 | ~x6 | x7) & (x6 | ~x7 | ~x2 | x3))) & (x2 | x3 | x5 | (x6 ^ x7)));
  assign n3534 = x3 ? (~x7 | ((x0 | x4 | ~x5 | ~x6) & (~x0 | ~x4 | (~x5 ^ ~x6)))) : ((~x5 ^ x6) | (x0 ? (x4 | ~x7) : (~x4 | x7)));
  assign n3535 = n3134 & (x0 ? ((~x5 & ~x6 & x3 & x4) | (~x3 & x6 & (x4 ^ x5))) : (~x4 & (x3 ? (x5 ^ ~x6) : (x5 & ~x6))));
  assign n3536 = ~n3538 & n3540 & (x3 ? (x1 | n3539) : n3537);
  assign n3537 = (x1 | ((~x0 | ~x6 | (x2 ? x7 : (~x4 | ~x7))) & (x6 | ~x7 | (x4 ? ~x2 : x0)))) & (x0 | ~x2 | (x4 ? (x6 | ~x7) : (~x6 | x7)));
  assign n3538 = ~n662 & ((~x0 & x4 & (x2 ^ ~x3)) | (~x2 & ~x4 & (x3 ? ~n857 : x0)));
  assign n3539 = (~x4 | x6 | x7 | ~x0 | ~x2) & (x0 | x2 | x4 | ~x6 | ~x7);
  assign n3540 = (x3 | ~x4 | ~x6 | ~x0 | ~x1 | x2) & (~x3 | (x0 & x1) | (x2 ? (x4 | x6) : (~x4 | ~x6)));
  assign z288 = n3542 | ~n3543 | n3544 | n3548 | (~x1 & ~n3547);
  assign n3542 = n664 & ((~x2 & ~x3 & ~x4 & x5 & x7) | (~x7 & (x2 ? (x3 ? (x4 & x5) : (x4 ^ x5)) : ((~x4 & ~x5) | (~x3 & x4 & x5)))));
  assign n3543 = x2 ? ((~x3 | x4 | ~x7 | x0 | ~x1) & (x1 | (x0 ? (x3 ? (x4 | ~x7) : (~x4 | x7)) : (x7 | (~x3 ^ ~x4))))) : (x3 ? ((x0 | ~x4 | ~x7) & (x1 | ((~x4 | ~x7) & (~x0 | x4 | x7)))) : (x0 ? (~x1 | (x4 ^ x7)) : (x1 | (~x4 ^ x7))));
  assign n3544 = x5 & ((~x4 & n1317 & ~n3546) | (~x3 & ~n3545));
  assign n3545 = (~x2 | ((x4 | ~x6 | x7 | ~x0 | x1) & (x0 | ~x1 | ~x4 | (x6 ^ x7)))) & (~x0 | x1 | x2 | x7 | (~x4 ^ ~x6));
  assign n3546 = (x6 | ~x7 | x1 | ~x2) & (~x1 | x2 | (~x6 ^ ~x7));
  assign n3547 = x0 ? (x2 ? ((x5 | ~x7 | x3 | x4) & (~x3 | ~x4 | (~x5 ^ x7))) : (x3 | (x4 ? (x5 | ~x7) : (x5 ^ x7)))) : ((~x2 | ~x3 | x4 | x5 | ~x7) & ((x5 ^ x7) | (x2 ? (x3 | ~x4) : (~x3 | x4))));
  assign n3548 = ~x5 & ((n1205 & ~n3550) | (~x6 & ~n3549));
  assign n3549 = (x2 | ((x0 | ~x1 | x3 | ~x4 | ~x7) & (~x0 | ~x3 | (x1 ? (x4 | ~x7) : (~x4 | x7))))) & (x0 | ~x1 | ~x2 | ~x7 | (~x3 ^ ~x4));
  assign n3550 = (~x1 | x2 | x3 | x4 | ~x7) & (~x2 | ((x1 | x3 | ~x4 | ~x7) & (~x1 | x7 | (~x3 ^ ~x4))));
  assign z289 = ~n3554 | ~n3558 | (x6 & (n3553 | (~x0 & ~n3552)));
  assign n3552 = (~x2 | ((x1 | x7 | (x3 ? (x4 | ~x5) : (~x4 | x5))) & (~x1 | ~x3 | ~x4 | ~x5 | ~x7))) & (~x1 | x2 | x3 | ((x5 | x7) & (x4 | ~x5 | ~x7)));
  assign n3553 = n651 & ((~x4 & ~x5 & ~x7 & x1 & x3) | (~x1 & x7 & (x3 ? (x4 ^ ~x5) : (x4 & ~x5))));
  assign n3554 = ~n3555 & ~n3557 & (x3 | (n3556 & (~n597 | ~n738)));
  assign n3555 = x5 & (x2 ? ((x3 & ~x4 & ~x0 & x1) | (~x3 & x4 & x0 & ~x1)) : ((x3 & x4 & ~x0 & x1) | (~x4 & (x0 ? (x1 ^ x3) : (~x1 & ~x3)))));
  assign n3556 = (~x4 | ~x5 | ~x6 | ~x0 | ~x1 | x2) & (x0 | x6 | ((~x2 | ~x4 | x5) & (~x1 | (x5 & (~x2 | ~x4)))));
  assign n3557 = ~n1323 & ((~x0 & ~x1 & x5 & (x2 ^ x4)) | (~x5 & (x0 ? (x1 ? (~x2 & ~x4) : (x2 & x4)) : (x1 ? (x2 & x4) : (~x2 & ~x4)))));
  assign n3558 = (~x3 | n3559) & (x6 | (~n1155 & (x1 | n3560)));
  assign n3559 = (x0 | ~x1 | x2 | x4 | ~x5 | x6) & (~x6 | ((x4 | x5 | x0 | x2) & (x1 | (x0 ? (~x2 | (~x4 ^ x5)) : (x5 ? ~x4 : (x2 & x4))))));
  assign n3560 = (~x3 | ((~x0 | x2 | ~x4 | x5 | x7) & (x0 | ~x2 | ~x7 | (~x4 ^ ~x5)))) & (~x0 | x3 | ~x5 | x7 | (x2 & x4));
  assign z290 = n3562 | n3569 | (~n620 & ~n3568);
  assign n3562 = x3 & (n3563 | ~n3565 | (~x1 & ~n3564));
  assign n3563 = ~x1 & (x0 ? (~x4 & x5 & (x2 ^ x6)) : (x4 & ~x5 & (x2 ^ ~x6)));
  assign n3564 = x0 ? (x4 | x5 | (x2 ? (~x6 | ~x7) : (x6 | x7))) : (~x4 | ~x5 | (x2 ? (x6 | x7) : (~x6 | ~x7)));
  assign n3565 = ~n3566 & ~n3567 & (~n757 | ~n750) & (~n924 | ~n1231);
  assign n3566 = ~x0 & ((x1 & ~x2 & x4 & x6 & x7) | (~x1 & ~x4 & (x2 ? (~x6 & ~x7) : (x6 & x7))));
  assign n3567 = (x2 ? (x6 & x7) : (~x6 & ~x7)) & (x0 ? (~x1 & x4) : (x1 & ~x4));
  assign n3568 = x2 ? (((~x3 ^ x5) | (x0 ? (x1 | ~x4) : (~x1 | x4))) & (x0 | ((x1 | (x3 ? (x4 | ~x5) : (~x4 | x5))) & (~x4 | ~x5 | ~x1 | ~x3)))) : ((x3 | (x0 ? (x1 ? (x4 | ~x5) : (~x4 | x5)) : (x1 ? x5 : (x4 | ~x5)))) & (~x4 | x5 | x0 | ~x1) & (~x3 | ((x1 | (x4 ^ x5)) & (~x0 | x4 | x5))));
  assign n3569 = ~x3 & (n3570 | n3571 | n3572 | n3573 | n3575);
  assign n3570 = n1558 & ((x4 & ~x6 & ~x7 & x1 & ~x2) | (~x1 & ~x4 & x7 & (~x2 ^ x6)));
  assign n3571 = x6 & ((~x4 & ~x5 & x0 & ~x1) | (~x0 & x4 & x5 & (~x1 ^ ~x2)));
  assign n3572 = ~n846 & ((~x7 & n664 & ~x2 & ~x4) | (x4 & x7 & n2003));
  assign n3573 = ~n627 & ((n537 & ~n3574) | (x0 & ~x1 & n540));
  assign n3574 = x0 ? (~x1 | x2) : (~x1 ^ ~x2);
  assign n3575 = ~x6 & ((~x0 & ~x1 & x5 & (x2 ^ x4)) | (x1 & (x4 ^ ~x5) & (x0 ^ x2)));
  assign z291 = ~n3581 | ~n3587 | (~x1 & ~n3577) | (~n800 & ~n3580);
  assign n3577 = (~x3 | n3579) & (n3578 | n2744) & (~n1263 | ~n1846);
  assign n3578 = ~x0 ^ ~x6;
  assign n3579 = (~x5 | ~x6 | ~x7 | x0 | ~x2 | ~x4) & (x2 | ((x0 | x4 | x5 | ~x6 | ~x7) & (~x0 | ((x4 | ~x5 | x6 | x7) & (~x6 | ~x7 | ~x4 | x5)))));
  assign n3580 = (x0 | ~x1 | ((~x4 | ~x6 | x2 | ~x3) & (x4 | x6 | ~x2 | x3))) & (x1 | ((x4 | x6 | x2 | x3) & (~x2 | ((x4 | ~x6 | x0 | ~x3) & (~x4 | (x0 ? (x3 ^ x6) : (~x3 | x6)))))));
  assign n3581 = n3583 & ~n3586 & (n620 | n3582) & (~x1 | n3585);
  assign n3582 = (x0 | (x1 ? ((x2 | x3 | x5) & (x4 | ~x5 | ~x2 | ~x3)) : (x4 | (x2 ? (x3 | x5) : (~x3 | ~x5))))) & (x2 | ~x4 | ((~x1 | x3 | x5) & (~x3 | ~x5 | ~x0 | x1)));
  assign n3583 = (n800 | n3584) & (x1 | n806 | (~n2314 & ~n1263));
  assign n3584 = x0 ? (x3 | x4 | (x1 ^ ~x2)) : (~x3 | ~x4 | (~x1 ^ ~x2));
  assign n3585 = (x0 | x2 | x3 | ~x5 | ~x7) & ((x0 & x2) | ((~x5 | ~x7 | x3 | ~x4) & (x5 | x7 | ~x3 | x4)));
  assign n3586 = ~n1429 & (n1574 | (~x4 & n610 & ~n910));
  assign n3587 = ~n3588 & (~x1 | (x0 ? (~n563 | ~n568) : n3589));
  assign n3588 = ~n806 & ((~x1 & ((~x2 & ~x3 & x6) | (x0 & x2 & x3 & ~x6))) | (~x0 & x1 & (x2 ? (~x3 & x6) : (x3 & ~x6))));
  assign n3589 = x3 ? (x5 | ((x4 | ~x6 | ~x7) & (~x2 | ~x4 | x6 | x7))) : (~x5 | x6 | x7 | (x2 & ~x4));
  assign z292 = ~n3596 | (x1 ? ~n3591 : (~n3594 | (~x4 & ~n3593)));
  assign n3591 = x0 ? (~n563 | ~n698) : n3592;
  assign n3592 = x7 ? ((x4 | ~x5 | x2 | x3) & ((x2 ^ ~x3) | (x4 ? (~x5 | x6) : (x5 | ~x6)))) : ((~x5 | x6 | ~x2 | x4) & (x2 | x5 | ~x6 | (~x3 ^ ~x4)));
  assign n3593 = x6 ? ((x0 | x5 | (x2 ? (~x3 | x7) : (x3 | ~x7))) & (~x5 | ((~x0 | (x2 ? (~x3 | ~x7) : (x3 | x7))) & (x0 | x2 | ~x3 | x7)))) : ((x0 | ~x2 | x3 | x5 | x7) & (~x0 | x2 | ~x3 | ~x5 | ~x7));
  assign n3594 = (~x4 | n3595) & (n1007 | (x0 ? (~x2 | (~x4 ^ x7)) : (x2 | (~x4 ^ ~x7))));
  assign n3595 = (~x0 | x2 | x3 | ~x5 | x6 | x7) & (x0 | ((x2 | x3 | x5 | x6 | ~x7) & (~x2 | ~x3 | (x5 ? (x6 | x7) : (~x6 | ~x7)))));
  assign n3596 = n3599 & (x5 ? n3598 : n3597);
  assign n3597 = x1 ? ((x2 | (x3 ? (x4 | x6) : (~x4 | ~x6))) & (x0 | ~x2 | x3 | x4 | x6)) : ((~x4 | x6 | x0 | ~x2) & (~x6 | ((~x0 | ~x2 | ~x3 | ~x4) & (x0 | x4 | (~x2 ^ x3)))));
  assign n3598 = (x1 | (x0 ? (x2 ? (x4 | x6) : (~x4 | ~x6)) : (~x4 | (x2 ? (~x3 | ~x6) : (x3 | x6))))) & (x0 | ~x1 | ~x2 | ((x4 | ~x6) & (~x3 | ~x4 | x6)));
  assign n3599 = x6 ? (x7 ? n3601 : n3600) : (x7 ? n3600 : n3601);
  assign n3600 = x2 ? ((~x4 | x5 | x0 | ~x1) & (x1 | (x0 ? (x3 ? (~x4 | ~x5) : (x4 | x5)) : (x4 | ~x5)))) : ((~x4 | ~x5 | ~x1 | x3) & (~x0 | x1 | x5 | (~x3 ^ x4)));
  assign n3601 = x0 ? ((~x1 | x2 | x3 | x4 | ~x5) & (x1 | x5 | (x2 ? (x3 | ~x4) : (~x3 ^ ~x4)))) : ((x1 | ~x2 | x3 | ~x4 | ~x5) & (~x3 | ((x1 | x2 | ~x4 | ~x5) & (~x1 | x4 | (~x2 ^ x5)))));
  assign z293 = n3603 | ~n3607 | (~n912 & ~n3605) | (~x7 & ~n3606);
  assign n3603 = ~x1 & ((n686 & n1263) | (x4 & ~n3604));
  assign n3604 = (x0 | ~x2 | ~x3 | ~x5 | ~x6 | x7) & (x6 | ~x7 | ((x3 | ~x5 | x0 | ~x2) & (~x0 | x5 | (~x2 ^ ~x3))));
  assign n3605 = (x7 | (x0 ? ((x1 | ~x2 | ~x3) & (~x1 | x2 | x3 | x4)) : (x1 | x2 | (~x3 & ~x4)))) & (x0 | ~x7 | (x1 ? (x2 ? (x3 | x4) : ~x3) : (~x2 | ~x3)));
  assign n3606 = (x3 | ~x4 | x5 | x0 | x1 | ~x2) & (~x1 | ((~x3 | ~x4 | ~x5 | x0 | ~x2) & (~x0 | x2 | x5 | (~x3 ^ x4))));
  assign n3607 = ~n3609 & n3610 & n3612 & (n846 | n3608);
  assign n3608 = ((x3 & x4) | ((x0 | (x1 ? (~x2 | x7) : (x2 | ~x7))) & (~x0 | x1 | ~x2 | ~x7))) & (x4 | ((x0 | ~x1 | x3 | x7) & (x1 | x2 | ((x3 | ~x7) & (~x0 | ~x3 | x7)))));
  assign n3609 = ~n1568 & ((x3 & x4 & x5 & x0 & ~x1) | (~x0 & ~x3 & (x1 ? (x4 & ~x5) : (~x4 & x5))));
  assign n3610 = ~n3611 & (~n723 | ~n814 | ~n677);
  assign n3611 = (~x1 ^ x7) & ((x3 & ~x5 & ~x0 & x2) | (~x3 & x5 & x0 & ~x2));
  assign n3612 = n3613 & (~n664 | ~n2825 | (~n753 & ~n1144));
  assign n3613 = x0 ? (x1 | ((~x5 | x7 | ~x2 | x3) & (x2 | ~x3 | x5 | ~x7))) : (~x1 | x2 | (x3 ? (x5 | x7) : (~x5 | ~x7)));
  assign z294 = n3615 | ~n3616 | ~n3618 | n3623 | (~n662 & ~n3622);
  assign n3615 = n3391 & (x2 ? (~x5 & ~n1403) : (~x3 & n1153));
  assign n3616 = (~x2 | x4 | ~x6 | n3068) & (x2 | ((~x4 | x6 | n3068) & (~x1 | n3617)));
  assign n3617 = (x4 | x5 | x6 | ~x0 | ~x3) & (x0 | ~x6 | (x3 ? (~x4 | ~x5) : (x4 | x5)));
  assign n3618 = ~n3620 & (n620 | n3619) & (x1 | n3621);
  assign n3619 = x1 ? ((x3 | x4 | ~x0 | x2) & (x0 | ~x2 | (x3 ? (x4 | x5) : ~x4))) : (~x3 | (x0 ? (x2 ? (~x4 | ~x5) : x4) : (x2 | ~x4)));
  assign n3620 = x4 & ((~x2 & ~x3 & x6 & ~x0 & ~x1) | (~x6 & ((x0 & x1 & ~x2 & ~x3) | (~x0 & x2 & (~x1 ^ x3)))));
  assign n3621 = (x3 | x6 | ((~x0 | (x2 ? (x4 | x5) : (~x4 | ~x5))) & (x4 | ~x5 | x0 | ~x2))) & (x0 | ~x3 | ~x6 | (x2 ? (~x4 | ~x5) : (x4 | x5)));
  assign n3622 = (x0 | ~x3 | (x4 & x5) | (x1 ^ ~x2)) & (x1 | x3 | ((x2 | (x5 ? x4 : ~x0)) & (~x0 | (x5 ? ~x2 : ~x4))));
  assign n3623 = ~x0 & (x4 ? (n605 & ~n3624) : ~n3625);
  assign n3624 = (x2 | x5 | x6 | x7) & (~x2 | ~x5 | ~x6 | ~x7);
  assign n3625 = (~x5 | ((x1 | x2 | ~x3 | ~x6 | x7) & (~x1 | ((x2 | x3 | ~x6 | x7) & (x6 | ~x7 | ~x2 | ~x3))))) & (x1 | x3 | x5 | ~x7 | (~x2 ^ x6));
  assign z295 = n3627 | n3632 | ~n3635 | (x5 ? ~n3634 : ~n3631);
  assign n3627 = ~x0 & (x1 ? (n3628 & ~n3629) : (~n3630 | (n549 & ~n3629)));
  assign n3628 = x2 & ~x7;
  assign n3629 = (~x3 | x4 | ~x5 | ~x6) & (x3 | ~x4 | x5 | x6);
  assign n3630 = (x7 | ((x2 | ~x3 | x4 | ~x5 | x6) & (x3 | ((x5 | ~x6 | x2 | ~x4) & (~x2 | (x4 ? (~x5 | x6) : (x5 | ~x6))))))) & (~x2 | ~x7 | ((x3 | (x4 ? (~x5 | ~x6) : (x5 | x6))) & (x5 | x6 | ~x3 | ~x4)));
  assign n3631 = x3 ? (x2 ? ((x4 | ~x7 | x0 | ~x1) & (~x4 | x7 | ~x0 | x1)) : ((~x4 | ~x7 | x0 | ~x1) & (x4 | (x0 ? (x1 ^ ~x7) : (x1 | x7))))) : ((~x0 | ~x1 | x2 | x4 | ~x7) & (x1 | ~x2 | (x0 ? (x4 ^ x7) : (~x4 | x7))));
  assign n3632 = x0 & ((~x1 & ~n3633) | (n1082 & n1231));
  assign n3633 = (x4 | ((~x2 | x3 | x5 | ~x6 | ~x7) & (x2 | x6 | (x3 ? (~x5 | ~x7) : (x5 | x7))))) & (~x2 | ~x4 | ~x7 | (x3 ? (x5 | ~x6) : (~x5 | x6)));
  assign n3634 = (x0 | ~x1 | x2 | ~x3 | ~x4 | x7) & (x1 | ((x3 | ~x4 | x7 | x0 | x2) & (~x2 | (~x3 ^ ~x4) | (x0 ^ x7))));
  assign n3635 = x1 ? ((~x4 | x7 | x2 | x3) & (x0 | ((~x2 | ~x4 | (~x3 ^ x7)) & (x4 | ((x3 | x7) & (x2 | ~x3 | ~x7)))))) : ((~x3 | (~x2 ^ x4) | (x0 ^ ~x7)) & (x2 | x3 | ~x7 | (~x0 & x4)));
  assign z296 = ~n3641 | (x2 ? (x3 ? ~n3639 : ~n3640) : ~n3637);
  assign n3637 = (x1 | n3638) & (x3 | ~n568 | ~x0 | ~x1);
  assign n3638 = (x3 | x4 | x5 | x6 | ~x7) & (~x0 | ~x5 | ((x6 | x7 | ~x3 | ~x4) & (x3 | (x4 ? (x6 | ~x7) : (~x6 | x7)))));
  assign n3639 = (x1 | ((x4 | ~x5 | x6 | x7) & (~x6 | ~x7 | ~x4 | x5))) & (x0 | ~x1 | ((~x6 | x7 | ~x4 | x5) & (x4 | ~x5 | x6 | ~x7)));
  assign n3640 = (~x0 | x1 | x4 | x5 | ~x6 | ~x7) & (x0 | ~x1 | ((~x4 | (x5 ? (~x6 | x7) : (x6 | ~x7))) & (~x6 | x7 | x4 | x5)));
  assign n3641 = ~n3643 & ~n3645 & (x3 ? n3646 : (n3642 & n3644));
  assign n3642 = ((x4 ^ x6) | ((x0 | ~x1 | ~x2 | x5) & (~x0 | x1 | x2 | ~x5))) & (x1 | x2 | x4 | x5 | ~x6) & (x0 | ((~x4 | ((~x5 | ~x6 | x1 | ~x2) & (~x1 | x6 | (x2 ^ x5)))) & (x1 | x5 | ~x6 | (x2 & x4))));
  assign n3643 = n1317 & ((~x1 & ~x2 & ~x4 & x5 & x6) | (x1 & ((~x2 & ~x4 & x5 & ~x6) | (x2 & (x4 ? (~x5 & ~x6) : (x5 & x6))))));
  assign n3644 = (~x0 | ~x1 | x2 | ~x4 | x5) & (x1 | ~x5 | ((~x2 | x4) & (x0 | x2 | ~x4)));
  assign n3645 = ~n1429 & ((x1 & ~x2 & ~x3 & ~x4) | (x0 & ~x1 & (x2 ? (~x3 & x4) : (x3 & ~x4))));
  assign n3646 = (x1 | x2 | ~x4 | x5) & ((~x4 ^ ~x5) | ((x0 | ~x1 | x2) & (x1 | ~x2)));
  assign z297 = ~n3648 | ~n3652;
  assign n3648 = (~n1416 | n3651) & (~x1 | n3650) & (n846 | n3649);
  assign n3649 = (~x0 & (x3 ? (x4 & x7) : ~x2)) | (~x2 & ((~x1 & ~x3 & x4) | (x0 & ~x4 & ~x7))) | (x3 & ((x0 & x1) | (x2 & x4))) | (x2 & ((x0 & (x1 | (x4 & ~x7))) | (~x3 & ~x4) | (x1 & x4 & ~x7)));
  assign n3650 = (x2 | x3 | x4 | x5 | ~x6) & (x0 | ((~x5 | x6 | ~x3 | ~x4) & (x3 | ((~x2 | x4 | ~x5 | x6) & (~x4 | x5 | ~x6)))));
  assign n3651 = (x2 | ~x3 | x4 | x5 | ~x6) & (x3 | ((x2 | ~x4 | ~x5 | x6) & (x1 | ((~x5 | ~x6 | x2 | x4) & (~x2 | (x4 ? (x5 | ~x6) : (~x5 | x6)))))));
  assign n3652 = (x1 | n3653) & (~x7 | (x0 ? n3655 : n3654));
  assign n3653 = x4 ? (x3 ? (~x5 | x6 | (x0 & ~x2)) : (x5 | (x0 ? (x2 ^ x6) : (x2 | ~x6)))) : (x0 ? ((x2 | x5 | ~x6) & (~x2 | x3 | ~x5 | x6)) : (x3 | (x2 ? (x5 | ~x6) : (~x5 | x6))));
  assign n3654 = (~x2 | ~x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (~x1 | ((~x2 | x3 | x4 | x5 | ~x6) & (x2 | ((x5 | x6 | x3 | x4) & (~x5 | ~x6 | ~x3 | ~x4)))));
  assign n3655 = (~x4 | ((x2 | x3 | ~x5 | x6) & (x1 | ((x2 | ~x5 | x6) & (x5 | ~x6 | ~x2 | ~x3))))) & (x1 | ~x2 | x4 | (x3 ? (~x5 | x6) : (x5 | ~x6)));
  assign z298 = ~n3658 | n3662 | n3663 | (~n800 & ~n3657);
  assign n3657 = (x3 | (x4 ? ((x0 | ((x2 | ~x6) & (~x1 | ~x2 | x6))) & (~x1 | x2 | ~x6) & (~x0 | x1 | ~x2 | x6)) : ((x2 | x6) & (x0 | ~x2 | ~x6)))) & ((~x2 ^ ~x6) | (x0 ? (x1 | x4) : (~x3 | ~x4)));
  assign n3658 = ~n3660 & n3661 & (n3659 | (n1215 & n846));
  assign n3659 = (~x2 | ~x3 | ~x4 | ~x0 | x1) & (x0 | ((x2 | ~x3 | x4) & (x3 | ~x4 | x1 | ~x2)));
  assign n3660 = ~n3458 & (x0 ? (~x1 & ~x4) : ((~x3 & ~x4) | (~x1 & x3 & x4)));
  assign n3661 = (~n1102 | n3341) & (~n565 | ~n720);
  assign n3662 = ~n630 & (x2 ? (~x4 & ((~x1 & x3) | (~x0 & (~x1 | x3)))) : ((~x3 & (x4 ? x1 : x0)) | (x4 & (~x0 | (~x1 & x3)))));
  assign n3663 = x4 & ((n1343 & n540 & n750) | (~x3 & ~n3664));
  assign n3664 = (~x1 | ((x6 | x7 | x2 | x5) & (~x5 | ~x6 | ~x7 | x0 | ~x2))) & (~x0 | ((x6 | x7 | x2 | x5) & (x1 | ~x5 | ~x6 | (~x2 ^ ~x7))));
  assign z299 = n3666 | n3670 | ~n3671 | (~x3 & ~n3669);
  assign n3666 = ~x0 & (x7 ? ~n3668 : ~n3667);
  assign n3667 = (x3 | ((x4 | ~x5 | x6) & (~x1 | ((~x4 | x5 | ~x6) & (x2 | ~x5 | x6))))) & (x1 | ~x3 | ((~x5 | x6 | ~x2 | ~x4) & (x4 | (x5 ^ x6))));
  assign n3668 = ((x5 ^ x6) | ((x1 | ~x3 | ~x4) & (~x1 | ~x2 | x3 | x4))) & (x1 | ~x3 | x4 | x5 | ~x6) & (~x4 | ((~x5 | ~x6 | ~x2 | ~x3) & (x1 | x3 | (x2 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n3669 = x4 ? ((x0 | (x1 ? (~x5 | ~x7) : (x5 | x7))) & (~x5 | ~x7 | ((~x1 | x2) & (~x0 | x1 | ~x2)))) : ((~x5 | (x0 ? (x7 | (x1 ^ ~x2)) : (~x7 | (x1 & x2)))) & (~x0 | x5 | ~x7 | (x1 ^ ~x2)));
  assign n3670 = ~n1862 & ((x3 & ~x5 & ~x0 & x1) | (x5 & ~n910 & x0 & ~x3));
  assign n3671 = (n620 | n3674) & (~n738 | n3672) & (~x3 | n3673);
  assign n3672 = ((~x5 ^ x7) | ((x2 | x3 | x4 | x6) & (~x3 | ~x4 | ~x6))) & (~x3 | ((x4 | (x5 ? (x6 | ~x7) : (~x6 | x7))) & (x6 | x7 | ~x4 | x5))) & (x3 | ((x5 | x6 | x7 | ~x2 | x4) & (x2 | ~x6 | ((~x5 | ~x7) & (~x4 | x5 | x7)))));
  assign n3673 = (~x4 | x5 | ~x7 | x0 | ~x1) & (x7 | ((x0 | ~x1 | (~x4 ^ ~x5)) & (x2 | ((x0 | ~x4 | ~x5) & (~x1 | x4 | x5)))));
  assign n3674 = (~x3 | x4 | ~x5 | x0 | ~x1) & (x3 | ((x0 | x1 | ~x2 | ~x4 | ~x5) & (x5 | (x0 ? (~x4 | (x1 ^ ~x2)) : (x4 | (x1 & x2))))));
  assign z300 = n3676 | ~n3681 | (x1 ? ~n3679 : ~n3680);
  assign n3676 = ~x0 & ((x5 & ~n3677) | (n1120 & ~n3678));
  assign n3677 = (~x2 | ((x6 | x7 | x1 | ~x4) & (~x3 | ((x6 | ~x7 | x1 | x4) & (~x1 | ~x6 | (x4 ^ x7)))))) & (~x1 | x2 | ((x6 | x7 | ~x3 | x4) & (x3 | ~x7 | (x4 & x6))));
  assign n3678 = (x3 | x4 | x7 | ~x1 | x2) & (x1 | (~x2 & ~x3) | (~x4 ^ ~x7));
  assign n3679 = (x2 | ((x4 | ~x5 | ~x6 | x0 | ~x3) & (~x0 | x5 | ((x4 | x6) & (x3 | ~x4 | ~x6))))) & (x0 | ~x5 | ((~x3 | ~x4 | x6) & (~x2 | ((x3 | x4 | ~x6) & (~x4 | x6)))));
  assign n3680 = (~x4 | ((~x5 | ~x6 | x0 | ~x2) & (x5 | (x0 ? ((~x2 & ~x3) | ~x6) : x6)))) & (x2 | x4 | ((x5 | ~x6 | x0 | x3) & (~x0 | ~x3 | ~x5 | x6)));
  assign n3681 = (n662 | n3684) & (n620 | n3683) & (~n738 | n3682);
  assign n3682 = (x5 | x6 | ((~x2 | ((x4 | ~x7) & (x3 | ~x4 | x7))) & (~x3 | ((x4 | ~x7) & (x2 | ~x4 | x7))))) & (x2 | ~x5 | ((~x3 | x4 | ~x6 | ~x7) & (x3 | x7 | (~x4 & ~x6))));
  assign n3683 = (~x4 | ((~x1 | ((x0 | x5) & (x3 | ~x5 | ~x0 | x2))) & (~x0 | x1 | ((x2 | x3 | x5) & (~x5 | (~x2 & ~x3)))))) & (x0 | x1 | x4 | ~x5 | (x2 & x3));
  assign n3684 = (x0 | x1 | x2 | ~x4 | ~x5) & (x4 | ((~x1 | ((x3 | ~x5 | ~x0 | x2) & (x0 | x5 | (~x2 & ~x3)))) & (~x0 | x1 | (x2 ? ~x5 : (x3 | x5)))));
  assign z301 = ~n3687 | (~x1 & ((~x2 & ~n3686) | (n943 & n1263)));
  assign n3686 = (x5 | ~x6 | x7 | x0 | x3 | x4) & (~x4 | x6 | ((~x5 | ~x7 | x0 | x3) & (~x0 | (x3 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n3687 = ~n3688 & ~n3689 & ~n3690 & n3691 & (n918 | n1009);
  assign n3688 = ~x0 & ((x1 & ~x2 & x3 & ~x5 & x7) | (x2 & ((~x5 & ~x7 & ~x1 & ~x3) | (x1 & ((x5 & ~x7) | (~x3 & ~x5 & x7))))));
  assign n3689 = x4 & n539 & ((n723 & n610) | (~x0 & ~n1875));
  assign n3690 = x0 & ((x1 & ~x2 & ~x3 & ~x5 & ~x7) | (x3 & x5 & x7 & ~x1 & x2));
  assign n3691 = (~x5 | (x6 ? n3694 : n3692)) & (x1 | n3693) & (x5 | (x6 ? n3692 : n3694));
  assign n3692 = (x0 | ~x1 | x2 | x3 | x4 | ~x7) & (x1 | (x0 ? (x7 | (x3 ? (x2 & x4) : ~x2)) : (~x7 | (~x2 & ~x3))));
  assign n3693 = (x0 | x2 | ~x4 | x5 | x7) & (~x0 | ~x5 | ((x4 | ~x7 | ~x2 | x3) & (x2 | (x3 ? (~x4 | ~x7) : (x4 | x7)))));
  assign n3694 = (x2 | (x3 & x4) | (x0 ? (x1 | ~x7) : (~x1 | x7))) & (x0 | ~x2 | ~x3 | (x1 ^ x7));
  assign z302 = ~n3700 | (~n662 & ~n3699) | (~x2 & (~n3696 | ~n3698));
  assign n3696 = x0 ? (~n605 | ~n568) : n3697;
  assign n3697 = (~x5 | ~x6 | ~x7 | x1 | x3 | ~x4) & (x4 | ((x1 | x3 | x5 | x6 | ~x7) & (~x1 | ~x5 | (x3 ? (x6 | ~x7) : (~x6 | x7)))));
  assign n3698 = (x6 | ((x0 | x1 | x3 | (~x4 & ~x5)) & (~x1 | (x0 ? x3 : (~x3 | ~x4))))) & (~x0 | x1 | ~x6 | (~x3 ^ (x4 & x5)));
  assign n3699 = (x0 | ~x1 | ~x2 | ~x3) & (x1 | ((x0 | x2 | ~x3) & (x3 | (x4 & x5) | (~x0 ^ x2))));
  assign n3700 = (~x2 | n3704) & (n3701 | n3702) & (n620 | n3703);
  assign n3701 = (~x1 | x2 | x4 | x5) & (x1 | ~x2 | ~x4 | ~x5);
  assign n3702 = x0 ? (~x3 | x6) : (x3 | ~x6);
  assign n3703 = (~x0 | x1 | ~x2 | (x3 & x4)) & (x2 | ((~x3 | ~x4 | ~x5 | ~x0 | x1) & (x0 | ~x1 | (x3 ? (x4 | x5) : ~x4))));
  assign n3704 = (~x4 | x5 | x6 | ~x0 | x1 | ~x3) & (x0 | (x1 ? (x3 | x6) : (~x3 | ~x6)));
  assign z303 = ~n3708 | ~n3710 | (~x2 & (~n3706 | ~n3707));
  assign n3706 = (x4 | ((x0 | ((x1 | x3 | ~x5 | x7) & (x5 | ~x7 | ~x1 | ~x3))) & (~x0 | ~x1 | ~x3 | x5 | x7))) & (~x0 | x1 | ~x4 | (x3 ? (x5 ^ x7) : (x5 | ~x7)));
  assign n3707 = ((~x3 ^ x7) | (x0 ? (x1 | x4) : (~x1 | ~x4))) & (x0 | x3 | x7 | (~x1 ^ x4));
  assign n3708 = (x3 | ((x0 | ~x1 | ~x2 | x7) & (~x0 | (x1 ? (x2 | x7) : (~x2 | ~x7))))) & n3709 & (x0 | ~x3 | (x1 ? (~x2 | ~x7) : (~x2 ^ x7)));
  assign n3709 = (~n943 | ~n1476) & (~n2205 | ~n923 | ~n1546);
  assign n3710 = (x0 | n3711) & (~n538 | ((x4 | ~x7 | x0 | x3) & (~x0 | ~x3 | (~x4 ^ x7))));
  assign n3711 = (n1545 | n3712) & (~n563 | ~n2237 | n3713);
  assign n3712 = (~x1 | ~x3 | x4 | x7) & (x1 | x3 | ~x4 | ~x7);
  assign n3713 = x1 ? (~x5 | ~x7) : (x5 | x7);
  assign z304 = x7 ? ~n3715 : ~n3717;
  assign n3715 = n531 & (~n750 | ~n1478) & (x3 | n3716);
  assign n3716 = (x0 | ~x1 | ~x2 | x4 | x5 | x6) & ((x0 ^ ~x6) | ((~x1 | x2 | x4 | ~x5) & (x1 | ~x4 | (~x2 ^ x5))));
  assign n3717 = ~n3718 & ~n3720 & (x6 ? (n785 | ~n2010) : n3719);
  assign n3718 = ~x0 & ((x1 & ((x3 & x4) | (~x4 & ~x5 & x2 & ~x3))) | (x3 & (x2 ? (~x4 & x5) : (x4 & ~x5))) | (~x1 & ((x3 & ~x4) | (x4 & x5 & x2 & ~x3))));
  assign n3719 = x0 ? (x3 | ((~x4 | x5 | x1 | ~x2) & (~x1 | x2 | x4 | ~x5))) : (x1 | ~x3 | ~x4 | (~x2 ^ x5));
  assign n3720 = x0 & ((x1 & ~x2 & ~x3 & ~x4 & ~x5) | (~x1 & ((x3 & x4 & x5) | (x2 & (x3 ^ ~x4)))));
  assign z305 = ~n3728 | (x6 ? ~n3725 : (n3723 | (~x2 & ~n3722)));
  assign n3722 = (x0 | x1 | x3 | x4 | x5 | ~x7) & (~x5 | (x0 ? (x7 | (x1 ? (x3 | ~x4) : (~x3 | x4))) : (~x3 | ~x7 | (~x1 ^ x4))));
  assign n3723 = ~x5 & n871 & ((n738 & n1835) | (~x0 & n3724));
  assign n3724 = x7 & (~x1 ^ ~x4);
  assign n3725 = (~n3726 | ~n677) & (~x2 | n3727);
  assign n3726 = x7 & x5 & ~x3 & x4;
  assign n3727 = (x0 | x1 | x3 | ~x4 | x5 | ~x7) & ((x3 ? (~x4 | ~x5) : (x4 | x5)) | (x0 ? (x1 | x7) : (~x1 | ~x7)));
  assign n3728 = ~n3729 & n3730 & ~n3731 & n3733 & (~n3336 | n3732);
  assign n3729 = ~n785 & ((~x0 & x1 & ~n571) | (~x1 & ~n783 & ~n2189));
  assign n3730 = (x2 | x4 | x5 | ~x0 | x1) & (x0 | ((~x1 | (x2 ? (x4 | ~x5) : (~x4 | x5))) & (x1 | ~x2 | ~x4 | ~x5)));
  assign n3731 = ~x1 & (((x3 ^ x5) & (x0 ? (x2 & x4) : (~x2 & ~x4))) | (~x0 & x2 & ~x3 & ~x4 & ~x5) | (x3 & x4 & x5 & x0 & ~x2));
  assign n3732 = (~x1 | x2 | x3 | x4 | ~x6) & (x1 | ~x2 | ~x3 | ~x4 | x6);
  assign n3733 = (~n677 | ~n921) & (x3 | ~n2095 | ~n694);
  assign z306 = (~x0 & ~n3735) | (x0 & ~n3739) | (x2 & ~n3743) | (~x2 & ~n3742);
  assign n3735 = (~x2 | n3738) & (n1323 | n3737) & (x2 | x4 | n3736);
  assign n3736 = x1 ? ((x3 | x5 | ~x6 | x7) & (x6 | ~x7 | ~x3 | ~x5)) : ((~x3 | x5 | ~x6 | x7) & (x3 | x6 | (~x5 ^ x7)));
  assign n3737 = x5 ? ((~x2 | x4 | x7) & (x1 | x2 | ~x4 | ~x7)) : ((x1 | ~x2 | ~x4 | ~x7) & (~x1 | (x2 ? (x4 | ~x7) : (~x4 | x7))));
  assign n3738 = (x1 | x3 | x4 | x5 | x6 | x7) & (~x5 | ~x6 | ~x7 | ~x1 | ~x3 | ~x4);
  assign n3739 = (n824 | n3740) & (x1 | n3741);
  assign n3740 = (~x1 | x2 | x3 | ~x4 | x6) & (x1 | ~x3 | (x2 ? (~x4 | ~x6) : (x4 | x6)));
  assign n3741 = (~x6 | ((x4 | x5 | ~x7 | ~x2 | x3) & (x2 | x7 | (x3 ? (~x4 | ~x5) : (x4 | x5))))) & (~x2 | x6 | ((x5 | ~x7 | ~x3 | x4) & (~x5 | x7 | x3 | ~x4)));
  assign n3742 = (((~x5 | ~x6) & (x4 | x5 | x6)) | (~x0 ^ x3)) & (x4 | ((~x5 | ~x6 | x1 | ~x3) & (~x1 | x3 | x5 | x6))) & (x0 | x1 | x3 | x5 | ~x6) & (~x4 | (x5 ? ((~x0 | x1 | ~x3 | x6) & (~x1 | (x3 ? x0 : ~x6))) : (x6 | ((x1 | x3) & (x0 | (x1 & x3))))));
  assign n3743 = (x5 | ((~x4 | (x0 ? (x1 | (~x3 ^ x6)) : (~x1 | (~x3 & ~x6)))) & (~x3 | ~x6 | (x0 & (x1 | x4))))) & (x3 | ~x5 | x6 | (x0 & (x1 | x4)));
  assign z307 = ~n3752 | (x2 ? ~n3747 : (x3 ? ~n3746 : ~n3745));
  assign n3745 = x7 ? (x0 ? ((~x1 | ~x4 | x6) & (x1 | x4 | x5 | ~x6)) : (x1 ? (x5 | ~x6) : (x4 ? (~x5 | ~x6) : x6))) : ((x4 | ((x5 | ~x6 | x0 | x1) & (~x0 | (x1 ? (~x5 | ~x6) : (x5 | x6))))) & (~x0 | ~x4 | x5 | ~x6) & (x0 | x6 | ((~x4 | ~x5) & (~x1 | (~x4 & ~x5)))));
  assign n3746 = x4 ? ((x1 | ((~x6 | ~x7 | ~x0 | ~x5) & (x0 | ((~x6 | x7) & (~x5 | x6 | ~x7))))) & (x0 | x5 | ((~x6 | x7) & (~x1 | x6 | ~x7)))) : ((x0 | x1 | x5 | (x6 ^ x7)) & ((~x6 ^ x7) | (x0 ? x1 : (~x1 | ~x5))));
  assign n3747 = ~n3749 & ~n3750 & (x1 ? (x0 | ~n3751) : n3748);
  assign n3748 = (x5 | ((x0 | x3 | x4 | x6 | ~x7) & (~x0 | ((~x6 | x7 | x3 | ~x4) & (~x3 | x4 | x6 | ~x7))))) & (x0 | x3 | ~x5 | (x4 ? (x6 | x7) : (~x6 | ~x7)));
  assign n3749 = ~n620 & ((~x1 & x4 & (x0 ? (~x3 & x5) : (x3 & ~x5))) | (~x0 & x3 & ~x4 & (x1 | x5)));
  assign n3750 = ~n662 & ((~x0 & x1 & x5 & (x3 ^ ~x4)) | (~x1 & ((x4 & ~x5 & ~x0 & ~x3) | (x0 & (x3 ? x4 : (~x4 & ~x5))))));
  assign n3751 = ~x3 & ~x5 & (x4 ? (~x6 & ~x7) : (x6 & x7));
  assign n3752 = (x1 | n3755) & (n1323 | n3754) & (x0 | ~x1 | n3753);
  assign n3753 = (x2 | ~x3 | x4 | x5 | ~x6) & (x3 | ((x4 | x5 | x6) & (~x2 | ~x4 | ~x5 | ~x6)));
  assign n3754 = x0 ? ((~x1 | x2 | x4 | x5) & (x1 | ~x5 | (~x2 ^ x4))) : (~x4 | (x1 ? (~x2 ^ x5) : (~x2 | ~x5)));
  assign n3755 = (x2 | (x0 ? ((~x5 | ~x6 | x3 | x4) & (x5 | x6 | ~x3 | ~x4)) : ((x3 | ~x4 | x5 | x6) & (~x5 | ~x6 | ~x3 | x4)))) & (x0 | ~x2 | x4 | (x3 ? (x5 | ~x6) : (~x5 | x6)));
  assign z308 = ~n3762 | (x2 ? (n3760 | (~x1 & ~n3761)) : ~n3757);
  assign n3757 = (~x5 | (n3758 & (~x0 | n662 | n1688))) & ~n3759 & (x0 | x5 | n662 | n1688);
  assign n3758 = (x1 | ((x4 | ~x6 | x7 | x0 | x3) & (~x0 | ((x3 | ~x4 | ~x6 | x7) & (x6 | ~x7 | ~x3 | x4))))) & (x0 | x3 | ((x4 | x6 | ~x7) & (~x1 | ((x6 | ~x7) & (~x4 | ~x6 | x7)))));
  assign n3759 = ~n3172 & (x1 ? n2205 : n1156);
  assign n3760 = ~n592 & ((x3 & ~x5 & ~x6 & x0 & ~x1) | (~x0 & ((~x1 & ~x3 & x5 & x6) | (x1 & (x3 ? (x5 & ~x6) : (~x5 & x6))))));
  assign n3761 = ((~x0 ^ ~x3) | ((~x6 | x7 | x4 | x5) & (x6 | ~x7 | ~x4 | ~x5))) & (x5 | ~x6 | ~x7 | ~x0 | x3 | ~x4) & (x0 | ~x3 | x4 | ~x5 | x6 | x7);
  assign n3762 = (~x1 | n3765) & (x1 | n3763) & (n927 | n3764);
  assign n3763 = (~x2 | (((x4 ? (x5 | ~x7) : (~x5 | x7)) | (x0 ^ x3)) & (x0 | ~x3 | ~x5 | (~x4 ^ x7)))) & (~x0 | x3 | x5 | (~x4 ^ x7)) & (x2 | ((~x0 | x5 | (~x4 ^ x7)) & (x3 | (x4 ? ((x5 | x7) & (x0 | ~x5 | ~x7)) : ((x5 | ~x7) & (~x0 | ~x5 | x7))))));
  assign n3764 = x0 ? (x3 | (x1 ? (x2 | x5) : (~x2 | ~x5))) : (~x3 | (x1 ? (x2 | x5) : (~x2 ^ x5)));
  assign n3765 = (~x0 | x2 | ~x3 | x4 | x5 | x7) & (x0 | (((~x4 ^ x7) | (x2 ? (~x3 ^ x5) : (~x3 | ~x5))) & (~x2 | ((x5 | x7 | x3 | x4) & (~x5 | ~x7 | ~x3 | ~x4))) & (x2 | x3 | ~x4 | x5 | ~x7)));
  assign z309 = ~n3772 | (x1 ? ~n3769 : (x3 ? ~n3768 : ~n3767));
  assign n3767 = x0 ? ((x6 | x7 | x4 | x5) & (~x4 | ((x5 | ~x6 | ~x7) & (x6 | x7 | x2 | ~x5)))) : ((~x2 | ~x6 | (x4 ? (x5 | x7) : (~x5 | ~x7))) & (x5 | x6 | ((x4 | ~x7) & (x2 | ~x4 | x7))));
  assign n3768 = (~x7 | ((x4 | ((~x5 | ~x6 | ~x0 | x2) & (x0 | (x2 ? (~x5 | x6) : (x5 | ~x6))))) & (~x0 | ~x2 | ~x4 | (~x5 ^ ~x6)))) & (~x5 | x7 | ((~x2 | (x0 ? (x4 | x6) : (~x4 | ~x6))) & (x0 | x2 | (~x4 ^ x6))));
  assign n3769 = (n824 | n3771) & (~x0 | ~n563 | ~n686) & (x0 | n3770);
  assign n3770 = (~x7 | ((~x2 | x3 | x4 | x5 | ~x6) & (x6 | ((x4 | ~x5 | x2 | ~x3) & (~x2 | ~x4 | (x3 ^ x5)))))) & (~x4 | x7 | ((~x5 | x6 | ~x2 | x3) & (x2 | ~x6 | (x3 ^ x5))));
  assign n3771 = (~x0 | x2 | x3 | ~x4 | x6) & (x0 | ~x2 | ~x3 | x4 | ~x6);
  assign n3772 = (x0 | n3775) & (n846 | n3774) & (~x0 | n3773);
  assign n3773 = (~x4 | ~x5 | ~x6 | ~x1 | x2 | x3) & (x1 | ((~x2 | (x3 ? (x5 | ~x6) : (~x5 | x6))) & (x4 | ((x3 | ~x5) & (x2 | ~x3 | x5)))));
  assign n3774 = (x2 | (x0 ? (x1 ? (x3 | x4) : (~x3 | ~x4)) : (~x1 | (~x3 ^ x4)))) & (x0 | ~x2 | (x1 ? (~x3 | ~x4) : (~x3 ^ x4)));
  assign n3775 = x1 ? (x5 ? (x6 | ((x3 | x4) & (x2 | ~x3 | ~x4))) : ((~x2 | (x3 ? (x4 | x6) : (~x4 | ~x6))) & (x2 | x3 | x4 | ~x6))) : (x2 ? ((x5 | ~x6 | x3 | x4) & (~x5 | x6 | ~x3 | ~x4)) : (x3 ? (x4 ? (x5 | ~x6) : (~x5 | x6)) : (~x5 | (~x4 & ~x6))));
  assign z310 = ~n3777 | ~n3782 | (~n620 & ~n3781);
  assign n3777 = (n1568 | n3780) & (~n1123 | n3778) & (n662 | n3779);
  assign n3778 = (x1 | ~x2 | x5 | (x3 ? (~x6 | x7) : (x6 | ~x7))) & (x2 | ((x5 | ~x6 | ~x7 | x1 | ~x3) & (~x1 | x3 | x7 | (~x5 ^ ~x6))));
  assign n3779 = x3 ? (~x5 | ((x1 | x2 | x4) & (x0 | (x1 ? (~x2 ^ x4) : (~x2 | ~x4))))) : (x5 | ((~x0 | (x1 ? (x2 | x4) : ~x4)) & (x1 | ~x2 | ~x4) & (x0 | ~x1 | (~x2 ^ x4))));
  assign n3780 = (x0 | ~x1 | ((x3 | ~x4 | ~x5 | x6) & (x5 | ~x6 | ~x3 | x4))) & (x1 | ((x0 | x3 | x4 | ~x5 | ~x6) & (~x0 | ~x3 | ~x4 | (x5 ^ x6))));
  assign n3781 = x3 ? (~x5 | ((x1 | ~x2 | x4) & (x0 | (x1 ? (x2 ^ x4) : (x2 | ~x4))))) : (x5 | (x0 ? (x1 ? (x2 | ~x4) : x4) : (~x4 | (~x1 ^ ~x2))));
  assign n3782 = ~n3784 & ~n3786 & (x1 | n3783) & (n2286 | n3785);
  assign n3783 = ((x3 ? (x4 | x5) : (~x4 | ~x5)) | ((x2 | x6) & (~x0 | ~x2 | ~x6))) & (~x2 | x3 | x4 | ~x5 | x6) & (x2 | x5 | ~x6 | ((~x3 | ~x4) & (x0 | x3 | x4)));
  assign n3784 = ~n1007 & ((x0 & x1 & ~x2 & ~x4) | (~x0 & (x1 ? (x2 ^ x4) : (x2 & x4))));
  assign n3785 = (~x5 | x6 | ~x0 | x1) & (x5 | ~x6 | x0 | ~x1);
  assign n3786 = n1701 & n610 & ((~n1116 & n873) | (n543 & n539));
  assign z311 = ~n3794 | (x0 & ~n3793) | (~x3 & ~n3788) | (x3 & ~n3792);
  assign n3788 = (n910 | n3790) & (x1 | n3789) & (x0 | ~x1 | n3791);
  assign n3789 = (~x5 | x6 | ~x7 | ~x0 | x2 | ~x4) & (x4 | ((x6 | ~x7 | x2 | x5) & (x0 | ~x6 | ((~x5 | ~x7) & (x2 | x5 | x7)))));
  assign n3790 = (x5 | x6 | x7 | ~x0 | ~x4) & ((x0 ? (~x4 | ~x5) : (x4 | x5)) | (~x6 ^ x7));
  assign n3791 = (~x2 | x4 | x5 | x6 | ~x7) & (~x6 | x7 | ~x4 | ~x5);
  assign n3792 = (x1 | ((~x0 | ~x4 | ~x5 | x6 | x7) & ((x5 ^ x7) | (x0 ? (~x4 | ~x6) : (x4 | x6))))) & (x0 | ((~x1 | ~x4 | ~x5 | x6 | x7) & (~x6 | ~x7 | x4 | x5)));
  assign n3793 = (~x1 | x2 | ~x3 | x4 | x5 | x7) & (x3 | ((x1 | ~x2 | x4 | x5 | ~x7) & (~x1 | x2 | ((x5 | ~x7) & (x4 | ~x5 | x7)))));
  assign n3794 = (~x4 & ((~x5 & x7) | (~x0 & ~x1 & (~x5 | x7)))) | (x1 & (x0 | (x4 & x5 & ~x7))) | (~x3 & (~x5 ^ x7)) | (x3 & (x5 ^ x7)) | (x0 & x4 & (x5 | ~x7));
  assign z312 = n932 | n3796 | ~n3800 | (~x0 & ~n3799);
  assign n3796 = ~x2 & (x1 ? ~n3798 : ~n3797);
  assign n3797 = x6 ? ((~x0 | x3 | ~x4 | ~x5 | ~x7) & ((~x4 ^ x7) | (x0 ? (x3 | x5) : ~x5))) : ((x3 | x4 | ~x5 | x7) & (~x0 | ~x3 | x5 | (~x4 ^ ~x7)));
  assign n3798 = (x5 | (x0 ? (x6 | ((x4 | x7) & (x3 | ~x4 | ~x7))) : (~x6 | ((~x3 | x4 | ~x7) & (~x4 | x7))))) & (x0 | ~x5 | x6 | ((~x3 | x4 | x7) & (~x4 | ~x7)));
  assign n3799 = x1 ? (~x4 | (x5 ? ~x6 : ((~x2 & ~x3) | x6))) : ((~x4 | ~x5 | x6) & (x2 | x3 | (x4 ? x6 : (x5 | ~x6))));
  assign n3800 = (~n534 | ~n2112) & (~x2 | n3801);
  assign n3801 = (x6 | (~x4 ^ ~x7) | (x0 ? (x1 | x5) : (~x1 | ~x5))) & (x0 | ~x6 | (~x1 ^ x5) | (~x4 ^ x7));
  assign z313 = ~n3806 | (~x2 & (~n3803 | ~n3805));
  assign n3803 = (~n698 | ~n937) & (x3 | n3804);
  assign n3804 = (~x5 | (((x4 ^ x6) | (x0 ? (x1 | ~x7) : (~x1 | x7))) & (x1 | x7 | (x0 ? (x4 | ~x6) : (~x4 | x6))))) & (x0 | ~x1 | x5 | (~x4 ^ (x6 & ~x7)));
  assign n3805 = x5 ? ((~x3 | ((~x6 | x7 | x0 | ~x1) & (x1 | (x6 ? ~x0 : x7)))) & (~x0 | ~x1 | x3 | (~x6 & x7))) : (((x0 ? (x1 | x3) : (~x1 | ~x3)) | (x6 ^ x7)) & (~x0 | x6 | ~x7 | (x1 ^ ~x3)));
  assign n3806 = (~x2 | ((x1 | ((~x5 | (x6 ^ x7)) & (~x0 | (x5 ? x7 : (x6 | ~x7))))) & (x0 | ~x1 | (x5 ? (~x6 | x7) : (x6 ^ x7))))) & (x0 | ((~x5 | x6 | ~x7) & (x1 | (x5 ? ~x7 : (~x6 | x7)))));
  assign z314 = ~n3810 | (~x2 & (n3809 | (~x5 & ~n3808)));
  assign n3808 = (~x6 | ((x0 | x3 | (x1 ? (~x4 | ~x7) : (x4 | x7))) & (~x0 | ~x1 | ~x3 | x4 | x7))) & (~x0 | ~x3 | x4 | x6 | (x1 ^ x7));
  assign n3809 = n1489 & n1163;
  assign n3810 = n946 & (~n947 | ((~x1 | x4 | ~x6 | ~x7) & (x1 | ~x4 | x6 | x7)));
  assign z315 = (~x2 & (~n3812 | (~x7 & ~n1655))) | ~n3813;
  assign n3812 = (x4 | ((x0 | x1 | x3 | x5 | ~x7) & (~x0 | ~x3 | x7 | (~x1 ^ x5)))) & (x0 | ~x1 | x3 | ~x4 | (x5 ^ x7));
  assign n3813 = (~x0 | x2 | x3 | (~x1 ^ x7)) & (x0 | (x1 ? (~x7 | (~x2 & ~x3)) : (~x3 | x7))) & ~n3814 & (x1 | ~x2 | x7);
  assign n3814 = ~n2805 & ~n620 & ~x4 & n670;
  assign z316 = n3816 | ~n3818 | ~n3819 | (n3628 & ~n3817);
  assign n3816 = ~x0 & ~x3 & ((~x4 & ~x5 & ~x1 & x2) | (x1 & x4 & (x2 ^ x5)));
  assign n3817 = (x0 | ~x1 | x3 | ~x4 | ~x5 | x6) & (~x0 | x1 | ~x3 | x4 | x5 | ~x6);
  assign n3818 = (x0 | x2 | ~x3) & (x1 | ((x2 | ~x3 | (~x4 & ~x5)) & (~x0 | ~x2 | x3)));
  assign n3819 = (x1 | x2 | ~x4 | ~n732) & (x4 | (x1 ? (~x2 | ~n732) : (n2805 | (~x2 ^ x6))));
  assign z317 = n2499 | n3822 | ~n3825 | (~x0 & ~n3821);
  assign n3821 = x3 ? (x4 | (x5 & x6) | (~x1 ^ ~x2)) : (~x4 | ~x5 | (x1 ? (~x2 | ~x6) : x2));
  assign n3822 = x2 & (n3823 | (x4 & n664 & n618));
  assign n3823 = x6 & n2512 & ((n2205 & n1317) | (x0 & n3824));
  assign n3824 = ~x5 & (~x3 ^ x7);
  assign n3825 = ~n3826 & ~n3827 & n3828 & (~x3 | ~n1449 | ~n738);
  assign n3826 = x4 & (x0 ? (~x1 & x3) : (~x5 & (x1 ^ ~x3)));
  assign n3827 = ~x0 & ~x4 & x5 & x6 & (x1 ^ ~x3);
  assign n3828 = (~n650 | ~n1120 | ~n534) & (~n720 | ~n686);
  assign z318 = ~n3833 | ~n3831 | ~n2516 | ~n3830;
  assign n3830 = (~n1546 | ~n1179) & (~n757 | ~n1176) & (~n1148 | n1139);
  assign n3831 = ~n3832 & (~n1102 | ((~x4 | x6 | ~x1 | x3) & (x1 | ~x3 | (~x4 ^ x6))));
  assign n3832 = ~x0 & x5 & ((x4 & x6 & x1 & x2) | (~x1 & ((~x2 & ~x4 & x6) | (x4 & ~x6))));
  assign n3833 = ~n3835 & (~x6 | (~n3834 & (~n814 | ~n534 | ~n691)));
  assign n3834 = ~n592 & ((~x0 & ~x1 & x2 & x3 & x5) | (x0 & ~x5 & (x1 ? (~x2 & ~x3) : x2)));
  assign n3835 = n1121 & (x4 ? (x7 & n2758) : (~x7 & (x3 ? n2758 : n534)));
  assign z319 = n3840 | n3842 | (~x3 & ~n3837) | (~x1 & ~n3839);
  assign n3837 = (~x2 | x6 | x7 | n627 | ~n664) & (x2 | n3838);
  assign n3838 = (x0 | ~x1 | (x6 & x7) | (~x4 ^ ~x5)) & (x1 | ((~x5 | ~x6 | ~x0 | x4) & (x0 | ~x4 | x5 | x6 | x7)));
  assign n3839 = (~x7 & ((~x0 & (x2 ? (x3 & x6) : (~x3 & ~x6))) | (~x2 & ((~x3 & x5 & ~x6) | (x0 & x6))) | (x0 & ~x5 & (x2 | x3)))) | (x0 & x7 & (x5 ^ ~x6)) | (~x2 & ~x3 & ~x5 & x6) | (~x0 & (x5 ^ x6));
  assign n3840 = x1 & ~n3841;
  assign n3841 = x0 ? (x2 | x3 | (~x5 ^ (x6 & x7))) : ((~x3 | ((x2 | ~x5) & (x6 | x7 | ~x2 | x5))) & (~x5 | ((~x6 | ~x7) & (~x2 | (~x6 & ~x7)))));
  assign n3842 = n544 & n904 & (x0 ? (~x2 & ~n868) : (x2 & n2095));
  assign z320 = n3844 | ~n3846 | ~n3848 | (~n620 & ~n3845);
  assign n3844 = n1943 & ((x3 & ~x5 & ~x6 & x0 & ~x2) | (~x0 & ~x3 & x5 & (~x2 ^ x6)));
  assign n3845 = x0 ? (x1 | x2 | x3 | (x4 & x5)) : (~x1 | ~x2 | (~x3 & ~x4));
  assign n3846 = (~n534 | ~n1590) & (x1 | ~x6 | n3847);
  assign n3847 = (~x0 | x2 | x3 | ~x4 | ~x5) & (~x3 | x4 | x5 | x0 | ~x2);
  assign n3848 = ~n3850 & (n662 | n3849);
  assign n3849 = x1 ? (x2 | x3 | (~x0 & (x4 | x5))) : ((~x0 | (~x2 & (~x3 | ~x4))) & (~x2 | ~x3 | (~x4 & ~x5)));
  assign n3850 = ~x0 & (x1 ? (~x6 & (~x2 ^ (~x3 & ~x4))) : (x6 & (~x2 | ~x3)));
  assign z321 = n3855 | ~n3857 | (x4 ? ~n3856 : (n3852 | n3854));
  assign n3852 = ~x2 & ~n3853;
  assign n3853 = (x5 | ~x6 | x7 | x0 | x1 | x3) & (~x7 | ((x0 | ~x1 | x3 | ~x5 | x6) & (~x0 | ~x3 | (x1 ? (x5 | x6) : (~x5 | ~x6)))));
  assign n3854 = n616 & ((n2155 & n2747) | (n2503 & n904));
  assign n3855 = n1123 & ((~x3 & ((x5 & ~x7 & ~x1 & ~x2) | (x1 & (x2 ? (x5 ^ ~x7) : (~x5 & x7))))) | (~x1 & x2 & x3 & (x5 ^ ~x7)));
  assign n3856 = (x3 | x7 | x0 | x2) & (~x7 | ((x2 | ~x3 | ~x0 | x1) & (x0 | ~x2 | (~x1 ^ x3))));
  assign n3857 = (~x7 | ((x0 | ~x1 | ~x2 | ~x3) & (~x0 | (x1 ? (x2 | x3) : ~x2)))) & n3858 & (x0 | x7 | ((x2 | ~x3) & (x1 | ~x2 | x3)));
  assign n3858 = ~n3859 & (~n943 | ~n1476) & (~n534 | ~n1979);
  assign n3859 = x0 & ~x1 & ~x2 & ~x4 & (x3 ^ x7);
  assign z322 = n3863 | ~n3864 | (~x4 & (n3862 | (x5 & ~n3861)));
  assign n3861 = x0 ? (x1 | ~x3 | (x2 ? (x6 | ~x7) : (~x6 | x7))) : (~x1 | x3 | (x2 ? (x6 | x7) : (~x6 | ~x7)));
  assign n3862 = n1120 & ((n651 & ~n1150) | (x2 & n598 & n2527));
  assign n3863 = n650 & ((~x2 & ~x5 & ~x6 & x0 & x1) | (~x1 & ((x0 & x5 & (~x2 ^ x6)) | (~x5 & ~x6 & ~x0 & x2))));
  assign n3864 = (x4 | x5 | ((x2 | ~x3 | ~x0 | x1) & (x0 | ~x2 | x3))) & (x1 | ~x2 | (x0 ? (~x3 | ~x4) : x3)) & (x2 | ((~x1 | x3 | ~x4) & ((~x1 & ~x4 & ~x5) | (~x0 ^ x3))));
  assign z323 = n3866 | n3869 | n3870 | ~n3871 | (~x4 & ~n3868);
  assign n3866 = ~x1 & ((~x4 & ~n3867) | (n1415 & n1163));
  assign n3867 = x0 ? (x7 | ((~x5 | x6 | ~x2 | ~x3) & (x2 | ~x6 | (~x3 ^ ~x5)))) : ((x2 | x3 | ~x5 | x6 | ~x7) & (~x2 | ~x3 | x5 | ~x6 | x7));
  assign n3868 = x1 ? (x2 | ((x0 | x3 | (~x5 ^ x6)) & (~x3 | (x0 ? (x5 | x6) : (~x5 | ~x6))))) : (x0 ? ((~x5 | ~x6 | ~x2 | x3) & (x2 | x6 | (~x3 ^ ~x5))) : ((~x5 | ~x6 | x2 | x3) & (x5 | x6 | ~x2 | ~x3)));
  assign n3869 = ~x4 & ((~x0 & ((~x1 & ~x2 & x3 & ~x5) | (x2 & (x1 ? (~x3 ^ x5) : (~x3 & x5))))) | (~x2 & ~x3 & x5 & x0 & x1));
  assign n3870 = n1943 & ((x0 & ~x2 & x3 & ~x5 & x6) | (~x0 & ~x3 & x5 & (x2 ^ x6)));
  assign n3871 = n3872 & (~x4 | ((x0 | (x1 ^ x3)) & (x3 | ((x1 | ~x2) & (~x0 | ~x1 | x2)))));
  assign n3872 = (~x5 | ~x6 | ~n534 | x3 | ~x4) & (x5 | ~n738 | ~x3 | x4);
  assign z324 = n3874 | n3876 | n3880 | ~n3881 | (~x2 & ~n3879);
  assign n3874 = ~x5 & ((n650 & n544 & n694) | (~x1 & ~n3875));
  assign n3875 = (x4 | ~x6 | x7 | x0 | ~x2 | ~x3) & (x3 | ((~x4 | ~x6 | ~x7 | x0 | ~x2) & (x2 | ((x6 | ~x7 | x0 | x4) & (~x0 | ~x6 | (x4 ^ x7))))));
  assign n3876 = x5 & ((~x6 & ~n3878) | (n738 & n2825 & ~n3877));
  assign n3877 = (~x4 | ~x7) & (~x3 | x4 | x7);
  assign n3878 = x0 ? (x1 | ((~x4 | x7 | x2 | x3) & (~x2 | ~x3 | (x4 ^ x7)))) : (x1 ? ((~x4 | ~x7 | x2 | ~x3) & (x4 | x7 | ~x2 | x3)) : (x2 | x3 | (x4 ^ x7)));
  assign n3879 = x0 ? (x4 | x6 | (x1 ? (~x3 | x5) : (x3 ^ x5))) : ((x3 | x4 | x5 | (x1 ^ ~x6)) & (~x5 | ((x3 | ~x4 | ~x6) & (~x1 | ((~x4 | ~x6) & (~x3 | x4 | x6))))));
  assign n3880 = (~x4 ^ x5) & ((x1 & (x0 ? (~x2 & ~x3) : x2)) | (~x0 & ((x2 & ~x3) | (~x1 & ~x2 & x3))));
  assign n3881 = n3882 & (~n538 | ((n783 | n1936) & (~n669 | ~n957)));
  assign n3882 = (x0 | ~x1 | x2 | ~x3 | x4 | x5) & (x1 | ((~x3 | ~x4 | ~x5 | x0 | ~x2) & (~x0 | x4 | x5 | (~x2 & ~x3))));
  assign z325 = n3884 | n3888 | ~n3890 | (~n1099 & ~n3887);
  assign n3884 = ~x2 & (x0 ? ~n3885 : ~n3886);
  assign n3885 = (~x4 | ((~x5 | x7 | x1 | ~x3) & (~x1 | x3 | x5 | ~x6 | ~x7))) & (x3 | x4 | x5 | x6 | ~x7) & (x1 | ((~x6 | x7 | x3 | x5) & (~x3 | ((~x5 | x6 | x7) & (~x6 | ~x7 | x4 | x5)))));
  assign n3886 = (x1 | x3 | ~x5 | x6 | x7) & (x5 | ((x3 | x4 | x6 | ~x7) & (~x1 | ~x3 | ~x4 | (~x6 ^ x7))));
  assign n3887 = (x0 | ((~x1 | ((x5 | ~x6) & (x2 | ~x5 | x6))) & (~x6 | ((x2 | x5) & (~x5 | ~x7 | x1 | ~x2))) & (x5 | ((~x2 | x6 | ~x7) & (x1 | (x7 ? x6 : ~x2)))))) & (x2 | ((~x0 | x1 | ~x5 | (~x6 ^ x7)) & (~x1 | x5 | (x6 ? x7 : ~x0)))) & (~x0 | x1 | ~x2 | (x5 ? (x6 | x7) : ~x6));
  assign n3888 = x2 & (n3889 | (~x4 & ~x5 & n738 & ~n2181));
  assign n3889 = ~n906 & ((x0 & ~x1 & x4 & x5 & ~x6) | (~x0 & ~x4 & (x1 ? (~x5 & ~x6) : (x5 & x6))));
  assign n3890 = ~n3893 & ~n3894 & (n3891 | n3494) & (x5 | n3892);
  assign n3891 = (x3 | x4 | x6 | x7) & (~x3 | ~x4 | ~x6 | ~x7);
  assign n3892 = (~x6 | (x0 ? ((x1 | ~x2 | ~x3 | ~x4) & (~x1 | x2 | x3 | x4)) : (~x3 | ~x4 | (~x1 ^ ~x2)))) & (x1 | x3 | x6 | (x0 ? (x2 | ~x4) : (~x2 | x4)));
  assign n3893 = ~n1687 & ((~x5 & ((~x1 & x2 & x7) | (~x0 & (~x1 | x2)))) | (~x2 & x5 & (x0 ? (~x1 & x7) : (x1 & ~x7))));
  assign n3894 = x5 & n538 & (n3895 | (n642 & n610));
  assign n3895 = x6 & x4 & ~x0 & x3;
  assign z326 = ~n3902 | (x2 ? ~n3899 : (x0 ? ~n3897 : ~n3898));
  assign n3897 = (x1 | (~x6 ^ x7)) & (x4 | x5 | x7 | ((~x3 | ~x6) & (~x1 | x3 | x6)));
  assign n3898 = (~x3 | ((x1 | x4 | x5 | x6 | x7) & (~x1 | ~x4 | (x6 ^ x7)))) & (x1 | x3 | (x6 ? ~x7 : (x7 | (~x4 & ~x5))));
  assign n3899 = x0 ? (x1 | ~n3900) : n3901;
  assign n3900 = x3 & (x6 ^ ~x7);
  assign n3901 = x7 ? (x1 ? ((~x5 | x6 | ~x3 | ~x4) & (x3 | x4 | ~x6)) : (x6 | (x4 ? x3 : (~x3 & ~x5)))) : ((~x6 | ((~x3 | (x1 ? (~x4 | ~x5) : (x4 | x5))) & (x1 | x3 | (~x4 & ~x5)))) & (~x1 | x3 | x6 | (x4 & x5)));
  assign n3902 = ~n3903 & ~n3904 & ~n3905 & (~n1120 | ~n616 | n739);
  assign n3903 = ~x0 & ((x1 & ~x2 & x3 & ~x4 & ~x6) | (x2 & ((~x1 & x3 & x4 & ~x6) | (x1 & x6 & (x3 ^ x4)))));
  assign n3904 = ~x3 & ((x0 & (x1 ? (~x2 & x6) : (x2 & ~x6))) | (~x0 & x1 & ~x2 & ~x6));
  assign n3905 = x6 & x3 & ~x2 & ~x0 & ~x1;
  assign z327 = n3907 | ~n3910 | (~x0 & ~n3909);
  assign n3907 = ~x1 & ((n2317 & n686) | (x3 & ~n3908));
  assign n3908 = (x0 | x2 | x4 | x5 | (x6 ^ x7)) & (~x5 | ((x0 | ~x2 | x4 | x6 | x7) & (~x4 | ~x6 | ~x7 | ~x0 | x2)));
  assign n3909 = (~x2 | ((~x1 | ~x3 | ~x4 | x5 | ~x7) & ((~x3 ^ x7) | (x1 ? (~x4 | ~x5) : (x4 | x5))))) & (x1 | x4 | ~x5 | (~x3 ^ ~x7));
  assign n3910 = ~n3911 & ~n3912 & (~n694 | ~n2692) & (~n1977 | n3913);
  assign n3911 = x0 & ((~x2 & ((~x1 & ~x7) | (x4 & x7 & x1 & ~x3))) | (~x1 & ((x3 & ~x7) | (x2 & ~x3 & x7))));
  assign n3912 = ~x0 & ((x4 & ((x3 & ~x7 & x1 & ~x2) | (~x1 & (~x3 ^ x7)))) | (x1 & (x3 ? (~x4 & x7) : (x2 ? (~x4 & ~x7) : x7))));
  assign n3913 = (~x0 | x2 | ~x3 | x4 | x6 | ~x7) & (x3 | (x6 ^ x7) | (x0 ? (x2 | x4) : (~x2 | ~x4)));
  assign z328 = ~n3921 | n3918 | n3916 | n3369 | n3915 | n3368;
  assign n3915 = ~x0 & ~x1 & ((x2 & ~x4 & ~x5) | (x4 & x5 & (~x2 | ~x3)));
  assign n3916 = x2 & ((n1880 & n1846) | (x7 & ~n3917));
  assign n3917 = x0 ? (x1 | ((~x5 | ~x6 | x3 | x4) & (x5 | x6 | ~x3 | ~x4))) : (~x1 | x4 | x5 | (~x3 ^ ~x6));
  assign n3918 = ~x2 & ((n605 & n2238 & ~n3920) | (x6 & ~n3919));
  assign n3919 = x0 ? ((x1 | ~x3 | ~x4 | ~x5 | x7) & (~x1 | x5 | (x3 ? (x4 | x7) : (~x4 | ~x7)))) : ((~x1 | x3 | x4 | ~x5 | x7) & (~x4 | x5 | ~x7 | x1 | ~x3));
  assign n3920 = x0 ? (~x5 | x7) : (x5 | ~x7);
  assign n3921 = n3922 & (~n1184 | (x0 ? (~x1 | ~n2984) : (x1 | (~n2984 & ~n2985))));
  assign n3922 = (~x1 | ((x3 | ~x4 | ~x5 | ~x0 | x2) & (x0 | ((~x2 | ((x4 | ~x5) & (~x3 | ~x4 | x5))) & (x4 | (x5 ? ~x3 : x2)))))) & (~x0 | x1 | ((x2 | ((~x4 | x5) & (x3 | x4 | ~x5))) & (~x4 | (x5 ? ~x2 : x3))));
  assign z329 = ~n3929 | (x0 ? ~n3924 : (x3 ? ~n3927 : ~n3928));
  assign n3924 = x4 ? n3925 : n3926;
  assign n3925 = ((x5 ^ x7) | ((x1 | ~x2 | ~x3 | x6) & (~x1 | x2 | x3 | ~x6))) & (x1 | x2 | ((~x6 | x7 | ~x3 | ~x5) & (x3 | x6 | (~x5 ^ x7))));
  assign n3926 = (~x3 | ((x1 | x6 | ~x7 | (x2 ^ x5)) & (x5 | ~x6 | x7 | ~x1 | x2))) & (x1 | ~x2 | x3 | ~x6 | (~x5 ^ x7));
  assign n3927 = x6 ? ((x5 ^ x7) | (x1 ? (~x2 | x4) : (x2 | ~x4))) : ((x1 | ~x2 | x4 | (~x5 ^ x7)) & (~x1 | x2 | ~x4 | ~x5 | ~x7));
  assign n3928 = (x5 | x6 | x7 | ~x1 | ~x2 | x4) & (x2 | (x1 ? (~x6 | (x4 ? (x5 | ~x7) : (~x5 | x7))) : (x6 | (x4 ? (x5 | x7) : (~x5 | ~x7)))));
  assign n3929 = ~n3376 & ~n3930 & ~n3931 & ~n3933 & (x0 | n3932);
  assign n3930 = ~n1099 & (x6 ? ~n3378 : (n539 & ~n2111));
  assign n3931 = n738 & ((~x2 & ~x3 & ~x4 & ~x5) | (x5 & ((~x2 & x3 & ~x4 & ~x6) | (x2 & (x3 ? (x4 & x6) : ~x6)))));
  assign n3932 = x2 ? ((x4 | ~x5 | ~x6 | ~x1 | x3) & (x5 | (x1 ? (~x3 | (~x4 & x6)) : (x3 | (x4 & x6))))) : ((~x1 | ~x3 | ~x4 | ~x5 | ~x6) & (x1 | ((x3 | ~x5 | ~x6) & (x5 | x6 | ~x3 | ~x4))));
  assign n3933 = ~n912 & ((x0 & ~x1 & ~x2 & n814) | (~x0 & (x1 ? (~x2 & n690) : (x2 & n814))));
  assign z330 = n3935 | ~n3937 | (~n662 & ~n3945) | (~x0 & ~n3944);
  assign n3935 = ~x3 & ((n587 & n1546) | (~x2 & ~n3936));
  assign n3936 = (~x0 | ((x1 | x4 | ~x5 | ~x6 | ~x7) & (~x1 | ~x4 | x5 | x6 | x7))) & (~x5 | ~x6 | ~x7 | x0 | ~x1 | ~x4);
  assign n3937 = ~n3939 & ~n3940 & ~n3941 & n3942 & (n620 | n3938);
  assign n3938 = (x4 | ((~x0 | ((x1 | ~x2 | x3) & (~x3 | x5 | ~x1 | x2))) & (~x2 | ((x0 | ~x1 | ~x3) & (x1 | x3 | x5))))) & (~x2 | ~x3 | x5 | x0 | ~x1) & (x2 | ((x0 | (x1 ? (x3 | ~x5) : (~x3 | ~x4))) & (~x4 | (x1 ? x3 : (~x3 | ~x5)))));
  assign n3939 = n738 & ((x4 & ~x5 & ~x6 & ~x2 & x3) | (~x4 & ((~x5 & x6 & x2 & x3) | (~x2 & (x3 ? (x5 & ~x6) : (~x5 & x6))))));
  assign n3940 = ~x0 & x3 & ((x1 & ~x2 & ~x4 & x6) | (~x1 & ~x6 & (~x2 ^ x4)));
  assign n3941 = ~x3 & ((x0 & ((x4 & x6 & ~x1 & x2) | (x1 & ~x2 & ~x4 & ~x6))) | (~x0 & x1 & x2 & x4 & ~x6));
  assign n3942 = (~n559 | ~n2609) & (~n3943 | n739) & (~n568 | ~n1229);
  assign n3943 = x7 & x6 & ~x0 & ~x5;
  assign n3944 = (~x4 | ~x5 | ~x6 | ~x1 | ~x2 | ~x3) & (x3 | ((x4 | ((~x1 | x6 | (x2 ^ x5)) & (~x5 | ~x6 | x1 | ~x2))) & (x1 | ~x4 | (x2 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n3945 = (x0 | ~x1 | ((~x4 | ~x5 | x2 | ~x3) & (x4 | x5 | ~x2 | x3))) & (x1 | (x4 ? ((x2 | x3 | x5) & (~x0 | (x2 ? (~x3 | x5) : x3))) : ((~x2 | ~x3 | ~x5) & (x0 | (x2 ? ~x3 : (x3 | ~x5))))));
  assign z331 = n3947 | n3949 | (x2 ? ~n3953 : ~n3952);
  assign n3947 = x0 & ((~x1 & ~n3948) | (n1082 & n762));
  assign n3948 = x2 ? (~x3 | ((x6 | ~x7 | x4 | x5) & (~x4 | ~x5 | (x6 ^ x7)))) : ((~x3 | ~x4 | ~x5 | ~x6 | x7) & (x4 | (x3 ? (x5 | (x6 ^ x7)) : (~x5 | (~x6 ^ x7)))));
  assign n3949 = ~x0 & ((n708 & ~n3951) | (~x5 & ~n3950));
  assign n3950 = (~x6 | (x2 ^ x7) | (x1 ? (~x3 | ~x4) : (x3 | x4))) & (x2 | x6 | ~x7 | ((x3 | x4) & (~x1 | ~x3 | ~x4)));
  assign n3951 = x1 ? ((x2 | ~x4 | ~x6 | ~x7) & (~x2 | x4 | x6 | x7)) : (~x4 | x7 | (x2 ^ x6));
  assign n3952 = x4 ? ((~x0 | ((x3 | ~x5 | x7) & (x5 | ~x7 | x1 | ~x3))) & (x0 | ((x7 | (x3 ^ x5)) & (x1 | ((x5 | x7) & (x3 | ~x5 | ~x7))))) & (x3 | x7 | (x1 ^ x5))) : ((x0 | (x3 ? ~x7 : (~x5 | x7))) & (~x5 | ~x7 | x1 | ~x3) & (~x0 | ((x3 | x5 | ~x7) & (~x1 | (x3 ? (x5 | x7) : ~x7)))));
  assign n3953 = (x1 & (x0 | (x3 & ~x5 & x7))) | (x4 & ((~x7 & (~x3 | x5)) | (~x0 & ~x1 & (~x7 | (~x3 & x5))))) | (~x4 & ((x7 & (x3 | ~x5)) | (x0 & (x7 | (x3 & ~x5))))) | (x0 & x3 & x7) | (x5 & ~x7 & ~x0 & ~x3);
  assign z332 = n3956 | n3957 | ~n3960 | (~x1 & ~n3955);
  assign n3955 = (x2 | ((~x4 | x5 | x0 | ~x3) & (~x5 | ~x6 | ~x0 | x4))) & (~x2 | ((x4 | ~x5 | (x0 ^ x3)) & (~x0 | x3 | x5 | (~x4 & x6)))) & (x0 | ((~x5 | ~x6 | x3 | ~x4) & (~x3 | x5 | x6))) & (~x0 | ((~x3 | ~x5 | ~x6) & (x3 | ~x4 | x5 | x6)));
  assign n3956 = ~n912 & ((~x0 & x2 & x3 & (x1 ^ x4)) | (~x2 & (x0 ? (x1 ? (~x3 & x4) : (x3 & ~x4)) : (x1 ? (x3 & x4) : (~x3 & ~x4)))));
  assign n3957 = x3 & ((x7 & ~n3958 & x0 & ~x1) | (~x0 & (x1 ? ~n3959 : (~x7 & ~n3958))));
  assign n3958 = (~x5 | x6 | x2 | ~x4) & (x5 | ~x6 | ~x2 | x4);
  assign n3959 = (~x5 | x6 | x7 | x2 | x4) & (~x2 | ~x4 | x5 | ~x6 | ~x7);
  assign n3960 = (~x1 | n3961) & (x3 | (x2 ? n3963 : n3962));
  assign n3961 = (~x0 | x2 | x3 | x4 | x5 | x6) & (x0 | (x4 ? (x3 ? (~x5 | (~x2 & ~x6)) : (x5 | x6)) : ((~x3 | x5 | x6) & (x3 | ~x5 | ~x6) & (x2 | (~x3 ^ x5)))));
  assign n3962 = ((x4 ? (x6 | ~x7) : (~x6 | x7)) | (x0 ? (~x1 | x5) : (x1 | ~x5))) & (~x6 | ((~x0 | x1 | ~x4 | x5 | x7) & (x0 | ~x1 | ~x7 | (~x4 ^ ~x5))));
  assign n3963 = (~x5 | x6 | x7 | ~x0 | x1 | ~x4) & (x0 | (x1 ? ((~x6 | x7 | ~x4 | x5) & (x4 | ~x5 | x6 | ~x7)) : (~x7 | (x4 ? (~x5 | x6) : (x5 | ~x6)))));
  assign z333 = n3965 | ~n3969 | (~n592 & ~n3967) | (~x0 & ~n3968);
  assign n3965 = ~x2 & ((~x3 & ~n3966) | (n559 & n937));
  assign n3966 = (x0 | ~x1 | x4 | x5 | ~x6 | ~x7) & (~x4 | ((~x1 | ((x6 | ~x7 | ~x0 | x5) & (x0 | ~x5 | (x6 ^ x7)))) & (~x0 | x1 | x7 | (~x5 ^ ~x6))));
  assign n3967 = (~x3 | ((x0 | ~x1 | x2 | ~x5 | x6) & (x5 | ~x6 | x1 | ~x2))) & (x0 | x1 | ~x2 | x5 | ~x6) & (x3 | ((~x0 | ~x1 | x2 | x5 | ~x6) & (x0 | ~x5 | (x1 ? (~x2 | x6) : (x2 | ~x6)))));
  assign n3968 = x1 ? ((x2 | x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (x5 | x6 | ~x2 | x4) & (~x5 | ((~x3 | x4 | ~x6) & (~x2 | ((x4 | ~x6) & (~x3 | ~x4 | x6)))))) : ((~x4 | x5 | x6) & (~x6 | ((~x2 | x3 | ~x4 | ~x5) & (x2 | ((x4 | x5) & (~x3 | ~x4 | ~x5))))));
  assign n3969 = ~n3971 & ~n3972 & (~n762 | ~n1620) & (n927 | n3970);
  assign n3970 = (x0 | ((~x5 | x6 | x1 | x3) & (x5 | ~x6 | ~x1 | ~x2))) & (x1 | ((~x5 | x6 | ~x2 | x3) & (x2 | ((~x3 | ~x5 | x6) & (x5 | ~x6 | ~x0 | x3)))));
  assign n3971 = ~n783 & ((~x1 & x2 & x3 & x5) | (x1 & ~x2 & (x0 ? (~x3 & x5) : (x3 & ~x5))));
  assign n3972 = n738 & (((x4 ^ ~x5) & (x2 ? (~x3 & x6) : (~x3 ^ x6))) | (~x2 & ~x3 & ~x4 & x5 & x6) | (x4 & ~x5 & ~x6 & (x2 | x3)));
  assign z334 = n3974 | ~n3979 | (x7 ? ~n3978 : ~n3977);
  assign n3974 = ~x5 & (x0 ? ~n3975 : ~n3976);
  assign n3975 = (x1 | ~x2 | ((~x6 | x7 | x3 | x4) & (x6 | ~x7 | ~x3 | ~x4))) & (x2 | x4 | x6 | ((x3 | x7) & (~x1 | ~x3 | ~x7)));
  assign n3976 = (x3 | x4 | ~x7 | ~x1 | x2) & (~x4 | ((x1 | x2 | x3 | x6 | x7) & (~x1 | ((x2 | x3 | ~x6 | x7) & (x6 | ~x7 | ~x2 | ~x3)))));
  assign n3977 = (x1 | (x2 ? (x5 ^ x6) : (x3 | (x0 ? (~x5 | x6) : (x5 | ~x6))))) & (x0 | ((~x2 | (x5 ^ x6)) & (x5 | x6 | ~x1 | x3)));
  assign n3978 = (~x1 & ((x5 & x6) | (~x0 & x2 & x3))) | (x2 & (x6 ? x5 : x3)) | (~x2 & ~x3 & (~x5 | ~x6)) | (~x5 & ~x6) | (x3 & x5 & x6) | (x0 & x1);
  assign n3979 = ~n3980 & (~n1132 | n3981) & (~x3 | ~n1156 | ~n1546);
  assign n3980 = ~x2 & (x3 ? (~x5 & ~x7 & (~x0 | ~x1)) : ((x5 & x7 & ~x0 & ~x1) | (x0 & ((~x5 & x7) | (x1 & x5 & ~x7)))));
  assign n3981 = x0 ? (x1 | (x4 ? ~x7 : (~x6 | x7))) : (~x1 | (x4 ? (x6 | ~x7) : x7));
  assign z335 = n3983 | ~n3986 | (~n857 & ~n3989) | (~x3 & ~n3990);
  assign n3983 = ~x6 & (n3985 | (~x4 & ~n3984));
  assign n3984 = (x7 | (x0 ? ((x1 | ~x2 | ~x3 | ~x5) & (~x1 | x2 | x3 | x5)) : (~x2 | ~x3 | (x1 ^ x5)))) & (x1 | ~x7 | ((x2 | ~x3 | ~x5) & (x0 | (x2 ? (x3 | x5) : ~x3))));
  assign n3985 = x3 & x4 & ((~x0 & x1 & x2 & ~x7) | (~x1 & ((~x2 & x7) | (x0 & x2 & ~x7))));
  assign n3986 = (n1387 | n3988) & (~n686 | ~n754) & (n1568 | n3987);
  assign n3987 = (x0 | ((~x3 | ~x6) & (~x1 | x3 | x4 | x5 | x6))) & (x1 | ((~x3 | ~x6) & (x4 | x5 | x6 | ~x0 | x3)));
  assign n3988 = (~x0 | x3 | x4 | x5 | ~x6) & (x0 | ~x3 | x6 | (~x4 & ~x5));
  assign n3989 = x2 ? (x6 | (x3 ^ (~x4 & ~x5))) : (x3 | ~x6);
  assign n3990 = (x2 | ~x6 | x0 | x1) & ((~x4 & ~x5) | ((x0 | x1 | ~x2 | x6) & (x2 | ~x6 | ~x0 | ~x1)));
  assign z336 = ~n3994 | (n597 & ~n3992) | (~x4 & ~n3993);
  assign n3992 = x3 ? ((x0 | ((~x6 | x7) & (~x1 | x6 | ~x7))) & (x6 | ~x7 | (x1 ? x2 : ~x0))) : (x0 ? ((x2 | ~x6 | ~x7) & (x1 | ((~x6 | ~x7) & (x2 | x6 | x7)))) : ((~x2 | x6 | x7) & (~x1 | ((x6 | x7) & (~x2 | ~x6 | ~x7)))));
  assign n3993 = (~x5 | (x3 ? (x7 | (x0 & x1)) : (~x7 | (~x0 ^ (x1 & x2))))) & (~x0 | x3 | x5 | x7 | (x1 ^ ~x2));
  assign n3994 = (x1 & ((x2 & ~x4) | (x0 & (x2 | ~x7)))) | (x3 & x7) | (~x3 & ~x7) | (~x4 & (x0 | ~x7));
  assign z337 = n3997 | ~n3998 | (~x2 & (n3996 | (n1543 & n1838)));
  assign n3996 = ~x5 & ((~n945 & ~n3172) | (n3098 & n1229));
  assign n3997 = x4 & ((x2 & ((~x5 & x6 & ~x0 & x1) | (x0 & ~x1 & x5))) | (~x0 & ~x1 & ~x2 & (x5 | x6)));
  assign n3998 = ~n4000 & (n910 | n3999) & (~n1156 | ~n648 | n3578);
  assign n3999 = (x0 | ~x4 | (~x5 & ~x6)) & (x4 | x5 | ((x6 | x7) & (~x0 | (x6 & x7))));
  assign n4000 = (x0 ? (~x1 & ~x2) : (x1 & x2)) & (x4 ? x5 : (~x5 & ~x6));
  assign z338 = n4002 | n4005 | ~n4006 | (n563 & ~n4004);
  assign n4002 = ~x2 & ((n650 & n1543 & n653) | (~x3 & ~n4003));
  assign n4003 = (~x0 | x1 | x4 | ~x5 | ~x6 | x7) & (x0 | x6 | ((x1 | ~x4 | x5 | x7) & (~x1 | ~x7 | (~x4 ^ x5))));
  assign n4004 = (x0 | x6 | (x1 ? (x5 | x7) : (~x5 | ~x7))) & (~x5 | ~x6 | ~x7 | ~x0 | x1);
  assign n4005 = ~n824 & ((x0 & x1 & ~x2 & ~x3 & x6) | (~x1 & (x2 | x3) & (~x0 ^ x6)));
  assign n4006 = (x0 | ~x5 | ~x6) & (x5 | x6 | (x0 ^ (~x1 | (~x2 & ~x3))));
  assign z341 = ~x2 & (n4008 | ~n4009);
  assign n4008 = ~x1 & (x3 ? ((x0 & (~x5 | ~x6)) | (~x4 & (x0 | (~x5 & ~x6)))) : ((x4 & (~x0 | (x5 & x6))) | (~x0 & (x5 | x6))));
  assign n4009 = (x1 | n550 | n4010) & (x0 | ~x1 | (n1099 & n4011));
  assign n4010 = x3 ? (~x6 | x7) : (x6 | ~x7);
  assign n4011 = (x5 | x6 | x7 | ~x3 | ~x4) & (x3 | x4 | ~x5 | ~x6 | ~x7);
  assign z342 = ~n4016 | (x3 & (n4014 | (n1843 & ~n4013)));
  assign n4013 = (~x6 | x7 | ~x2 | x4) & (x6 | ~x7 | x2 | ~x4);
  assign n4014 = ~x1 & (x0 ? n4015 : (n2503 & n1148));
  assign n4015 = x4 & ((~x6 & ~x7 & x2 & ~x5) | (x6 & x7 & ~x2 & x5));
  assign n4016 = ~n4017 & ~n4018 & n4019 & (~n664 | ~n1343 | n2587);
  assign n4017 = ~x0 & ((x1 & ~x2 & x3 & x4 & x5) | (~x1 & ((x4 & ~x5 & x2 & ~x3) | (~x2 & x3 & ~x4 & x5))));
  assign n4018 = x2 & ((~x0 & x1 & ~x3) | (~x1 & ((~x3 & ~x4) | (x0 & (~x3 | ~x4)))));
  assign n4019 = ~n598 | (~n4020 & (~n1812 | ~n568));
  assign n4020 = x4 & ~x2 & x3;
  assign z343 = n4022 | ~n4027 | (x0 ? ~n4026 : ~n4025);
  assign n4022 = x7 & ((n664 & ~n4024) | (~x1 & ~n4023));
  assign n4023 = (~x4 | ((~x3 | ~x5 | ~x6 | ~x0 | x2) & (x6 | ((~x0 | (x2 ? (~x3 | x5) : (x3 | ~x5))) & (x0 | ~x2 | x3 | ~x5))))) & (x0 | x2 | x4 | x5 | (~x3 ^ ~x6));
  assign n4024 = (~x2 | ~x3 | x4 | x5 | ~x6) & (x2 | ((x3 | x4 | ~x5 | ~x6) & (x5 | x6 | ~x3 | ~x4)));
  assign n4025 = x1 ? ((~x2 | x3 | x4 | ~x5 | x6) & (~x4 | x5 | ~x6 | x2 | ~x3)) : (x2 ? (~x4 | (x3 ? (x5 | x6) : (~x5 | ~x6))) : (x3 | x4 | (~x5 ^ x6)));
  assign n4026 = (x4 | ~x5 | x6 | ~x1 | x2 | x3) & (x1 | ((x2 | ((~x5 | ~x6 | x3 | ~x4) & (x5 | x6 | ~x3 | x4))) & (~x2 | ~x3 | ~x4 | x5 | ~x6)));
  assign n4027 = (x4 | ((x3 | ((x0 | ~x1 | ~x2 | x5) & (~x0 | (x1 ? (x2 | x5) : ~x2)))) & (x0 | ~x3 | ((x1 | (~x2 & ~x5)) & (~x2 | ~x5))))) & (x1 | ((x0 | x2 | ~x3 | ~x4) & (~x0 | ~x2 | (x3 ? (~x4 | ~x5) : x5)))) & (x0 | ~x4 | ((x2 | ~x3 | ~x5) & (~x1 | (x2 ? ~x3 : (x3 | x5)))));
  assign z344 = n4030 | ~n4036 | (~x2 & ~n4033) | (x0 & ~n4029);
  assign n4029 = (~x1 | x2 | x3 | x4 | ~x5 | ~x6) & (x1 | ((~x5 | x6 | x3 | x4) & (~x3 | x5 | (x2 ? (x4 ^ x6) : (x4 | ~x6)))));
  assign n4030 = x2 & ((~x1 & ~n4032) | (~x0 & x1 & ~n4031));
  assign n4031 = (~x3 | x4 | x5 | ~x6 | ~x7) & (~x5 | x6 | x7 | x3 | ~x4);
  assign n4032 = (~x5 | x6 | ~x7 | x0 | x3 | ~x4) & (~x3 | x5 | ((x4 | ~x6 | x7) & (~x0 | ~x4 | x6 | ~x7)));
  assign n4033 = (~x5 | x7 | n4034 | ~x0 | x3) & (~x3 | (n4035 & (~x7 | n4034 | x0 | x5)));
  assign n4034 = x1 ? (~x4 | x6) : (x4 | ~x6);
  assign n4035 = (x0 | ~x1 | x4 | x5 | ~x6 | x7) & (x1 | ~x4 | ((x5 | x6 | x7) & (~x6 | ~x7 | ~x0 | ~x5)));
  assign n4036 = ~n4038 & (x0 ? n4037 : n4039);
  assign n4037 = (x2 | ((x4 | ~x5 | x1 | ~x3) & (~x4 | x5 | ~x1 | x3))) & (x1 | ((x3 | x4 | x5) & (~x2 | ~x4 | ~x5)));
  assign n4038 = ~x0 & (((x1 ^ ~x2) & (x3 ? (~x4 & x5) : (x4 & ~x5))) | (x1 & ~x2 & x4 & x5) | (~x1 & x2 & (x3 ? (x4 & x5) : (~x4 & ~x5))));
  assign n4039 = ((x4 ^ x6) | ((~x1 | x2 | ~x3 | x5) & (x1 | ~x2 | (~x3 ^ x5)))) & (x1 | x2 | x3 | x4 | ~x5 | ~x6) & (~x1 | ~x2 | ((~x5 | ~x6 | x3 | x4) & (x5 | x6 | ~x3 | ~x4)));
  assign z345 = ~n4047 | (x3 ? (~n4042 | (x7 & ~n4041)) : ~n4043);
  assign n4041 = (x0 | ~x1 | x2 | x4 | x5 | ~x6) & (~x4 | ((x5 | x6 | x0 | x2) & (~x0 | x1 | ((x5 | x6) & (x2 | ~x5 | ~x6)))));
  assign n4042 = (x1 | ~x2 | n2351) & (x0 | ((~x2 | n2351) & (x1 | (n2351 & (~x2 | ~n1449 | ~n544)))));
  assign n4043 = n4046 & (x2 | n4044) & (n1041 | n4045);
  assign n4044 = (~x6 | ((x0 | ~x1 | x4 | ~x5 | ~x7) & (x7 | ((x0 | ~x1 | ~x4 | ~x5) & (~x0 | x1 | (~x4 ^ ~x5)))))) & (x0 | x5 | x6 | (x1 ? (~x4 | x7) : (x4 | ~x7)));
  assign n4045 = (~x2 | x5 | x7 | x0 | ~x1) & (x1 | ((x5 | x7 | x0 | x2) & (~x0 | (x2 ? (x5 | x7) : (~x5 | ~x7)))));
  assign n4046 = x0 ? (~x1 | x2 | (~n686 & ~n1163)) : (~x2 | (~n1163 & (x1 | ~n686)));
  assign n4047 = x3 ? ((n1799 | n850) & (~n3290 | ~n534)) : n4048;
  assign n4048 = (x2 | (x0 ? ((x5 | x6) & (~x1 | ~x5 | ~x6)) : ((~x4 | ~x5 | x6) & (~x1 | x4 | x5)))) & (~x5 | ~x6 | x0 | x1) & (~x2 | (((x0 & x1) | ((~x5 | ~x6) & (x4 | x5 | x6))) & (x1 | (x0 ? (~x4 | ~x5) : (x5 | x6)))));
  assign z346 = ~n4055 | (x0 ? ~n4050 : (x2 ? ~n4054 : ~n4053));
  assign n4050 = (~x4 | n4051) & (x1 | x4 | n4052);
  assign n4051 = (~x1 | x2 | x3 | ~x6 | x7) & (x1 | ((~x6 | ~x7 | x2 | ~x5) & (x5 | (~x2 & ~x3) | (~x6 ^ x7))));
  assign n4052 = (x2 | ~x5 | ~x6 | (~x3 ^ x7)) & (x5 | ((~x3 | x6 | x7) & (~x2 | ((x6 | x7) & (x3 | ~x6 | ~x7)))));
  assign n4053 = (x3 | ~x5 | ((~x1 | (x4 ? (~x6 | ~x7) : (x6 | x7))) & (~x6 | x7 | x1 | x4))) & (~x7 | ((x1 | ((~x3 | ~x4 | x6) & (x4 | x5 | ~x6))) & (x5 | ((~x4 | x6) & (~x3 | x4 | ~x6))))) & (x5 | x7 | ((~x4 | ~x6) & (~x3 | x4 | x6)));
  assign n4054 = (x3 | x5 | x6 | ((x4 | x7) & (~x1 | ~x4 | ~x7))) & (~x6 | ((~x4 | x5 | x7) & (~x3 | ((~x4 | x7) & (~x5 | ~x7 | x1 | x4)))));
  assign n4055 = ~n4058 & n4059 & (x4 ? (x1 | n4057) : n4056);
  assign n4056 = (x2 | (x0 ? ((x1 | x5 | (x3 ^ x6)) & (~x5 | ~x6 | ~x1 | x3)) : ((~x3 | ~x5 | ~x6) & (x5 | x6 | ~x1 | x3)))) & (x0 | ~x2 | ((~x3 | x5 | x6) & (~x5 | ~x6 | x1 | x3)));
  assign n4057 = (x0 | x2 | x3 | ~x5 | x6) & (~x0 | ((~x2 | x3 | ~x5 | x6) & (x2 | (x3 ? (~x5 | x6) : (x5 | ~x6)))));
  assign n4058 = (n616 | n1415 | n1180) & (n1163 | (~x4 & ~n1215));
  assign n4059 = (x0 | ~x1 | x2 | ~x4 | ~x5 | x6) & (x4 | ((~x2 | ~x5 | ~x6 | x0 | ~x1) & (~x0 | ((~x5 | ~x6 | x1 | ~x2) & (~x1 | x2 | x5 | x6)))));
  assign z347 = (~x0 & ~n4061) | (~n846 & ~n4064) | ~n4067 | (x0 & ~n4065);
  assign n4061 = x1 ? n4063 : n4062;
  assign n4062 = (~x4 | ((x2 | ((~x6 | x7 | ~x3 | ~x5) & (x6 | ~x7 | x3 | x5))) & (~x6 | ~x7 | ~x2 | x5))) & (~x2 | ~x7 | ((~x5 | x6 | (x3 & x4)) & (~x3 | x5 | ~x6)));
  assign n4063 = (x4 | ((x2 | ~x3 | x5 | x6 | ~x7) & (~x2 | x3 | ~x5 | ~x6 | x7))) & (~x2 | ~x3 | (x5 ? (x6 | ~x7) : ((~x6 | ~x7) & (~x4 | x6 | x7))));
  assign n4064 = x0 ? ((~x1 | x2 | x3 | x4 | x7) & (x1 | ~x3 | (~x2 ^ x7))) : ((~x1 | ((~x4 | ~x7 | x2 | x3) & (x4 | x7 | ~x2 | ~x3))) & (x3 | ((~x2 | ~x4 | x7) & (x1 | (x2 ? x7 : (x4 | ~x7))))));
  assign n4065 = (x1 | n4066) & (~x1 | x2 | x3 | ~x7 | n912);
  assign n4066 = (~x3 | ((x5 | ~x6 | x7 | x2 | x4) & (~x2 | ~x4 | ~x5 | x6 | ~x7))) & (x2 | x3 | ~x7 | (x4 ? (~x5 | ~x6) : (~x5 ^ x6)));
  assign n4067 = ~n4069 & ~n4070 & n4071 & (~x7 | n4068);
  assign n4068 = (x0 | ((~x3 | ~x4 | ~x5 | x1 | ~x2) & (~x1 | x2 | (x3 ? (~x4 | x5) : (x4 | ~x5))))) & (x1 | ~x2 | x5 | ((x3 | x4) & (~x0 | ~x3 | ~x4)));
  assign n4069 = ~x1 & ((x3 & ((x5 & ~x7 & x0 & ~x2) | (~x0 & ~x5 & (x2 ^ x7)))) | (x0 & ~x3 & ~x7 & (~x2 ^ x5)));
  assign n4070 = ~x7 & n897 & ((x1 & ~n2241) | (n1449 & n605));
  assign n4071 = x3 ? (x4 | n4072) : ((~n1156 | ~n750) & (~x4 | n4072));
  assign n4072 = (~x5 | x7 | x0 | x2) & (~x0 | x5 | (x1 ? (x2 | x7) : (~x2 | ~x7)));
  assign z348 = n4074 | n4076 | (x2 ? ~n4080 : ~n4079);
  assign n4074 = x1 & ((n559 & n2314) | (~x0 & ~n4075));
  assign n4075 = x4 ? (x7 | ((~x5 | x6 | x2 | x3) & (~x2 | ~x3 | (~x5 ^ x6)))) : ((x2 | ~x3 | x5 | ~x6 | ~x7) & (x3 | ((~x6 | ~x7 | x2 | ~x5) & (~x2 | x7 | (~x5 ^ ~x6)))));
  assign n4076 = ~x1 & (x5 ? ~n4078 : ~n4077);
  assign n4077 = x4 ? ((x0 | x2 | ~x3 | x6 | x7) & (~x7 | (~x0 ^ x6) | (~x2 ^ ~x3))) : ((x0 | ~x2 | x3 | x6 | ~x7) & (~x0 | x2 | ~x3 | ~x6 | x7));
  assign n4078 = (x0 | ~x2 | ~x3 | x4 | x6 | x7) & (x3 | ((~x4 | ((x6 | ~x7 | x0 | x2) & (~x0 | ~x6 | (x2 & x7)))) & (x0 | x4 | (x2 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n4079 = x6 ? ((~x0 | (x1 ? (x3 | x4) : (~x3 | ~x7))) & (~x4 | ~x7 | ~x1 | x3) & (x1 | ((x3 | x4 | ~x7) & (~x4 | x7 | x0 | ~x3)))) : ((x0 | ((~x1 | (x3 ? x7 : x4)) & (~x3 | (x7 ? (x1 & ~x4) : x4)))) & (x7 | ((x1 | x3 | ~x4) & (~x0 | ((x3 | ~x4) & (x1 | (x3 & ~x4)))))));
  assign n4080 = x0 ? (x1 | ((~x3 | ~x6 | (~x4 & x7)) & (x6 | (x3 & (x4 | ~x7))))) : (x6 ? (x3 ? ((x4 | ~x7) & (~x1 | (x4 & ~x7))) : ((~x4 | x7) & (x1 | (~x4 & x7)))) : ((~x1 | x3 | ~x7) & (~x4 | x7 | x1 | ~x3)));
  assign z349 = ~n4088 | n4087 | n4086 | n4084 | n4082 | n4083;
  assign n4082 = ~x0 & (x1 ? (x2 ? (x3 ? (~x4 & ~x7) : (x4 & x7)) : (~x7 & (x3 ^ ~x4))) : ((x4 & ~x7 & x2 & ~x3) | (~x2 & (x3 ? (~x4 ^ x7) : (~x4 & x7)))));
  assign n4083 = ~n1007 & ((x2 & ~x4 & ~x7 & ~x0 & ~x1) | (x0 & x7 & (x1 ? (~x2 & ~x4) : (x2 & x4))));
  assign n4084 = ~n4085 & ~x7 & n738;
  assign n4085 = x2 ? ((x5 | ~x6 | ~x3 | ~x4) & (x3 | (x4 ? (~x5 | x6) : (x5 | ~x6)))) : ((~x3 | x4 | ~x5 | x6) & (x5 | ~x6 | x3 | ~x4));
  assign n4086 = x0 & ((x3 & ~x4 & x7 & ~x1 & x2) | (~x2 & ((x4 & x7 & ~x1 & x3) | (~x3 & (x1 ? (~x4 ^ x7) : (~x4 & x7))))));
  assign n4087 = n664 & ((x7 & ((~x2 & x3 & ~x4 & ~x5) | (x5 & (x2 ? (x3 ^ ~x4) : (~x3 & x4))))) | (x2 & ~x5 & ~x7 & (x3 ^ ~x4)));
  assign n4088 = (x1 | n4089) & (x0 | (~n4091 & (~x4 | n4090)));
  assign n4089 = x2 ? (((~x4 ^ x5) | (x0 ? (x3 | x7) : (~x3 | ~x7))) & (x0 | x3 | x4 | x5 | ~x7) & (~x0 | ~x3 | ~x4 | ~x5 | x7)) : ((~x0 | ~x3 | x4 | (x5 ^ x7)) & (x3 | ~x4 | ((~x5 | x7) & (x0 | x5 | ~x7))));
  assign n4090 = (x1 | ~x2 | ~x3 | ~x5 | (~x6 ^ x7)) & (x2 | x5 | ((~x1 | x3 | (x6 ^ x7)) & (x6 | x7 | x1 | ~x3)));
  assign n4091 = n733 & ((~x1 & x2 & x3 & n1120) | (x1 & (x2 ? (~x3 & n1120) : (x3 & n1121))));
  assign z350 = n4095 | ~n4096 | (~x4 & (n4094 | (~x7 & ~n4093)));
  assign n4093 = ((x0 ? (x1 | x6) : (~x1 | ~x6)) | (x2 ? (x3 | x5) : (~x3 | ~x5))) & (x3 | ~x5 | x6 | x0 | x1 | ~x2) & (~x0 | ~x1 | x2 | ~x6 | (~x3 ^ x5));
  assign n4094 = n549 & ((~x0 & ~x1 & x3 & ~x5 & x6) | (~x3 & ((x5 & ~x6 & ~x0 & x1) | (x0 & ~x5 & (x1 ^ x6)))));
  assign n4095 = n664 & (x4 ? ((x2 & (x3 ^ x5)) | (~x5 & ~x6 & ~x2 & ~x3)) : ((~x2 & (x3 ? ~x5 : (x5 & x6))) | (x5 & x6 & x2 & x3)));
  assign n4096 = ~n4099 & ~n4100 & (~n2326 | n4098) & (x1 | n4097);
  assign n4097 = x2 ? ((~x0 | (x3 ? (x4 | ~x5) : (~x4 | x6))) & (x3 | ~x4 | ~x5 | x6) & (x0 | x5 | (x3 ? (~x4 | x6) : x4))) : (x0 ? ((~x5 | ~x6 | x3 | x4) & (~x3 | (~x4 ^ ~x5))) : ((x3 | ~x4 | x5) & (~x5 | ~x6 | ~x3 | x4)));
  assign n4098 = (x6 | (~x0 ^ x3) | (x1 ? (~x5 | ~x7) : (x5 | x7))) & (x1 | ~x3 | ~x6 | ~x7 | (~x0 ^ x5));
  assign n4099 = ~n783 & ((n616 & n2417) | (n2573 & (n610 | n1743)));
  assign n4100 = ~n1323 & (x0 ? (~x5 & (x1 ? n1148 : n710)) : (~x1 & x5 & (n710 | n1148)));
  assign z351 = n4102 | ~n4105 | (n1317 & ~n4112) | (~x2 & ~n4111);
  assign n4102 = ~x3 & (n4104 | (~x1 & ~n4103));
  assign n4103 = x2 ? ((x4 ? (~x6 | ~x7) : (x6 | x7)) | (~x0 ^ x5)) : (x5 | ((~x6 | ~x7 | x0 | x4) & (~x0 | x7 | (~x4 ^ x6))));
  assign n4104 = n664 & ((~x2 & x4 & x5 & ~x6 & x7) | (~x4 & ((x6 & ~x7 & x2 & ~x5) | (~x2 & x5 & (x6 ^ ~x7)))));
  assign n4105 = ~n4106 & ~n4108 & (n846 | n4110) & (~x2 | n4107);
  assign n4106 = ~n850 & (n720 | (~x0 & (n1386 | n758)));
  assign n4107 = ((x5 ^ x6) | ((~x0 | x1 | ~x3 | ~x4) & (x0 | (x1 ? x3 : (~x3 | x4))))) & (x0 | x3 | ~x4 | x5 | x6) & (x1 | (x0 ? ((x5 | ~x6 | ~x3 | x4) & (x3 | ~x5 | (x4 & x6))) : ((~x5 | x6 | ~x3 | ~x4) & (x3 | x5 | ~x6))));
  assign n4108 = ~n4109 & (x1 ? ~n1477 : (x3 & ~n850));
  assign n4109 = x0 ? (x2 | x7) : (~x2 | ~x7);
  assign n4110 = x0 ? (x4 | ((~x3 | ~x7 | x1 | ~x2) & (~x1 | x2 | x3 | x7))) : (x1 | x2 | ~x4 | (~x3 ^ x7));
  assign n4111 = ((x5 ^ x6) | ((x3 | ~x4 | x0 | ~x1) & (x1 | (x0 ? (~x3 ^ ~x4) : (~x3 | x4))))) & (x0 | ((~x1 | x3 | x4 | x5 | ~x6) & (x1 | ~x3 | ~x4 | ~x5 | x6))) & (~x0 | ((~x1 | ~x3 | x4 | x5 | x6) & (x1 | ((x3 | ~x4 | ~x5 | x6) & (x5 | ~x6 | ~x3 | x4)))));
  assign n4112 = (x5 | ~x6 | x7 | x1 | x2 | x4) & (~x1 | ((~x2 | ~x4 | x5 | x6 | ~x7) & (x2 | ~x5 | x7 | (~x4 ^ x6))));
  assign z352 = ~n4119 | (x1 ? (n4114 | (~x0 & ~n4118)) : ~n4115);
  assign n4114 = n2314 & n686;
  assign n4115 = (~x7 | n4116) & (x0 | x7 | n4117);
  assign n4116 = x2 ? (x0 ? ((~x5 | ~x6 | x3 | x4) & (x5 | x6 | ~x3 | ~x4)) : (x4 ? (x3 ? (~x5 | x6) : (x5 | ~x6)) : (x5 | x6))) : (x6 | (x0 ? (x3 ? (x4 | x5) : ~x5) : (x4 | ~x5)));
  assign n4117 = (x2 | ~x5 | ((~x4 | ~x6) & (x3 | x4 | x6))) & (~x4 | x5 | ~x6 | (~x2 & ~x3));
  assign n4118 = (~x6 | ((x4 | x5 | ~x7 | x2 | ~x3) & (~x2 | ~x4 | ~x5 | (~x3 & x7)))) & (x2 | x3 | ((x5 | x6 | ~x7) & (x4 | ~x5 | x7))) & (~x5 | x6 | ~x7 | ~x2 | x4);
  assign n4119 = (~x6 | (x7 ? n4120 : n4121)) & (n1311 | n4122) & (x6 | (x7 ? n4121 : n4120));
  assign n4120 = (x2 & ((x0 & (x1 | (~x4 & x5))) | (x1 & x3 & x5) | (~x5 & ((~x1 & x4) | (~x0 & ~x3 & ~x4))))) | (~x2 & (x4 ? ((x0 & x3) | (~x1 & x5) | (x1 & ~x3 & ~x5)) : ((~x0 & (x3 ^ x5)) | (~x1 & ~x3 & ~x5)))) | (x1 & ~x4 & (x3 | x5)) | (x4 & x5 & ~x0 & ~x1);
  assign n4121 = x1 ? (x4 | ((x3 | ~x5 | ~x0 | x2) & (x0 | ~x3 | (~x2 ^ x5)))) : ((x3 | ~x4 | ~x5 | x0 | ~x2) & (x5 | ((~x0 | ~x4 | (~x2 ^ x3)) & (x2 | x4 | (x0 & x3)))));
  assign n4122 = (~x0 | x1 | ~x5 | (~x2 & ~x3)) & (~x1 | x5 | (x0 ? (x2 | x3) : (~x2 ^ x3)));
  assign z353 = ~n4126 | (~x2 & (x5 ? ~n4125 : ~n4124));
  assign n4124 = x3 ? ((~x6 | ~x7 | x0 | x1) & (~x0 | ((x1 | ~x6 | x7) & (x6 | ~x7 | ~x1 | x4)))) : ((~x0 | ((x1 | ~x6 | ~x7) & (x6 | x7 | ~x1 | ~x4))) & (~x6 | ~x7 | x1 | ~x4) & (x0 | x4 | ((~x6 | x7) & (~x1 | x6 | ~x7))));
  assign n4125 = (x0 | ~x1 | x3 | x4 | x6 | x7) & (x1 | ((~x7 | (x0 ? (x3 | (~x4 ^ ~x6)) : (x6 | (~x3 & ~x4)))) & (~x3 | x7 | (x0 ? x6 : (x4 | ~x6)))));
  assign n4126 = ~n4130 & (n846 | n4129) & (x1 ? n4128 : n4127);
  assign n4127 = (~x0 | ((~x2 | x4 | (x3 ? (x5 | x7) : (~x5 | ~x7))) & (x3 | ~x4 | x5 | x7) & (x2 | ((x3 | x5 | x7) & (~x5 | ~x7 | ~x3 | ~x4))))) & (x2 | x3 | ~x4 | x5 | x7) & (x0 | ((x4 | ((~x5 | x7 | ~x2 | ~x3) & (x2 | (x3 ? (x5 | x7) : (~x5 | ~x7))))) & (~x2 | x3 | ((x5 | ~x7) & (~x4 | ~x5 | x7)))));
  assign n4128 = (~x3 | ~x5 | ~x7 | x0 | ~x2) & (x2 | ((x3 | ((~x4 | x5 | ~x7) & (~x0 | ((x5 | ~x7) & (~x4 | ~x5 | x7))))) & (x0 | ~x3 | ((~x5 | x7) & (x4 | x5 | ~x7)))));
  assign n4129 = x1 ? ((x3 | x4 | x7 | ~x0 | x2) & (x0 | (x2 ? (x3 | ~x7) : (~x4 | (x3 ^ x7))))) : ((x0 | ~x2 | x3 | x4 | x7) & (~x3 | (x0 ? (x2 ? (~x4 | x7) : (x4 | ~x7)) : (x2 ? ~x7 : (~x4 | x7)))));
  assign n4130 = x2 & ((~n912 & ~n4131) | (~x7 & ~n4132));
  assign n4131 = x0 ? (x1 | ~x7 | (~x3 & ~x4)) : (~x1 | x7 | (~x3 ^ x4));
  assign n4132 = (x0 | ~x1 | ((~x5 | x6 | x3 | x4) & (x5 | ~x6 | ~x3 | ~x4))) & (x1 | ((x0 | ~x3 | ~x4 | ~x5 | x6) & (~x0 | x4 | ~x6 | (x3 ^ x5))));
  assign z354 = ~n4137 | (x0 & ~x2 & ~n4134) | (~x0 & (~n4136 | (~x2 & ~n4135)));
  assign n4134 = (x5 | x7 | ((x1 | x3 | ~x4 | ~x6) & (~x1 | (x3 ? (x4 | ~x6) : (~x4 | x6))))) & (x1 | x4 | ~x5 | ~x7 | (x3 ^ x6));
  assign n4135 = (x1 | ~x3 | x4 | x5 | ~x6 | x7) & (~x5 | ((x1 | ~x3 | x4 | x6 | x7) & (~x7 | (x1 ? (x3 ? (~x4 | x6) : (x4 | ~x6)) : (~x4 | (x3 ^ x6))))));
  assign n4136 = x1 ? ((~x2 | x3 | x4 | x6 | ~x7) & (x2 | ~x3 | ~x4 | ~x6 | x7)) : ((x2 | x3 | ~x4 | ~x6 | x7) & (~x3 | ((x6 | ~x7 | x2 | x4) & (~x2 | (x4 ? (x6 | ~x7) : (~x6 | x7))))));
  assign n4137 = ~n4141 & n4142 & (~x2 | (~n4138 & ~n4140));
  assign n4138 = ~n4139 & (n1897 | (x4 & n723));
  assign n4139 = (x3 | ~x6 | x0 | ~x1) & (~x0 | x1 | (~x3 ^ ~x6));
  assign n4140 = n1317 & (x1 ? (x4 & n1902) : (n762 | n1231));
  assign n4141 = ~n662 & ((~x2 & ((x0 & (x1 ? (~x3 & ~x4) : (x3 & x4))) | (~x3 & x4 & ~x0 & x1))) | (~x0 & x2 & ~x4 & (~x1 ^ x3)));
  assign n4142 = n4143 & (~n738 | (x2 ? n1306 : (x3 | n1311)));
  assign n4143 = x1 ? ((x3 | ~x4 | ~x6 | ~x0 | x2) & (x0 | (x3 ^ x6) | (x2 ^ x4))) : (((x3 ? (~x4 | x6) : (x4 | ~x6)) | (x0 ^ x2)) & (x3 | ~x4 | ~x6 | x0 | ~x2) & (~x3 | x4 | x6 | ~x0 | x2));
  assign z355 = ~n4149 | (x1 ? ~n4145 : (n4147 | (~x6 & ~n4148)));
  assign n4145 = (x6 | n4146) & (x0 | ~n665 | ~n762);
  assign n4146 = (x2 | ((x0 | x3 | x4 | ~x5 | ~x7) & (x5 | ((~x4 | ~x7 | x0 | ~x3) & (~x0 | (x3 ? (x4 | ~x7) : (~x4 | x7))))))) & (x0 | ~x2 | ((x3 | ~x5 | (x4 ^ x7)) & (x5 | x7 | ~x3 | ~x4)));
  assign n4147 = ~n2354 & ((~x2 & ((~x6 & x7 & x0 & ~x4) | (~x0 & x4 & (x6 ^ x7)))) | (x0 & x2 & ~x6 & (~x4 ^ x7)));
  assign n4148 = (x0 | ~x2 | ~x3 | (x4 ? (~x5 | x7) : (x5 | ~x7))) & (~x0 | x2 | x3 | ~x4 | ~x5 | x7);
  assign n4149 = n4151 & ((x0 & (x1 | (n4152 & n4153))) | (n4150 & (x1 | (~x0 & n4152))));
  assign n4150 = x2 ? (((x5 ^ x7) | (x1 ? (x3 | x4) : (~x3 | ~x4))) & (x4 | ~x5 | x7 | x1 | ~x3) & (~x4 | x5 | ~x7 | ~x1 | x3)) : (x1 ? ((x5 | ~x7 | x3 | x4) & (~x5 | x7 | ~x3 | ~x4)) : ((~x4 | (x3 ? (x5 | ~x7) : (~x5 | x7))) & (~x3 | x4 | (x5 ^ x7))));
  assign n4151 = ((x4 ^ x7) | ((~x0 | ~x1 | x2 | x3) & (x0 | ~x2 | (x1 ^ x3)))) & (x0 | ~x1 | x2 | (x3 ? (x4 | ~x7) : (~x4 | x7)));
  assign n4152 = (~x0 | ((~x4 | x7 | x2 | ~x3) & (~x2 | x3 | x4 | ~x7))) & (x0 | x2 | x3 | x4 | ~x7);
  assign n4153 = ((x2 ? (~x3 | x4) : (x3 | ~x4)) | (~x5 ^ ~x7)) & ((x2 ^ x4) | (x3 ? (x5 | ~x7) : (~x5 | x7)));
  assign z356 = ~n4158 | (x2 & ~n4157) | (x1 & (n4156 | (~x2 & ~n4155)));
  assign n4155 = (x5 | ((x0 | x3 | ~x4 | ~x6 | ~x7) & (~x0 | x7 | (x3 ? (x4 | ~x6) : (~x4 | x6))))) & (x0 | ~x5 | ((x3 | x4 | ~x6 | x7) & (~x3 | ~x7 | (x4 ^ x6))));
  assign n4156 = ~x7 & n616 & ((x3 & x4 & ~x5 & ~x6) | (~x3 & x5 & (~x4 ^ x6)));
  assign n4157 = (x1 | (x0 ? ((~x5 | ~x6 | x3 | x4) & (x6 | (x3 ? (~x4 ^ ~x5) : (~x4 | x5)))) : ((~x5 | x6 | x3 | x4) & (x5 | ~x6 | ~x3 | ~x4)))) & (x0 | ~x1 | x6 | (x3 ? (x4 | ~x5) : (~x4 ^ ~x5)));
  assign n4158 = n4163 & (x2 | n4159) & (x1 | (~n4160 & n4161));
  assign n4159 = x4 ? ((x1 | (x3 ^ x5) | (x0 ^ x6)) & (x0 | ~x1 | (x3 ? (x5 | x6) : (~x5 | ~x6)))) : (x1 ? (x0 ? (x6 | (~x3 ^ x5)) : (~x6 | (x3 ^ x5))) : ((x0 | (x3 ? (x5 | x6) : (~x5 | ~x6))) & (~x0 | ~x3 | x5 | ~x6)));
  assign n4160 = ~n783 & ((~x0 & ~x2 & ~x3 & x5 & x7) | (x0 & x2 & ~x7 & (x3 ^ ~x5)));
  assign n4161 = (x2 | ~x3 | n4162) & (n1019 | ((~x0 | x2 | x3 | x7) & (x0 | ~x2 | (~x3 ^ x7))));
  assign n4162 = (x0 | ~x4 | x5 | x6 | ~x7) & (~x0 | x4 | ~x5 | ~x6 | x7);
  assign n4163 = ((x2 ? (x5 | ~x6) : (~x5 | x6)) | (x0 ? (x1 | ~x3) : (~x1 | x3))) & ((x1 ? (~x5 | ~x6) : (x5 | x6)) | (x0 ? (x2 | x3) : (~x2 | ~x3))) & (x0 | x1 | ~x6 | (x2 ? (x3 | ~x5) : (~x3 | x5)));
  assign z357 = ~n4169 | (~n620 & ~n4165) | (~x2 & ~n4166);
  assign n4165 = x2 ? ((x1 | (x0 ? (~x4 | (x3 & ~x5)) : (x4 | (~x3 & x5)))) & (x0 | ((~x3 | x4 | x5) & (~x4 | ~x5 | ~x1 | x3)))) : (((~x4 ^ x5) | (x0 ? (x1 | ~x3) : (~x1 | x3))) & ((x1 ^ x3) | (x0 ? (x4 | x5) : (~x4 | ~x5))));
  assign n4166 = n4168 & (x1 | n4167) & (n1215 | (~n1035 & ~n2010));
  assign n4167 = (x3 | (x0 ? ((x6 | x7 | x4 | x5) & (~x6 | ~x7 | ~x4 | ~x5)) : (~x5 | ((x6 | x7) & (x4 | ~x6 | ~x7))))) & (~x0 | ~x3 | ((x4 | ~x5 | x6 | x7) & (~x6 | ~x7 | ~x4 | x5)));
  assign n4168 = (~x0 | ~x1 | x3 | n1451) & (x0 | (x1 ? (x3 | ~n1846) : (~x3 | n1451)));
  assign n4169 = x2 ? (n4170 & n4173) : n4172;
  assign n4170 = (x1 | n4171) & (x0 | ~x1 | (n4031 & (n662 | n2136)));
  assign n4171 = x0 ? ((x4 | ((x5 | ~x6 | ~x7) & (x6 | x7 | ~x3 | ~x5))) & (x3 | ((x5 | x6 | x7) & (~x6 | ~x7 | ~x4 | ~x5)))) : ((~x4 | ((~x5 | x6 | x7) & (~x6 | ~x7 | x3 | x5))) & (~x3 | ((~x5 | ~x6 | ~x7) & (x6 | x7 | x4 | x5))));
  assign n4172 = ((x0 ? (x1 | ~x3) : (~x1 | x3)) | (x4 ? (~x5 | ~x6) : (x5 | x6))) & ((~x1 ^ x5) | ((~x4 | x6 | x0 | ~x3) & (x4 | ~x6 | ~x0 | x3))) & (~x4 | ~x5 | x6 | ~x0 | ~x1 | x3) & (x0 | x1 | x5 | ((x4 | ~x6) & (x3 | ~x4 | x6)));
  assign n4173 = (x1 | (x3 ? (~x4 | x5) : (x4 | ~x5)) | (x0 ^ ~x6)) & (x0 | ~x1 | (~x4 ^ x6) | (x3 ^ x5));
  assign z358 = ~n4178 | (~x2 & (~n4176 | (~x3 & ~n4175) | ~n4177));
  assign n4175 = (x0 | ((x1 | x4 | x5 | x6 | ~x7) & (~x5 | ((~x6 | x7 | x1 | ~x4) & (~x1 | (x4 ? (x6 | x7) : ~x6)))))) & (x5 | x7 | ((~x1 | x4 | x6) & (~x0 | x1 | ~x6)));
  assign n4176 = (x0 | x1 | ~x3 | ~n1163) & (n1002 | ((~x0 | x3 | (x1 ^ x6)) & (~x3 | ((x1 | ~x6) & (x0 | ~x1 | x6)))));
  assign n4177 = (x3 | ((x4 | ~x5 | x7 | x0 | x1) & ((~x4 ^ x7) | (x0 ? (x1 | ~x5) : (~x1 | x5))))) & (x1 | ~x3 | ((x4 | x5 | ~x7) & (~x0 | ~x4 | (x5 ^ x7))));
  assign n4178 = ~n4180 & ~n4181 & (n824 | n4183) & (~x2 | n4179);
  assign n4179 = ((~x5 ^ x7) | ((x1 | ~x3 | ~x4) & (x0 | ~x1 | x3 | x4))) & (x1 | x3 | x4 | x5 | x7) & (~x4 | ~x5 | ~x7 | x0 | ~x1 | ~x3);
  assign n4180 = ~n906 & (x1 ? ((~x4 & ~x5 & x0 & ~x2) | (~x0 & x4 & (x2 ^ x5))) : ((x2 & ~x4 & x5) | (x4 & ~x5 & ~x0 & ~x2)));
  assign n4181 = ((~x1 & ~x6) | (~x0 & x1 & x6)) & (n4182 | (x2 & ~n3065));
  assign n4182 = ~x2 & x3 & ~x4 & (x5 ^ ~x7);
  assign n4183 = (x3 | ~x4 | x6 | ~x0 | ~x1 | x2) & (~x2 | (~x3 ^ x4) | ((x1 | ~x6) & (x0 | ~x1 | x6)));
  assign z359 = ~n4189 | (x5 ? ~n4185 : (x3 ? ~n4188 : ~n4187));
  assign n4185 = x2 ? (x4 | n1799 | (~n869 & ~n3900)) : n4186;
  assign n4186 = x3 ? (~x4 | ((x1 | x6 | x7) & (x0 | ((x6 | x7) & (x1 | ~x6 | ~x7))))) : (x7 ? ((~x0 | ((x4 | x6) & (~x1 | ~x4 | ~x6))) & (x6 | (x4 ? (x0 & x1) : ~x1))) : ((x1 | ~x4 | ~x6) & (x0 | (x1 ? ~x6 : (x4 | x6)))));
  assign n4187 = (x0 & ((x6 & x7) | (x1 & x4))) | (~x4 & (x2 | (~x0 & ~x1 & (~x6 | ~x7)))) | (~x6 & ~x7) | (x1 & x6 & x7) | (x4 & (~x2 | (x6 & x7)));
  assign n4188 = (x0 | ~x2 | ~x4 | x6 | x7) & (x2 | ((~x0 | ~x1 | x4 | x6 | x7) & (~x7 | (x0 & x1) | (~x4 ^ ~x6))));
  assign n4189 = ~n4190 & ~n4191 & (~n1317 | (~x2 & ~n2237) | (x2 & n1019));
  assign n4190 = ~x3 & ((~x2 & ((~x5 & ~x6 & ~x0 & x4) | (x0 & x6 & (x4 ^ x5)))) | (~x0 & x2 & (x4 ? (x5 & x6) : ~x6)));
  assign n4191 = n738 & ((x3 & (x2 ? (x4 & ~x6) : (~x4 & x6))) | (x2 & ((x6 & ~n2500) | (~x3 & ~x4 & ~x6))));
  assign z360 = ~n4197 | (~n800 & ~n4196) | (~x2 & (n4193 | ~n4194));
  assign n4193 = n1156 & (x1 ? (x0 ? (~x4 & ~x6) : (x3 ? x4 : (~x4 & x6))) : ((x3 & x4 & ~x6) | (x0 & (x3 ^ ~x4))));
  assign n4194 = ~n4195 & (~n3098 | ~n1229) & (~n1449 | ~n544 | ~n1880);
  assign n4195 = ~x0 & ((~x6 & x7 & ~x3 & ~x4) | (x3 & x6 & (x1 ? (~x4 & ~x7) : (x4 & x7))));
  assign n4196 = x3 ? (x6 | ((x1 | x2 | x4) & (x0 | (x2 ^ x4)))) : (x0 ? ((x1 | ~x2 | ~x4) & (~x1 | x2 | x4 | ~x6)) : (~x6 | ((~x2 | ~x4) & (x1 | x2 | x4))));
  assign n4197 = ~n4201 & (n824 | n4200) & (~x2 | (~n4198 & ~n4199));
  assign n4198 = ~x0 & ((x3 & x4 & x5 & x6 & ~x7) | (~x3 & ~x6 & (x4 ? (~x5 & x7) : ~x7)));
  assign n4199 = ~x7 & n738 & (x3 ? (x4 & x5) : (~x4 & ~x6));
  assign n4200 = (x0 & x1 & (x3 | ~x4)) | (x4 & (x2 | (x3 & x6))) | (~x4 & (~x2 | (~x3 & ~x6)));
  assign n4201 = ~n592 & (n4202 | (n2467 & (n616 | n1176)));
  assign n4202 = ~x6 & x5 & ~x3 & x0 & ~x2;
  assign z361 = (x3 & ~n4204) | (~x0 & ~n4207) | ~n4212 | (~x3 & ~n4208);
  assign n4204 = x1 ? n4206 : n4205;
  assign n4205 = (x7 | (x4 ? ((x2 | x5 | x6) & (~x0 | ((x5 | x6) & (x2 | ~x5 | ~x6)))) : (x5 | ~x6 | (x0 & ~x2)))) & (~x2 | ~x5 | ~x7 | ((~x4 | x6) & (x0 | x4 | ~x6)));
  assign n4206 = (x5 | ~x6 | x7 | ~x0 | x2 | x4) & (x0 | (x2 ? ((~x6 | x7 | x4 | x5) & (x6 | ~x7 | ~x4 | ~x5)) : (~x4 | x7 | (~x5 ^ ~x6))));
  assign n4207 = (~x6 | ((x1 | ((~x3 | ~x4 | ~x5) & (x2 | x3 | x4 | x5))) & (~x3 | ~x5 | (x4 ? ~x2 : (~x1 & x2))))) & (~x3 | ~x4 | x6 | (~x2 ^ x5));
  assign n4208 = ~n4209 & ~n4210 & ~n4211 & ((x0 & x2) | n2351 | (~x0 & ~x2));
  assign n4209 = n738 & ((~x2 & ~x4 & x5 & x6 & ~x7) | (x7 & ((~x2 & x4 & x5 & x6) | (x2 & ~x5 & (x4 ^ x6)))));
  assign n4210 = ~x0 & x4 & x7 & ((~x5 & ~x6) | (~x2 & x5 & x6));
  assign n4211 = n924 & n1449 & n544;
  assign n4212 = (~n1021 | ~n4214) & (n4213 | (n1799 & ~n694));
  assign n4213 = (~x3 | x4 | x5 | x6) & (x3 | (x4 ? (x5 | ~x6) : (~x5 | x6)));
  assign n4214 = x5 & ((~x2 & x4 & ~x6) | (x6 & (x2 | ~x4)));
  assign z362 = ~n4218 | (~x4 & (n1916 | n4217 | (~x0 & ~n4216)));
  assign n4216 = (x1 | x3 | x5 | x6 | ~x7) & (x2 | ((~x5 | ((x3 | ~x6 | ~x7) & (x1 | x6 | x7))) & (~x7 | (x1 ? (x3 | ~x6) : (x6 | (x3 & x5))))));
  assign n4217 = ~n857 & ((~x6 & ((x2 & ((~x5 & x7) | (~x3 & x5 & ~x7))) | (x3 & (x5 ? ~x2 : x7)))) | (~x2 & x5 & (x3 ? x7 : (x6 & ~x7))));
  assign n4218 = ~n4219 & ~n4223 & ((x0 & ~n1122) | n4225 | (~x0 & ~n2527));
  assign n4219 = x4 & ((~x3 & ~n4220) | (~n800 & ~n4221) | (x3 & ~n4222));
  assign n4220 = x2 ? (~x5 | ((x1 | ~x6 | ~x7) & (x0 | (x6 ^ x7)))) : ((x7 | (x0 ? (~x5 | (~x1 ^ x6)) : (x5 | (x1 & ~x6)))) & (~x0 | ~x7 | (x1 ? (x5 | ~x6) : (~x5 | x6))));
  assign n4221 = (x1 | ((~x6 | (~x2 ^ x3)) & (~x0 | ((~x3 | ~x6) & (x2 | x3 | x6))))) & (x0 | ((x3 | ~x6) & (~x2 | (x6 ? ~x1 : ~x3))));
  assign n4222 = (x1 | ((~x0 | x7 | (x2 ? (~x5 | x6) : x5)) & (~x6 | ~x7 | ((~x2 | ~x5) & (x0 | (~x2 & ~x5)))))) & (x0 | ~x6 | ~x7 | ((~x2 | ~x5) & (~x1 | x2 | x5)));
  assign n4223 = ~n4224 & (n1621 | (~x4 & ~n630));
  assign n4224 = (x0 & (x2 ? x1 : x3)) | (~x2 & ((x1 & x3) | (~x0 & ~x1 & ~x3)));
  assign n4225 = (x1 | ~x2 | x4 | ~x5 | ~x6) & (~x1 | x2 | ~x4 | (~x5 ^ ~x6));
  assign z365 = n1700 | ~n1702 | n4227 | n4231 | (~n927 & ~n4230);
  assign n4227 = x6 & ((n1119 & ~n4229) | (~x0 & ~n4228));
  assign n4228 = (x4 | ~x5 | x7 | ~x1 | x2 | ~x3) & ((x2 ^ ~x7) | ((x4 | ~x5 | x1 | ~x3) & (~x4 | x5 | ~x1 | x3)));
  assign n4229 = (~x3 | ~x5 | ~x7 | x1 | ~x2) & (x3 | ((x5 | x7 | ~x1 | x2) & (x1 | ((x5 | ~x7) & (x2 | ~x5 | x7)))));
  assign n4230 = (~x0 | x1 | x2 | ~x3 | ~x5 | x6) & (x0 | ~x2 | ((~x5 | x6 | ~x1 | ~x3) & (x5 | ~x6 | x1 | x3)));
  assign n4231 = ~x6 & ((n2205 & n650 & n677) | (~x3 & ~n4232));
  assign n4232 = (x0 | ~x1 | ~x7 | (x2 ? (~x4 | x5) : (x4 | ~x5))) & (~x0 | x1 | ~x4 | x5 | x7);
  assign z366 = ~n1715 | n4235 | (n642 & ~n4234);
  assign n4234 = (~x3 | ~x5 | ~x7 | ~x0 | x1 | x2) & (x0 | ((x1 | x5 | ((x3 | ~x7) & (x2 | ~x3 | x7))) & (~x5 | ((~x1 | (x3 ^ x7)) & (~x2 | ~x3 | ~x7)))));
  assign n4235 = x4 & ((n1365 & ~n4237) | (~x5 & ~n4236));
  assign n4236 = x0 ? (x6 | ((x3 | ~x7 | ~x1 | x2) & (~x3 | x7 | x1 | ~x2))) : (~x6 | ((x1 | ((~x3 | x7) & (~x2 | x3 | ~x7))) & (x2 | ((~x3 | x7) & (~x1 | x3 | ~x7)))));
  assign n4237 = (~x2 | ~x3 | ~x7 | x0 | ~x1) & (~x0 | x1 | ((~x2 | x3 | x7) & (~x3 | ~x7)));
  assign z367 = n4239 | ~n4244 | (x1 & ~n4243) | (~n927 & ~n4242);
  assign n4239 = ~x2 & (x3 ? (~x6 & ~n4241) : ~n4240);
  assign n4240 = (~x0 | x1 | x4 | ~x5 | ~x6 | x7) & (x0 | ((x1 | ~x4 | x5 | x6 | x7) & (~x7 | ((x1 | x4 | x5 | x6) & (~x1 | (x4 ? (x5 | ~x6) : (~x5 | x6)))))));
  assign n4241 = (x4 | x5 | x7 | ~x0 | ~x1) & ((~x4 ^ x7) | (x0 ? (x1 | ~x5) : (x1 ^ x5)));
  assign n4242 = (~x1 | ((x3 | x5 | x6 | ~x0 | x2) & (~x3 | ~x5 | ~x6 | x0 | ~x2))) & (~x6 | ((~x3 | x5 | x0 | x2) & (x1 | (x0 ? (~x5 | (~x2 & ~x3)) : (~x2 | x5)))));
  assign n4243 = (~x4 | x5 | ~x6 | x0 | ~x2) & (x2 | ((x4 | ~x5 | ~x6 | x0 | ~x3) & (x3 | ((~x5 | x6 | x0 | ~x4) & (~x0 | (x4 ? ~x6 : (~x5 | x6)))))));
  assign n4244 = n4247 & (x1 | n4246) & (~x2 | x6 | n4245);
  assign n4245 = (~x4 | x5 | ~x7 | ~x0 | x1 | ~x3) & (x0 | ((x1 | x3 | x4 | x5 | ~x7) & (~x5 | (~x1 & ~x3) | (~x4 ^ x7))));
  assign n4246 = (x0 | x2 | x3 | x4 | x5 | ~x6) & (~x3 | x6 | ((x0 | (x2 ? (x4 | x5) : (~x4 | ~x5))) & (x4 | ~x5 | ~x0 | ~x2)));
  assign n4247 = (x1 | (x0 ? (x4 ? (x5 | ~x6) : (x6 | (x3 & x5))) : (~x5 | ((x4 | ~x6) & (x3 | ~x4 | x6))))) & (x0 | x4 | ((~x1 | x5 | x6) & (x3 | ~x5 | ~x6)));
  assign z368 = x3 ? (n4252 | ~n4253) : (~n4250 | (~x5 & ~n4249));
  assign n4249 = (~x1 | x2 | x4 | ~x6 | x7) & (x6 | ((~x0 | x1 | x4 | x7) & (x0 | ~x4 | (x1 ? (x2 | ~x7) : (~x2 | x7)))));
  assign n4250 = n4251 & (~n2573 | (x0 ? (x1 | ~n1690) : (~x1 | n2176)));
  assign n4251 = (x0 | ((~x6 | ((x1 | ~x5 | (x2 & x7)) & (x5 | (~x1 & ~x2) | ~x7))) & (x6 | ~x7 | x1 | x5) & (~x1 | ((x5 | x6 | x7) & (~x2 | (x5 ? (x6 | ~x7) : x7)))))) & (x1 | x2 | ~x5 | x6 | x7) & (~x0 | ((x2 | ((~x5 | x6 | x7) & (~x1 | (x5 ? ~x6 : (x6 | ~x7))))) & (x1 | (x5 ? (x6 & (~x2 | ~x7)) : (~x6 | x7)))));
  assign n4252 = ~n620 & ((~x0 & x5 & (~x1 ^ ~x2)) | (x0 & ~x1 & x2 & n2095));
  assign n4253 = ~n4254 & n4256 & (x5 | ~n541 | n4255);
  assign n4254 = ((~x0 & ~x5 & (~x1 ^ ~x2)) | (x0 & ~x1 & x2 & x5)) & (~x6 ^ x7);
  assign n4255 = (~x6 | x7 | x1 | ~x2) & (x6 | ~x7 | ~x1 | x2);
  assign n4256 = ((x0 ? (x1 | x2) : (~x1 | ~x2)) | (~x5 ^ ~x7)) & (x0 | x1 | x2 | (~x5 ^ x7));
  assign z369 = (~x1 & (n4259 | (x0 & ~n4258))) | ~n4261 | (~x0 & x1 & ~n4260);
  assign n4258 = (~x2 | ((x3 | ~x6 | ~x7) & (~x3 | x4 | x5 | x6 | x7))) & (~x6 | ~x7 | ((x3 | (x4 & x5)) & (x2 | x4 | x5))) & (x3 | x6 | x7 | (~x4 & ~x5));
  assign n4259 = ~x3 & n616 & (n837 | ((x4 | x5) & ~n662));
  assign n4260 = (x5 | ~x6 | ~x7 | ~x2 | ~x3 | x4) & (x3 | ((x6 | x7 | x4 | x5) & (x2 | ((~x5 | ~x6 | ~x7) & (~x4 | (x6 ^ x7))))));
  assign n4261 = (~x3 | n4263) & (n620 | n4262) & (~n694 | ~n699);
  assign n4262 = (x2 | ((~x0 | ((~x3 | x4 | x5) & (~x1 | x3 | ~x4))) & (x3 | ((~x5 | (~x1 ^ x4)) & (x0 | (x1 & x4)))))) & (x0 | ~x1 | ~x2 | (x3 & (x4 | x5)));
  assign n4263 = (x1 & (x2 ^ x6)) | ((x0 | ~x1) & (x2 ^ ~x6)) | (~x4 & ~x5 & (x0 | (x2 & x6)));
  assign z370 = ~n4267 | (n597 & ~n4265) | (~x4 & ~n4266);
  assign n4265 = x3 ? (x0 ? (x1 | ((~x6 | ~x7) & (x2 | x6 | x7))) : ((~x2 | x6 | x7) & (~x1 | ((x6 | x7) & (~x2 | ~x6 | ~x7))))) : ((~x0 | x6 | ~x7 | (x1 & x2)) & (~x6 | x7 | (x0 & x1)));
  assign n4266 = (~x5 | ((x0 | ((x3 | x7) & (~x3 | ~x7 | ~x1 | ~x2))) & (x2 | x3 | x7) & (x1 | ((x3 | x7) & (~x0 | ~x3 | ~x7))))) & (~x0 | ~x3 | x5 | x7 | (x1 ^ ~x2));
  assign n4267 = (x1 & ((x2 & ~x4) | (x0 & (x2 | x7)))) | (~x3 & x7) | (x3 & ~x7) | (~x4 & (x0 | ~x7));
  assign z371 = n4269 | n4272 | n4273 | ~n4274 | (~x5 & ~n4271);
  assign n4269 = ~x4 & (n1244 | (~x5 & ~n4270));
  assign n4270 = (x0 | x1 | x2 | ~x3 | x6 | x7) & (x3 | ((x0 | ~x1 | ~x2 | x6 | ~x7) & (~x0 | ~x6 | (x1 ? (x2 | ~x7) : (~x2 | x7)))));
  assign n4271 = (x1 | ((x6 | ~x7 | x0 | x4) & (~x2 | ((x6 | x7 | x0 | ~x4) & (~x0 | ~x6 | (~x4 ^ x7)))))) & (x0 | x2 | x6 | ((x4 | ~x7) & (~x1 | ~x4 | x7)));
  assign n4272 = ~x5 & ((~x2 & ~x4 & x6 & x0 & ~x1) | (x2 & x4 & ~x6 & ~x0 & x1));
  assign n4273 = ~x4 & ((~x1 & x5) | (~x0 & (x5 | x6)));
  assign n4274 = ~x0 | ~x4 | (x1 ? (~n563 | ~n653) : ~n730);
  assign z372 = n4277 | ~n4278 | (~x3 & (n4276 | (n698 & n750)));
  assign n4276 = n873 & ((x6 & ~n868 & x0 & x2) | (~x0 & ~x2 & n757));
  assign n4277 = ~n800 & ((~n2156 & (x0 ^ ~x6)) | (~x0 & ~x6 & (n742 | n811)));
  assign n4278 = n4279 & (n912 | n1362) & (x2 | ~n1120 | ~n664);
  assign n4279 = n4280 & (~n1156 | ~n605 | (x0 ? (~x2 | ~x6) : (x2 | x6)));
  assign n4280 = x0 ? (~x5 | x6 | (x1 ? (x2 | x3) : ~x2)) : (x1 | x5 | (~x6 & (x2 | ~x3)));
  assign z373 = ~n4284 | n4288 | (x5 ? (~x0 & ~n4289) : ~n4282);
  assign n4282 = x0 ? ((~n742 | ~n1844) & (~n672 | ~n811)) : n4283;
  assign n4283 = (x1 | x3 | x4 | x6 | ~x7) & ((~x6 ^ x7) | ((~x1 | x2 | ~x3) & (~x2 | x3 | (x1 & x4))));
  assign n4284 = n4287 & ~n4286 & (~n732 | n4285 | x4 | ~x5);
  assign n4285 = x1 ? (~x2 | ~x6) : (x2 | x6);
  assign n4286 = (~x0 | (x6 ^ ~x7)) & (~n2156 | (n538 & n1838)) & (x0 | (~x6 ^ ~x7));
  assign n4287 = (x0 | ~x3 | (x1 ? (~x2 | ~x6) : (x2 | x6))) & (~x0 | x1 | x2 | ~x6);
  assign n4288 = ~x3 & ((x0 & ~x1 & x2 & ~x4 & x6) | (~x0 & x4 & (x1 ? (x2 & x6) : (~x2 & ~x6))));
  assign n4289 = (x2 | ~x3 | ~x4 | ~x6 | x7) & ((~x6 ^ x7) | ((~x1 | x2 | ~x3) & (x1 | ~x2 | x3 | x4)));
  assign z374 = ~n4295 | ~n4294 | ~n4293 | n4291 | ~n4292;
  assign n4291 = ~x7 & ((~x0 & ~x1 & ~x2 & x3 & ~x4) | (~x3 & ((x0 & ~x1 & x2 & ~x4) | (~x0 & x4 & (x1 ^ ~x2)))));
  assign n4292 = (~n738 | ~n3134) & (~n698 | ~n754);
  assign n4293 = ~x2 | (x0 ? (x1 | ~n3726) : (~x1 | ~n2527));
  assign n4294 = ~x7 | ((x0 | (x1 ^ ~x2)) & (x1 | ~x2 | ~x3) & (~x1 | x2 | x3));
  assign n4295 = (x0 | (n4296 & (x1 | ~n665 | ~n568))) & (x1 | ~n4297);
  assign n4296 = (x3 | x4 | ((~x5 | x7 | x1 | x2) & (~x1 | ~x2 | (~x5 ^ x7)))) & (x1 | x2 | ~x3 | ~x4 | (x5 ^ x7));
  assign n4297 = n916 & ((~x0 & ~x2 & n3098) | (x0 & x2 & x4 & ~n662));
  assign z375 = n4299 | n4302 | ~n4303 | (~x4 & ~n4301);
  assign n4299 = ~x2 & ((n686 & n937) | (x5 & ~n4300));
  assign n4300 = (x0 | ~x1 | x3 | ~x6 | (x4 ^ x7)) & (x1 | x6 | ((~x4 | x7 | x0 | ~x3) & (~x0 | (x3 ? (x4 | ~x7) : (~x4 | x7)))));
  assign n4301 = (~x3 | x5 | ~x6 | x0 | x1 | ~x2) & (x2 | ((~x0 | ~x3 | (x1 ? (x5 | x6) : (~x5 | ~x6))) & (x3 | ~x5 | x6 | x0 | ~x1)));
  assign n4302 = ~x0 & ((~x4 & ~x5 & x1 & ~x3) | (~x1 & x3 & (x2 ? (~x4 & x5) : (x4 & ~x5))));
  assign n4303 = (~x1 | (x0 ? (x2 | x3) : (~x3 | ~x4))) & (x2 | (x0 ? ((x3 | x4) & (x1 | ~x3 | ~x4)) : ((~x3 | x4) & (x1 | x3 | ~x4)))) & n4304 & (~x3 | ~x4 | x0 | ~x2);
  assign n4304 = n4305 & (~n1176 | ~n2112) & (~n587 | ~n1180);
  assign n4305 = ~x0 | x1 | x3 | (x2 ? x4 : (~x4 | x5));
  assign z376 = ~n4310 | (~x2 & (~n4309 | (x5 ? ~n4308 : ~n4307)));
  assign n4307 = (~x0 | ~x1 | ~x3 | x4 | ~x6 | x7) & (~x7 | ((x0 | x1 | x3 | x4 | x6) & ((~x0 ^ x3) | (x1 ? (~x4 | x6) : (x4 | ~x6)))));
  assign n4308 = (x0 | ~x1 | x3 | ~x4 | ~x6 | x7) & (x1 | ~x3 | ((x6 | x7 | x0 | ~x4) & (~x0 | (x4 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n4309 = (~x0 | ((~x1 | x3 | ~x4 | ~x5) & (x4 | x5 | x1 | ~x3))) & (x1 | x3 | x4 | ~x5) & (x0 | ((x1 | x4 | ~x5) & (~x4 | (x1 ? (x3 ^ x5) : (~x3 | x5)))));
  assign n4310 = ~n4312 & ~n4313 & ~n4314 & n4315 & (x5 | n4311);
  assign n4311 = x1 ? (x2 | ((~x4 | ~x6 | x0 | ~x3) & (~x0 | (x3 ? (x4 | x6) : (~x4 | ~x6))))) : ((~x0 | ~x2 | x3 | ~x4 | x6) & (x0 | x4 | (x2 ? (~x3 | x6) : (x3 | ~x6))));
  assign n4312 = x2 & ((~x0 & x1 & ~x3 & ~x4 & ~x5) | (~x1 & x3 & (x0 ? (x4 ^ x5) : (x4 & x5))));
  assign n4313 = ~x3 & ((~x0 & x1 & ~x2 & ~x4) | (~x1 & (x0 ? (x2 ^ x4) : (x2 & x4))));
  assign n4314 = n1701 & ((x0 & ~x1 & x2 & x3 & ~x6) | (~x0 & x1 & ~x3 & (~x2 ^ x6)));
  assign n4315 = (~x2 | ~n650 | ~n664) & (~n943 | ~n1180);
  assign z377 = ~n4318 | n4324 | (x1 ? (~x6 & ~n4323) : ~n4317);
  assign n4317 = x3 ? ((x5 | ~x6 | x0 | ~x4) & (~x0 | x6 | (~x4 ^ ~x5))) : ((x4 | ((~x5 | ~x6 | ~x0 | ~x2) & (x0 | ((~x5 | x6) & (~x2 | x5 | ~x6))))) & (~x0 | ~x4 | x5 | (x2 ^ ~x6)));
  assign n4318 = ~n4320 & n4322 & (~n2003 | n4319) & (n571 | n4321);
  assign n4319 = (x3 | x4 | ~x5 | x6 | ~x7) & (~x4 | ((~x3 | (x5 ? (~x6 | x7) : (x6 | ~x7))) & (~x6 | ~x7 | x3 | ~x5)));
  assign n4320 = ~x0 & ((~x5 & ~x6 & ~x1 & x3) | (x6 & (x1 ? (x3 ^ ~x5) : (~x3 & x5))));
  assign n4321 = (x0 | ~x2 | ~x7 | (~x1 ^ x5)) & (x2 | x5 | x7 | ~x0 | ~x1);
  assign n4322 = (~x3 | x5 | ~x6 | ~x0 | x1) & (x2 | x3 | ((~x0 | (x1 ? (~x5 | ~x6) : (x5 | x6))) & (~x5 | x6 | x0 | ~x1)));
  assign n4323 = (x0 | ~x2 | x3 | ~x4 | ~x5) & (x4 | (x0 ? (x2 | (~x3 ^ x5)) : ((~x3 | ~x5) & (~x2 | x3 | x5))));
  assign n4324 = ~x2 & ((~x0 & ~n4325) | (~x7 & n738 & ~n4326));
  assign n4325 = x5 ? (x7 | ((x1 | ~x3 | ~x4 | x6) & (~x1 | x3 | ~x6))) : ((x3 ^ ~x7) | (x1 ? (~x4 | x6) : (x4 | ~x6)));
  assign n4326 = (x5 | ~x6 | x3 | x4) & (~x5 | (x3 ? (x4 ^ x6) : (~x4 | x6)));
  assign z378 = ~n4330 | (~x1 & (x0 ? ~n4329 : ~n4328));
  assign n4328 = (~x2 | ~x4 | ~x6 | ~x7) & (x5 | ((~x2 | (x4 ^ x6)) & (~x4 | ~x6 | ~x7) & (~x3 | x4 | x6 | x7)));
  assign n4329 = (x2 | x3 | ~x4 | ~x6 | ~x7) & (x4 | x7 | (x2 ? (x3 ? (x5 | ~x6) : (~x5 | x6)) : (x6 | (x3 ^ x5))));
  assign n4330 = ~n4333 & ~n4334 & (n620 | n4331) & (~n664 | n4332);
  assign n4331 = (x4 | ((x5 | ((x0 | (x2 ? ~x1 : ~x3)) & (x2 | (x3 ? ~x1 : (~x0 & x1))))) & (x0 | x1 | ~x5 | (~x2 & ~x3)))) & (~x5 | ((x0 | ~x1 | x2 | x3) & (~x0 | x1 | (~x4 & (x2 | x3)))));
  assign n4332 = (~x2 | ~x4 | x5 | ~x6 | ~x7) & (x2 | x3 | x6 | ((x5 | x7) & (x4 | (x5 & x7))));
  assign n4333 = ~n1862 & ((x2 & (x0 ? ~x1 : (x1 & ~x3))) | (x0 & (x1 ? (~x2 & ~x3) : (x3 & ~x5))) | (~x1 & ~x3 & x5) | (~x0 & ((~x2 & x5) | (x1 & (x5 | (~x2 & x3))))));
  assign n4334 = ~n1311 & ((x2 & ((~x0 & x1 & x5) | (~x3 & ~x5 & x0 & ~x1))) | (x3 & x5 & ~x0 & x1) | (~x2 & ((~x3 & x5 & ~x0 & ~x1) | (x0 & (x1 ? (~x3 & x5) : (x3 & ~x5))))));
  assign z379 = ~n4336 | n4343 | (~x4 & (x0 | ~n4341) & (~x0 | ~n4342));
  assign n4336 = ~n4339 & ~n4340 & (n912 | n4337) & (x1 | n4338);
  assign n4337 = x7 ? ((~x0 | ((x1 | ~x2 | ~x3 | ~x4) & (~x1 | x2 | x3))) & (~x1 | x2 | (x3 ? x0 : ~x4))) : ((x1 | x2 | x3) & (x0 | ((~x1 | ~x2 | ~x3 | ~x4) & (x1 | x2 | x4))));
  assign n4338 = (~x0 | ((~x2 | x3 | x4 | x5 | ~x7) & (~x5 | x7 | x2 | ~x3))) & (x0 | ~x7 | ((~x4 | x5 | ~x2 | ~x3) & (x2 | x3 | ~x5))) & (~x5 | x7 | (x2 ? (x3 | x4) : (~x3 | ~x4)));
  assign n4339 = ~n1099 & ((~x2 & ~x5 & ~x7 & x0 & x1) | (x2 & ((~x1 & ~x5 & x7) | (~x0 & (x1 ? (x5 ^ ~x7) : (x5 & ~x7))))));
  assign n4340 = n664 & ((x2 & x5 & x7 & (x3 ^ ~x4)) | (~x5 & ((x2 & ~x3 & ~x4 & ~x7) | (~x2 & (x3 ? (x4 & ~x7) : (~x4 & x7))))));
  assign n4341 = (~x7 | ((~x1 | ~x2 | x3 | x5 | ~x6) & (x1 | (x2 ^ ~x3) | (~x5 ^ ~x6)))) & (~x1 | x7 | ((~x5 | x6 | ~x2 | ~x3) & (x2 | ((x5 | x6) & (x3 | ~x5 | ~x6)))));
  assign n4342 = (~x1 | x2 | x3 | x5 | x6 | x7) & (x1 | (~x5 ^ ~x6) | (x2 ? (~x3 | x7) : ~x7));
  assign n4343 = x4 & ((~n846 & ~n4344) | (~x1 & ~n4345));
  assign n4344 = (x2 | x3 | x7 | x0 | ~x1) & (x1 | ((x0 | x2 | ~x3 | ~x7) & (~x0 | (x2 ? (~x3 | x7) : (x3 | ~x7)))));
  assign n4345 = x0 ? ((x2 | ~x3 | x5 | x6 | ~x7) & (~x2 | x3 | ~x5 | ~x6 | x7)) : (~x3 | ~x6 | x7 | (x2 ^ x5));
  assign z380 = n4349 | ~n4352 | (x0 ? ~n4347 : (n4350 | n4351));
  assign n4347 = (~n742 | ~n1621) & (x2 | n4348);
  assign n4348 = (x1 | ~x3 | ~x4 | ~x5 | x6) & (~x1 | x4 | x5 | x7 | (~x3 ^ x6));
  assign n4349 = ~n620 & ((x2 & (x0 ? (~x1 & (x3 ^ x4)) : (x3 & (x1 | x4)))) | (~x0 & ~x2 & ~x3 & (~x1 | ~x4)));
  assign n4350 = ~n1361 & (x2 ? (~x6 & ~n918) : (x3 & n767));
  assign n4351 = ~n3891 & x1 & n2895;
  assign n4352 = ~n4354 & n4355 & (n1116 | n2290) & (n662 | n4353);
  assign n4353 = (x2 | ((~x1 | ~x4 | (~x0 ^ x3)) & (~x0 | x1 | ~x3 | (x4 & x5)))) & (x0 | ~x2 | x3 | x4 | (x1 & x5));
  assign n4354 = x7 & n2825 & ((x0 & x1 & ~x3 & ~x4) | (~x0 & x3 & (x1 ^ x4)));
  assign n4355 = (~n1546 | ~n1967) & (~n738 | n1809 | ~x4 | ~x6);
  assign z381 = ~n4357 | n4367 | (~n662 & ~n4366);
  assign n4357 = ~n4358 & ~n4360 & ~n4361 & n4362 & (x3 | n4359);
  assign n4358 = n1317 & ((x4 & ~x5 & ~x7 & ~x1 & ~x2) | (x1 & ((~x2 & ~x4 & ~x5 & ~x7) | (x2 & x7 & (x4 ^ x5)))));
  assign n4359 = x0 ? ((~x1 | x2 | x4 | x5 | x7) & (~x4 | ~x5 | ~x7 | x1 | ~x2)) : (x1 | ~x5 | (x2 ? (~x4 | x7) : (x4 | ~x7)));
  assign n4360 = x7 & ((x0 & x1 & ~x2 & ~x3 & x4) | (~x0 & ((~x1 & ~x2 & ~x3 & x4) | ((~x1 ^ ~x2) & (x3 ^ ~x4)))));
  assign n4361 = ~x1 & ~x4 & (x0 ? (~x3 ^ x7) : (x3 & ~x7));
  assign n4362 = ~n4363 & ~n4365 & (~n558 | ~n1621) & (n800 | n4364);
  assign n4363 = ~x7 & x4 & ~x3 & ~x0 & x1;
  assign n4364 = (~x0 | x1 | x2 | ~x3 | ~x4) & (~x2 | x3 | x4 | x0 | ~x1);
  assign n4365 = x0 & ~x1 & x4 & ~x7 & (x2 ^ ~x3);
  assign n4366 = x0 ? (x3 | ((~x4 | x5 | x1 | ~x2) & (~x1 | x2 | x4 | ~x5))) : (~x3 | ((x1 | x2 | ~x4 | ~x5) & (~x1 | x4 | (~x2 ^ x5))));
  assign n4367 = x7 & ((n616 & n2238 & ~n4368) | (~x2 & ~n4369));
  assign n4368 = x1 ? (~x3 | ~x5) : (x3 | x5);
  assign n4369 = (~x0 | ((x1 | x3 | ~x4 | ~x5 | ~x6) & (~x1 | ~x3 | x4 | x5 | x6))) & (x0 | x1 | x3 | x4 | x5 | ~x6);
  assign z382 = n4371 | n4376 | (x1 ? ~n4375 : ~n4374);
  assign n4371 = x7 & (x1 ? (x4 & ~n4373) : ~n4372);
  assign n4372 = x0 ? (~x2 | ((x5 | ~x6 | x3 | x4) & (~x3 | (x4 ? (~x5 | ~x6) : (x5 | x6))))) : (x2 | ((x3 | x5 | x6) & (~x5 | ~x6 | ~x3 | x4)));
  assign n4373 = (~x0 | x2 | x3 | ~x5 | x6) & (x0 | (~x3 ^ x6) | (~x2 ^ x5));
  assign n4374 = (~x0 | ((x4 | ~x5 | ~x6) & (x3 | ~x4 | x5 | x6))) & (~x4 | ((~x2 | x3 | x5 | x6) & (x2 | ((x0 | (x6 ? x3 : ~x5)) & (x3 | ~x5 | x6) & (x5 | (~x3 & ~x6)))))) & (~x2 | x4 | (~x5 & (~x3 | ~x6)));
  assign n4375 = (x4 & ((~x5 & ~x6) | (~x2 & (~x5 | ~x6)) | (~x3 & (~x5 | (~x0 & ~x2))))) | (x3 & ((x0 & (x5 | x6)) | (x6 & ((~x4 & x5) | (x2 & (~x4 | x5)))))) | (x2 & ~x4 & x5) | (x0 & (x2 | (~x4 & x5 & x6)));
  assign n4376 = ~x7 & ((n730 & n814 & n1546) | (x6 & ~n4377));
  assign n4377 = x0 ? (x2 | ((~x4 | ~x5 | x1 | x3) & (x4 | x5 | ~x1 | ~x3))) : (~x2 | ~x4 | (x1 ? (~x3 | ~x5) : (x3 | x5)));
  assign z383 = ~n4380 | ~n4384 | (x1 & (n4114 | (~x0 & ~n4379)));
  assign n4379 = ((~x3 ^ x6) | ((~x5 | x7 | x2 | ~x4) & (~x2 | (x4 ? (x5 | x7) : (~x5 | ~x7))))) & (~x6 | ((x5 | ~x7 | x2 | x4) & (~x4 | ~x5 | x7 | ~x2 | ~x3)));
  assign n4380 = n4383 & (n800 | n4382) & (~x4 | n4381);
  assign n4381 = x2 ? ((x0 | x1 | x3 | x5 | x6) & (~x5 | (~x3 ^ x6) | (x0 ^ ~x1))) : ((~x0 | x1 | x3 | x5 | ~x6) & (x0 | ((~x3 | x5 | ~x6) & (~x5 | x6 | x1 | x3))));
  assign n4382 = (x0 | x1 | x2 | ~x3 | x4 | ~x6) & (~x0 | ~x4 | ((~x3 | ~x6 | x1 | ~x2) & (~x1 | x2 | x3 | x6)));
  assign n4383 = (x3 | ((x6 | (~x2 ^ x5) | (x0 ^ ~x1)) & (x2 | ~x6 | (x0 ? (~x1 | x5) : (x1 | ~x5))))) & (x1 | ~x3 | ((x0 | ~x5 | (~x2 ^ ~x6)) & (x5 | ~x6 | ~x0 | x2)));
  assign n4384 = (x4 | n4385) & (x1 | (x2 ? n4386 : n4387));
  assign n4385 = x3 ? (x5 ? ((x0 ^ ~x1) | (~x2 ^ ~x6)) : (x6 | (x0 ? (~x1 | x2) : ~x2))) : ((~x0 | ~x1 | x2 | ~x5 | x6) & (x0 | ~x6 | ((~x2 | x5) & (~x1 | x2 | ~x5))));
  assign n4386 = (x0 | x3 | x4 | x5 | x6 | ~x7) & ((x5 ^ x7) | (~x3 ^ x6) | (~x0 ^ x4));
  assign n4387 = (~x0 | ~x3 | ~x4 | x5 | x6 | ~x7) & (x3 | (x0 ? (~x6 | (x4 ? (~x5 | x7) : (x5 | ~x7))) : (x6 | (x4 ? (x5 | x7) : ~x7))));
  assign z384 = n4389 | ~n4394 | (~n662 & ~n4393) | (n664 & ~n4392);
  assign n4389 = ~x1 & (x5 ? ~n4390 : ~n4391);
  assign n4390 = x2 ? ((~x0 | ~x3 | ~x4 | x6 | ~x7) & (x0 | x3 | (x4 ? (x6 | ~x7) : ~x6))) : ((~x4 | (x0 ? (x3 ? (~x6 | ~x7) : (x6 | x7)) : (x3 | ~x6))) & (x0 | ~x3 | x4 | (~x6 ^ x7)));
  assign n4391 = (x4 | ~x6 | x7 | ~x0 | x2 | x3) & (x6 | ((~x3 | x4 | x0 | ~x2) & (x2 | ((~x4 | x7 | x0 | ~x3) & (~x0 | x4 | (~x3 & ~x7))))));
  assign n4392 = (x3 | ((~x6 | ((x2 | (x4 ? x5 : (~x5 | ~x7))) & (x5 | ((~x4 | x7) & (~x2 | x4 | ~x7))))) & (~x2 | ~x4 | x6 | (~x5 ^ x7)))) & (x2 | ~x3 | ((x6 | ~x7 | ~x4 | x5) & (x4 | x7 | (~x5 ^ x6))));
  assign n4393 = ((x0 ^ ~x3) & (x1 | (x4 & x5))) | (x0 & ((~x1 & ~x3 & ~x4) | (x2 & x4 & ~x5))) | (x1 & ((x2 & x4 & x5) | (~x3 & ~x4 & ~x5))) | (~x3 & ((x2 & (x4 ^ x5)) | (~x1 & ~x2 & x4 & x5))) | (~x2 & ~x4 & ~x5) | (~x0 & x3 & ((~x2 & ~x4) | (~x1 & ~x5 & (~x2 | ~x4))));
  assign n4394 = ~n4397 & ~n4398 & (~n3724 | ~n4395) & (x3 | n4396);
  assign n4395 = ~x6 & x3 & ~x0 & ~x2;
  assign n4396 = (x4 | ~x6 | x7 | x0 | ~x1) & (x1 | ((x0 | ~x2 | ~x4 | ~x6 | x7) & (~x0 | ((~x6 | x7 | ~x2 | x4) & (x2 | ~x4 | x6 | ~x7)))));
  assign n4397 = ~n2176 & ((~x0 & x2 & x3 & (x1 ^ x5)) | (~x2 & x5 & (x1 ? ~x3 : x0)));
  assign n4398 = ~n4010 & (x0 ? ((x1 & ~x2 & ~x4 & ~x5) | (~x1 & x2 & (x4 | x5))) : ((x1 & x2 & x4 & x5) | (~x1 & ~x2 & ~x4 & ~x5)));
  assign z385 = ~n4405 | (~x6 & ~n4400) | (~n824 & ~n4404);
  assign n4400 = (n1130 | n4402) & (x2 | n4401) & (~x2 | ~x7 | n4403);
  assign n4401 = (x4 | x5 | ~x7 | x0 | x1 | ~x3) & (x3 | ((~x0 | x1 | (x4 ? (x5 | ~x7) : (~x5 | x7))) & (~x1 | ((~x5 | x7 | ~x0 | ~x4) & (x0 | ~x7 | (~x4 ^ ~x5))))));
  assign n4402 = (~x1 | x2 | ~x3 | x5 | ~x7) & (x1 | ((x2 | ~x3 | ~x5 | ~x7) & (~x2 | (x3 ? (~x5 | x7) : (x5 | ~x7)))));
  assign n4403 = (~x0 | x1 | ~x3 | ~x4 | x5) & (x0 | x4 | (x1 ? (~x3 ^ x5) : (~x3 | ~x5)));
  assign n4404 = x0 ? ((x1 | (x2 ? (x3 ? x4 : (~x4 | x6)) : (~x3 ^ ~x4))) & (x2 | x3 | (x4 ? ~x1 : x6))) : ((~x1 | (x2 ? (x3 | ~x4) : (~x3 | x4))) & (x1 | x2 | x3 | ~x4) & (~x2 | ((~x3 | ~x4 | x6) & (x1 | (~x3 ^ ~x4)))));
  assign n4405 = (~x1 | n4408) & (~n544 | n4406) & (x1 | n4407);
  assign n4406 = (x1 | (((~x0 ^ x4) | (x2 ? (x3 | x5) : (~x3 | ~x5))) & (x0 | x4 | (x2 ? (~x3 | ~x5) : (~x3 ^ x5))))) & (x0 | ~x1 | ((x2 | ~x4 | (~x3 ^ x5)) & (x4 | ~x5 | ~x2 | x3)));
  assign n4407 = ((x0 ^ ~x2) | ((x3 | ~x4 | ~x5 | x7) & (x5 | ~x7 | ~x3 | x4))) & (x0 | x2 | x3 | x4 | x5 | ~x7) & (~x0 | ~x2 | ~x3 | ~x4 | ~x5 | x7) & ((x0 ? (~x2 | x3) : (x2 | ~x3)) | (x4 ? (x5 | ~x7) : (~x5 | x7)));
  assign n4408 = (~x0 | x2 | x3 | x4 | x5 | ~x7) & (x0 | (((~x2 ^ ~x3) | (x4 ? (x5 | ~x7) : (~x5 | x7))) & (~x2 | x3 | x4 | x5 | ~x7) & (x2 | ~x3 | ~x4 | ~x5 | x7)));
  assign z386 = ~n4411 | n4418 | (~x2 & ~n4410) | (~n1185 & ~n4417);
  assign n4410 = (~x0 | ~x1 | ~x3 | x4 | x5 | x6) & (x1 | ((x5 | ~x6 | x3 | x4) & (x0 | ((~x5 | x6 | ~x3 | ~x4) & (x3 | x5 | ~x6)))));
  assign n4411 = ~n4413 & ~n4414 & ~n4415 & n4416 & (n1041 | n4412);
  assign n4412 = (x0 | ~x2 | ((~x5 | ~x7 | x1 | x3) & (~x1 | x5 | (~x3 ^ x7)))) & (x2 | ((~x0 | ((x5 | ~x7 | x1 | ~x3) & (~x1 | x3 | ~x5 | x7))) & (~x3 | ~x5 | ~x7 | x0 | ~x1)));
  assign n4413 = ~n846 & (((x0 ? (~x1 & x2) : (x1 & ~x2)) & (x3 ^ ~x4)) | (x0 & ~x1 & ~x2 & ~x3 & x4) | (~x0 & ((x3 & ~x4 & x1 & x2) | (~x1 & (x2 ? (~x3 & x4) : (x3 & ~x4))))));
  assign n4414 = ~n2730 & ((x0 & ~x1 & x2 & x5 & ~x7) | (~x0 & ~x2 & x7 & (x1 ^ x5)));
  assign n4415 = n616 & ((n3290 & n605) | (n3291 & n758));
  assign n4416 = (n1477 | (x0 ? (x1 | ~x2) : (~x1 | x2))) & (n850 | (~x1 ^ x3) | (~x0 ^ x2));
  assign n4417 = (x4 | x5 | x7 | ~x0 | ~x1 | x2) & (x1 | ((x0 | ~x2 | x4 | x5 | ~x7) & (~x4 | ((x5 | ~x7 | x0 | x2) & (~x0 | (x2 ? (x5 | x7) : (~x5 | ~x7)))))));
  assign n4418 = ~x7 & ((~n4419 & n724) | (~x1 & ~n4420));
  assign n4419 = (x2 | x3 | x4 | x5) & (~x2 | ~x3 | ~x4 | ~x5);
  assign n4420 = (x0 | ~x2 | ~x3 | ~x4 | ~x5 | x6) & (x2 | x3 | ((x4 | ~x5 | x6) & (x5 | ~x6 | ~x0 | ~x4)));
  assign z387 = n4423 | n4426 | ~n4427 | (~n662 & ~n4422);
  assign n4422 = (x0 | (x2 ? ((~x1 | ((~x4 | x5) & (~x3 | x4 | ~x5))) & (~x3 | ~x4 | x5) & (x1 | ((~x4 | ~x5) & (x3 | x4 | x5)))) : ((x1 | ((x4 | ~x5) & (x3 | ~x4 | x5))) & (~x1 | ~x4 | ~x5) & (x4 | (~x3 ^ x5))))) & (~x1 | x2 | x3 | ~x4 | ~x5) & (~x0 | ((x4 | x5 | x2 | x3) & (x1 | ((x2 | ~x3 | ~x4 | x5) & (x3 | x4 | ~x5) & (~x2 | (x3 ? x4 : (~x4 | x5)))))));
  assign n4423 = ~x2 & (x1 ? ~n4425 : ~n4424);
  assign n4424 = (~x6 | ((~x0 | ((~x5 | ~x7 | x3 | ~x4) & (~x3 | x4 | x5 | x7))) & (~x4 | ~x5 | x7 | x0 | x3))) & (x0 | ~x3 | ~x4 | ~x5 | x6 | x7);
  assign n4425 = (x5 | ~x6 | x7 | ~x0 | ~x3 | x4) & (x0 | x3 | x6 | ~x7 | (~x4 & ~x5));
  assign n4426 = ~n2176 & ((~x0 & (x2 ? ((x3 & x5) | (x1 & (x3 | x5))) : (~x5 & (~x1 | ~x3)))) | (~x1 & ((~x2 & ~x3 & ~x5) | (x0 & (x2 ^ (x3 & x5))))));
  assign n4427 = ~n4429 & ~n4430 & (~n1176 | ~n1163) & (~n616 | n4428);
  assign n4428 = (x1 | ~x3 | x4 | x5 | ~x6 | x7) & (~x4 | ~x7 | ((x5 | x6 | x1 | ~x3) & (~x1 | ~x5 | (~x3 ^ x6))));
  assign n4429 = ~n1465 & (x0 ? (x1 ? (~x2 & ~x3) : (x2 & x3)) : ((~x2 & x3) | (~x1 & x2 & ~x3)));
  assign n4430 = ~x0 & ((n4431 & n767) | (~x1 & n2326 & n768));
  assign n4431 = x1 & ~x4;
  assign z388 = ~n4437 | (x5 ? ~n4435 : (n4434 | (~x1 & ~n4433)));
  assign n4433 = (~x7 | ((x0 | x2 | x3 | x4 | ~x6) & (x6 | ((x3 | ~x4 | (x0 & ~x2)) & (~x0 | x4 | (~x2 ^ ~x3)))))) & (~x3 | ~x4 | ~x6 | x7 | (~x0 & x2));
  assign n4434 = n664 & ((x2 & x3 & ~x4 & x6 & ~x7) | (~x3 & (x2 ? (x4 ? (x6 & ~x7) : (~x6 & x7)) : (~x7 & (~x4 | ~x6)))));
  assign n4435 = (x3 | n4436) & (~n3895 | (x1 ? x7 : ~n549));
  assign n4436 = (~x4 | (x0 ? (x7 | (x1 ? (x2 | ~x6) : (~x2 | x6))) : (~x1 | ~x7 | (~x2 & x6)))) & (x0 | x2 | x4 | (x1 ? ~x7 : (~x6 | x7)));
  assign n4437 = (~x6 | (x7 ? n4438 : n4440)) & (n2181 | n4439) & (x6 | (x7 ? n4440 : n4438));
  assign n4438 = (x2 | ((~x0 | (x1 ? (x3 | x5) : (x4 | ~x5))) & (~x4 | ((x1 | x3 | ~x5) & (x0 | ~x1 | ~x3))))) & (x0 | ((~x4 | x5 | x1 | x3) & (~x1 | ((~x3 | x5) & (x4 | ~x5 | ~x2 | x3))))) & (x1 | ((~x3 | x4 | ~x5) & (~x2 | (x3 ^ x5))));
  assign n4439 = (x2 | ((~x4 | x5 | x0 | ~x1) & (~x0 | (x1 ? (x4 | x5) : ~x5)))) & (x1 | ((~x4 | ~x5) & (x4 | x5 | x0 | ~x2)));
  assign n4440 = (x2 | ((x4 | x5 | x1 | ~x3) & (~x0 | x3 | (x1 ? (x4 | ~x5) : (~x4 | x5))))) & (x1 | ~x2 | x3 | x4 | ~x5) & (x0 | ~x3 | ((~x1 | x4 | ~x5) & (~x4 | x5 | x1 | ~x2)));
  assign z389 = ~n4444 | (~x6 & (x1 ? ~n4443 : ~n4442));
  assign n4442 = (~x7 | (x3 ? ((x2 | x4 | x5) & (x0 | (x2 ? (~x4 | x5) : x4))) : ((x4 | x5 | x0 | ~x2) & (~x0 | (x2 ? (x4 | ~x5) : ~x4))))) & (~x5 | ((x3 | ~x4 | ~x0 | x2) & (x7 | ((x0 | ~x2 | x3 | x4) & (~x0 | ~x3 | (x2 ^ x4))))));
  assign n4443 = (x2 | ((~x4 | ((x5 | x7 | x0 | ~x3) & (~x0 | x3 | (x5 & x7)))) & (x0 | ~x3 | x4 | (~x5 & ~x7)))) & (x0 | ~x2 | ((~x5 | x7 | x3 | x4) & (~x3 | ~x4 | (~x5 ^ x7))));
  assign n4444 = ~n4446 & ~n4449 & ~n4450 & n4451 & (~x4 | n4445);
  assign n4445 = x6 ? ((~x5 | ((x1 | x2 | x7) & (x0 | ~x1 | ~x2 | ~x7))) & (x1 | ~x2 | ~x7 | (~x0 & x5))) : (x7 | ((x1 | x5) & (x0 | ~x2 | (x1 & x5))));
  assign n4446 = x6 & ((x5 & n538 & ~n4448) | (~x2 & ~n4447));
  assign n4447 = x1 ? ((~x4 | ~x7 | ~x0 | x3) & (x0 | x7 | (x3 ? (~x4 | x5) : (x4 | ~x5)))) : ((~x0 | x4 | ~x5 | (~x3 ^ ~x7)) & (~x4 | ((~x3 | x5 | ~x7) & (x0 | (x3 ? ~x7 : (x5 | x7))))));
  assign n4448 = (x0 | ~x3 | ~x4 | ~x7) & (x3 | ((~x4 | x7) & (~x0 | x4 | ~x7)));
  assign n4449 = ~n630 & ((~x0 & ((x2 & ~x4) | (x1 & ~x2 & ~x3))) | (~x4 & ((~x1 & x2 & x3) | (x0 & ~x2 & ~x3))));
  assign n4450 = ~n800 & ((~x0 & x1 & n641) | (x0 & ~x1 & x2 & n642));
  assign n4451 = (x0 | ((x4 | n4453) & (x3 | ~x7 | n4452))) & (x7 | n4452 | ~x0 | ~x3);
  assign n4452 = (~x1 | x2 | x4 | x5 | ~x6) & (x1 | ((~x2 | ~x4 | ~x5 | ~x6) & (x2 | x5 | (x4 ^ x6))));
  assign n4453 = (~x1 | ~x2 | x5 | x6 | ~x7) & (x2 | ~x5 | ((~x6 | ~x7) & (x1 | x6 | x7)));
  assign z390 = n4455 | ~n4460 | (~n800 & ~n4459) | (~n824 & ~n4458);
  assign n4455 = x7 & (x1 ? ~n4457 : (~n868 & ~n4456));
  assign n4456 = x0 ? (x2 ? (x3 | ~x6) : (~x3 | x6)) : (x2 | (~x3 ^ ~x6));
  assign n4457 = (~x0 | x2 | ~x3 | x4 | x5 | x6) & (x0 | ((~x2 | x3 | x4 | ~x5 | ~x6) & (x2 | ((~x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (x3 | ~x4 | x5 | x6)))));
  assign n4458 = x2 ? ((x0 | ((~x1 | (x6 ? ~x4 : x3)) & (~x6 | (x4 ? x3 : (x1 & ~x3))))) & (x1 | ((~x0 | ~x3 | ~x6) & (x6 | ((x3 | x4) & (~x0 | (x3 & x4))))))) : ((~x0 | ~x1 | x3 | x4 | ~x6) & (x0 | ~x3 | x6 | (x1 & ~x4)));
  assign n4459 = (x0 | ~x2 | ~x3 | x6 | (x1 & ~x4)) & (x2 | ((~x0 | ((x3 | x6) & (x1 | ~x3 | ~x6))) & (x4 | x6 | ~x1 | x3) & (~x6 | ((x1 | x3 | ~x4) & (x0 | (x3 & (~x1 | x4)))))));
  assign n4460 = (n2842 | n4463) & (~x2 | ~n598 | ~n4461) & (x2 | n4462);
  assign n4461 = x4 & x5 & (x3 ^ ~x6);
  assign n4462 = (~x4 | x5 | ~x6 | x0 | x1 | ~x3) & (x3 | ((x0 | x1 | ~x4 | x5 | x6) & (~x0 | ~x5 | ~x6 | (x1 ^ x4))));
  assign n4463 = (~x2 | (x3 ? (~x5 | x6) : (x5 | ~x6))) & (x2 | ~x3 | x5 | x6);
  assign z391 = ~n4470 | (x2 ? ~n4465 : (x4 ? ~n4469 : ~n4468));
  assign n4465 = x5 ? n4467 : (n662 | n4466);
  assign n4466 = (~x0 | x1 | ~x3 | ~x4) & (x0 | (x1 ? (~x3 | x4) : (x3 | ~x4)));
  assign n4467 = (x4 | ~x6 | ~x7 | x0 | ~x1 | ~x3) & (x1 | (x0 ? ((x6 | x7 | x3 | x4) & (~x6 | ~x7 | ~x3 | ~x4)) : (x3 | (x4 ? (x6 | x7) : (~x6 | ~x7)))));
  assign n4468 = (~x3 | (x6 ^ x7) | (x0 ? (x1 | ~x5) : (~x1 | x5))) & (x1 | x3 | ((x6 | x7 | ~x0 | x5) & (x0 | ((~x6 | ~x7) & (~x5 | x6 | x7)))));
  assign n4469 = (x0 | ~x1 | x3 | ~x5 | x6 | x7) & (x5 | ((~x0 | ((~x6 | ~x7 | x1 | ~x3) & (~x1 | x3 | x6 | x7))) & (x0 | x1 | x3 | x6 | x7)));
  assign n4470 = (~x6 | ((x7 | n4471) & (x3 | ~x7 | n4472))) & n4473 & (x6 | ((~x7 | n4471) & (~x3 | x7 | n4472)));
  assign n4471 = x0 ? ((x2 | (x1 ? (x3 ? (x4 | x5) : ~x4) : (x3 | x5))) & (x1 | x3 | (x5 ? (~x2 & x4) : ~x4))) : (x1 ? ((~x2 | x3 | x4) & (~x4 | ~x5 | x2 | ~x3)) : (~x3 | ((x2 | x4 | ~x5) & (~x4 | (~x2 & x5)))));
  assign n4472 = (x0 | ~x1 | ~x2 | x4 | ~x5) & (~x4 | ((x0 | ~x1 | x2 | ~x5) & (~x0 | x1 | (x2 ^ x5))));
  assign n4473 = n4474 & (x1 | n4475) & (~n975 | n4476);
  assign n4474 = (x0 | ~x1 | ~x2 | ~x4 | (~x3 ^ x6)) & (x4 | (x0 ? ((~x3 | ~x6 | x1 | ~x2) & (~x1 | x2 | x3 | x6)) : ((x3 | ~x6 | ~x1 | x2) & (~x3 | x6 | x1 | ~x2))));
  assign n4475 = (((x2 | ~x3 | ~x4 | ~x5) & (~x2 | x3 | x4 | x5)) | (x0 ^ ~x6)) & (x2 | (x3 ? (x4 | x5) : (~x4 | ~x5)) | (x0 ^ x6));
  assign n4476 = (x5 | ~x6 | x3 | ~x4) & (~x3 | x6 | (x4 ^ ~x5));
  assign z392 = (~x3 & (n2893 | n4479)) | ~n2896 | (~x0 & n4478);
  assign n4478 = x1 & ((x2 & (~x4 ^ x7) & (x3 | ~x5)) | (x3 & x7 & ((x4 & ~x5) | (~x2 & ~x4 & x5))));
  assign n4479 = n658 & ((~x0 & ~x2 & n2743) | (~x4 & n723 & x0 & x2));
  assign z393 = ~n4481 | n4485 | (~x6 & (~n4484 | (~x7 & ~n4483)));
  assign n4481 = x2 ? n2906 : n4482;
  assign n4482 = (~x3 & ((~x0 & ((x5 & x6) | (x1 & ~x4 & ~x6))) | (x5 & x6 & (x1 | ~x4)))) | (~x5 & ~x6) | (x3 & (~x5 | (x0 & x1))) | (x4 & ((x3 & ~x6) | (~x0 & x1 & ~x5)));
  assign n4483 = (x0 | ~x1 | x2 | x3 | x4 | ~x5) & (x1 | ((x0 | ~x2 | x3 | x4 | x5) & (~x0 | ~x3 | ~x4 | (~x2 ^ ~x5))));
  assign n4484 = (x2 | ~n1144 | ~x0 | ~x1) & (n2241 | ((x1 | x2 | ~x7) & (x0 | ((x2 | ~x7) & (~x1 | ~x2 | x7)))));
  assign n4485 = x6 & ((n923 & ~n4486) | (n650 & n691 & n1546));
  assign n4486 = x2 ? ((x0 | ~x5 | ~x7) & (x1 | ((~x5 | ~x7) & (~x0 | x5 | x7)))) : ((~x1 | ~x5 | x7) & (x0 | ((~x5 | x7) & (~x1 | x5 | ~x7))));
  assign z394 = ~n4496 | n4495 | n4493 | n4492 | n4488 | n4491;
  assign n4488 = x4 & ((x5 & ~n4489) | (n916 & ~n4490));
  assign n4489 = (x0 | ~x1 | x3 | ~x6 | ~x7) & (x1 | ((~x0 | ~x2 | x3 | (x6 ^ x7)) & (x2 | ~x3 | ((~x6 | x7) & (x0 | x6 | ~x7)))));
  assign n4490 = (~x2 | x6 | x7 | ~x0 | x1) & (x0 | ~x1 | x2 | (~x6 ^ ~x7));
  assign n4491 = ~n2091 & ((~x0 & x1 & n1449) | (~x1 & (n2095 | (x0 & n1449))));
  assign n4492 = ~n622 & ((~x0 & ~x1 & x2 & x3 & x6) | (~x3 & ~x6 & ((x1 & ~x2) | (~x0 & (x1 | ~x2)))));
  assign n4493 = ~n4494 & (x0 ? n641 : n642);
  assign n4494 = (~x1 | x2 | x3 | ~x5 | ~x7) & (x1 | ((~x3 | x5 | x7) & (~x2 | (x3 ? x7 : (x5 | ~x7)))));
  assign n4495 = ~n2954 & ((x3 & x4 & x5) | (~x2 & (x3 ? x4 : (~x4 & ~x5))));
  assign n4496 = (~x0 | n4499) & (n1471 | n4497) & (x0 | n4498);
  assign n4497 = (x4 | x5 | x7 | ~x0 | x2) & (x0 | ((~x4 | ~x5 | ~x7) & (~x2 | x4 | x5 | x7)));
  assign n4498 = (x1 | ((x2 | x3 | x4 | ~x6) & (~x2 | ~x3 | ~x4 | ~x5 | x6))) & (~x1 | ~x3 | ~x4 | x5 | x6) & ((x2 ? (x3 | ~x6) : (~x3 | x6)) | (x5 ? x4 : (~x1 & ~x4)));
  assign n4499 = (x2 | ((x4 | x6 | x1 | ~x3) & (~x1 | x3 | ~x6 | (x4 & x5)))) & (x1 | x4 | ((~x2 | x3 | ~x6) & (~x3 | x5 | x6)));
  assign z395 = ~n4505 | (x1 ? ~n4503 : (x3 ? ~n4501 : ~n4502));
  assign n4501 = (x4 | ((x0 | x6 | ~x7 | (x2 ^ x5)) & (~x6 | ((~x0 | (x2 ? (x5 | x7) : (~x5 | ~x7))) & (~x5 | x7 | x0 | ~x2))))) & (~x2 | ~x4 | (x6 ^ x7) | (~x0 ^ x5));
  assign n4502 = (x0 | ~x2 | ~x4 | ~x5 | x6 | x7) & (x2 | (x0 ? (~x5 | (x4 ? x6 : (~x6 | x7))) : (x5 | (x4 ? (~x6 | ~x7) : (~x6 ^ x7)))));
  assign n4503 = (~n2317 | ~n1231) & (x5 | n4504);
  assign n4504 = x6 ? ((x4 ^ x7) | (x0 ? (x2 | x3) : (x2 ^ ~x3))) : ((x4 | ~x7 | ~x0 | x2) & (x0 | ((~x4 | x7 | x2 | ~x3) & (~x2 | x4 | ~x7))));
  assign n4505 = ~n4507 & ~n4508 & (~n3726 | ~n924) & (x5 | n4506);
  assign n4506 = (x2 | x3 | ~x7 | x0 | ~x1) & (x1 | (x0 ? (x2 | x3 | (~x4 ^ x7)) : (~x2 | ((x4 | ~x7) & (~x3 | ~x4 | x7)))));
  assign n4507 = ~n927 & ((~x2 & ((x3 & n738) | (n664 & n985))) | (n738 & (x3 ? n985 : x2)));
  assign n4508 = (~x0 | (x1 & ~x2)) & (~x1 | x2 | (x0 & ~x3)) & (n745 | n746) & (x1 | ~x2 | ~x3);
  assign z396 = ~n4520 | n4519 | n4517 | n4515 | n4510 | n4512;
  assign n4510 = x5 & ((n537 & n814 & n534) | (~x3 & ~n4511));
  assign n4511 = (~x0 | x1 | x2 | ~x4 | ~x6 | x7) & (x6 | ((x0 | ~x1 | x2 | x4 | x7) & (x1 | ((~x4 | x7 | x0 | ~x2) & (~x0 | (x2 ? (x4 | x7) : (~x4 | ~x7)))))));
  assign n4512 = ~x5 & (x4 ? ~n4514 : ~n4513);
  assign n4513 = x1 ? (x2 | ((~x6 | ~x7 | x0 | x3) & (~x0 | ~x3 | (x6 & x7)))) : (x0 ? (x2 | (x3 ? (~x6 | ~x7) : (x6 | x7))) : (~x2 | x6 | (x3 ^ x7)));
  assign n4514 = (x0 | x1 | x2 | x3 | x6 | x7) & (~x6 | ((~x0 | ~x1 | x2 | x3 | x7) & (x0 | ~x3 | ~x7 | (~x1 ^ ~x2))));
  assign n4515 = ~x1 & ~n4516;
  assign n4516 = (x0 | x3 | x5 | x6 | ~x7) & (x2 | ((x6 | ~x7 | x3 | x5) & (~x0 | ~x5 | x7 | (x3 ^ x6))));
  assign n4517 = ~n627 & ~n4518;
  assign n4518 = (~x3 | x6 | ~x7 | ~x0 | x1 | ~x2) & (x0 | ((~x1 | ((~x6 | x7 | ~x2 | x3) & (x2 | ~x3 | x6 | ~x7))) & (x1 | x2 | x3 | ~x6 | x7)));
  assign n4519 = ~x1 & ((~x0 & x2 & x3 & x5 & ~x6) | (~x2 & ((x0 & (x3 ? (x5 & ~x6) : (~x5 & x6))) | (~x5 & ~x6 & ~x0 & x3))));
  assign n4520 = n4521 & (n918 | ((~x2 | x6 | ~x0 | x1) & (x0 | (x1 ? (~x2 ^ ~x6) : (x2 | ~x6)))));
  assign n4521 = ~n4522 & n4523 & (~n537 | ~n708 | ~n694);
  assign n4522 = ~x0 & ((x1 & (x2 ? (~x5 & ~x6) : (x5 & x6))) | (~x5 & x6 & ~x1 & x2));
  assign n4523 = ~x0 | ((~x1 | x2 | x3 | x5 | x6) & (~x5 | ~x6 | x1 | ~x2));
  assign z397 = ~n4527 | (~x1 & (x0 ? ~n4525 : ~n4526));
  assign n4525 = x2 ? ((x3 | ~x4 | x5 | ~x6 | ~x7) & (~x3 | x4 | ~x5 | x6 | x7)) : (~x4 | ((~x6 | ~x7 | ~x3 | x5) & (x6 | x7 | x3 | ~x5)));
  assign n4526 = (x5 | x6 | x7 | x2 | x3 | ~x4) & (x4 | ~x7 | ((x2 | (x3 ? (~x5 | ~x6) : (x5 | x6))) & (~x5 | ~x6 | ~x2 | x3)));
  assign n4527 = n4529 & (n620 | n4528) & (x1 ? n4533 : n4532);
  assign n4528 = (~x1 | ((x2 | x3 | (x4 ? ~x0 : ~x5)) & (x0 | (x2 ? (x3 ? (x4 | x5) : ~x4) : (x3 | x4))))) & (x2 | ((~x3 | ((x1 | x4) & (~x0 | x5 | (x1 & x4)))) & (x1 | x3 | ~x4 | (x0 & ~x5))));
  assign n4529 = (n662 | n4530) & (x3 | ~n539 | n4531);
  assign n4530 = (x1 | ((x4 | x5 | ~x2 | ~x3) & (x3 | ((~x0 | x2 | (~x4 ^ x5)) & (~x2 | ~x4 | (x0 & ~x5)))))) & (x0 | ~x1 | x2 | (x3 ? x4 : (~x4 | ~x5)));
  assign n4531 = (x0 | ~x4 | x5 | ~x6 | ~x7) & (x4 | ((~x0 | ~x5 | x6 | x7) & (x0 | (x5 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n4532 = x6 ? ((x3 | x4 | ((~x2 | x5) & (~x0 | (~x2 & x5)))) & (x2 | ~x3 | ~x4 | (x0 & ~x5))) : ((~x2 | ~x3 | ~x4) & (x0 | ~x5 | (x2 ? ~x3 : (x3 | x4))));
  assign n4533 = (x6 | ((x3 | x4 | x5 | ~x0 | x2) & (x0 | (x2 ? (x3 | x4) : (~x3 | ~x4))))) & (x0 | ~x2 | ~x3 | ~x6 | (~x4 & ~x5));
  assign z398 = n4537 | ~n4539 | ~n4540 | (~x1 & (~n4535 | ~n4536));
  assign n4535 = x4 ? (~x5 | ((~x0 | (x2 ? (x3 | x7) : (~x3 | ~x7))) & (x3 | x7 | x0 | x2))) : ((x0 | ~x2 | ~x3 | (x5 ^ x7)) & (x3 | ((x5 | ~x7 | x0 | ~x2) & (~x0 | x2 | (~x5 ^ x7)))));
  assign n4536 = (x0 | x2 | x3 | x4 | ~x7) & (~x0 | ((~x3 | x4 | x7) & (~x2 | ~x7 | (~x3 ^ ~x4))));
  assign n4537 = ~x6 & ((n664 & ~n4538) | (n814 & n534 & n691));
  assign n4538 = x2 ? (x4 | ~x5 | (~x3 ^ x7)) : (x5 | (x3 ? (~x4 | x7) : ~x7));
  assign n4539 = (~x4 | ~x7 | x0 | ~x3) & (x7 | ((x3 | ~x4 | ~x0 | x2) & (x0 | (x2 ? (x3 | ~x4) : (~x3 | x4)))));
  assign n4540 = (~x1 | n4541) & (~x6 | (~n4543 & (x1 | n4542)));
  assign n4541 = (x0 | x2 | x3 | ~x5 | x7) & (x4 | ((~x3 | ~x5 | ~x7 | x0 | ~x2) & (x5 | (x0 ^ ~x2) | (~x3 ^ x7))));
  assign n4542 = ((~x0 ^ ~x2) | ((x3 | ~x4 | x5 | x7) & (~x5 | ~x7 | ~x3 | x4))) & (~x4 | x5 | ~x7 | ~x0 | x2 | ~x3) & (x0 | ~x2 | x3 | x4 | ~x5 | x7);
  assign n4543 = ~x3 & n539 & ((x5 & ~x7 & x0 & ~x4) | (~x0 & ((~x5 & ~x7) | (~x4 & x5 & x7))));
  assign z399 = ~n4549 | (x7 ? (x0 ? ~n4548 : ~n4547) : ~n4545);
  assign n4545 = (~n924 | ~n1179) & (x1 | n4546);
  assign n4546 = (~x2 | ((x4 | x5 | x6 | ~x0 | x3) & (x0 | ~x4 | (x3 ? (x5 | ~x6) : (~x5 | x6))))) & (~x0 | x2 | x5 | ~x6 | (~x3 ^ x4));
  assign n4547 = (x6 | (x1 ? (~x3 | (x2 ? (x4 | ~x5) : (~x4 | x5))) : (x3 | (x2 ? (x4 | ~x5) : x5)))) & (x4 | ~x5 | ~x6 | (x1 ? (~x2 | x3) : (x2 | ~x3)));
  assign n4548 = (x4 | ~x5 | x6 | ~x1 | x2 | x3) & (x1 | ((x2 | x3 | ~x4 | ~x5 | x6) & (~x2 | ((x3 | ~x4 | x5 | x6) & (~x5 | ~x6 | ~x3 | x4)))));
  assign n4549 = ~n4552 & n4553 & (x2 | (n4550 & n4551));
  assign n4550 = (~x1 | ((x3 | ~x4 | x5 | ~x6) & (x0 | ~x5 | (x3 ? (~x4 | ~x6) : (x4 | x6))))) & (~x0 | x1 | ((~x5 | x6 | x3 | x4) & (~x3 | (x4 ? ~x6 : (x5 | x6)))));
  assign n4551 = (x3 | ((~x5 | x6 | x0 | ~x4) & (~x0 | (x4 ? (x5 | x6) : (~x5 | ~x6))))) & (x0 | ~x3 | ~x4 | x5 | ~x6);
  assign n4552 = ~n1323 & ((~x0 & ((~x1 & ((x4 & ~x5) | (x2 & ~x4 & x5))) | (x2 & x4 & ~x5) | (~x2 & ((x4 & x5) | (x1 & ~x4 & ~x5))))) | (~x1 & x4 & (x5 ? x0 : x2)));
  assign n4553 = ~x2 | ((~x4 | n1772 | ~x0 | x1) & (x0 | (n3629 & (~x1 | ~x4 | n1772))));
  assign z400 = n4555 | ~n4556 | n4565 | n4566 | (x2 & ~n4563);
  assign n4555 = ~n846 & (x0 ? ((~x1 & x2 & x3 & x4) | (x1 & ~x2 & ~x3 & ~x4)) : ((~x1 & ~x2 & x3 & x4) | (x2 & (x1 ? (x3 ^ x4) : (~x3 & ~x4)))));
  assign n4556 = n4558 & n4559 & ~n4561 & (x2 ? n4562 : n4557);
  assign n4557 = (~x3 | x4 | x5 | x0 | x1) & (~x4 | ~x5 | ~x0 | x3);
  assign n4558 = (~x3 | ~x4 | (x5 ? ~n750 : (~x6 | ~n1887))) & (x3 | x4 | ~x5 | x6 | ~n1887);
  assign n4559 = (~n2609 | ~n4560) & (~n975 | (~n1120 & (x3 | ~n1121)));
  assign n4560 = ~x4 & x6 & (x5 ^ x7);
  assign n4561 = ~x1 & (x0 ? ((~x2 & x3 & x5 & ~x6) | (~x5 & x6 & x2 & ~x3)) : ((~x5 & x6 & ~x2 & ~x3) | (x5 & ~x6 & x2 & x3)));
  assign n4562 = (~x0 | x1 | ~x3 | x4 | x5 | x6) & (x0 | x3 | ((~x5 | ~x6 | x1 | ~x4) & (x5 | x6 | ~x1 | x4)));
  assign n4563 = (x3 | n4564) & (~x3 | x4 | ~x6 | ~n738 | n824);
  assign n4564 = (~x0 | x1 | x4 | x5 | x6 | ~x7) & (x0 | ((~x1 | x4 | x5 | ~x6 | x7) & (~x5 | x6 | ~x7 | x1 | ~x4)));
  assign n4565 = ~n806 & ((~x2 & ~x3 & ~x6 & x0 & x1) | (~x0 & ((~x1 & ~x2 & x3 & x6) | (x2 & (x1 ? (x3 ^ x6) : (~x3 & ~x6))))));
  assign n4566 = ~n1002 & ((~x0 & x1 & ~x2 & x3 & ~x6) | (~x1 & ((~x3 & (x0 ? (x2 ^ x6) : (~x2 & ~x6))) | (x3 & x6 & ~x0 & x2))));
  assign z401 = ~n4570 | ~n4574 | (~x1 & ~n4568) | (~n620 & ~n4569);
  assign n4568 = (~x4 | ~x5 | ~x6 | x0 | ~x3) & (x3 | ((x5 | ~x6 | x0 | x4) & (~x0 | x2 | x6 | (~x4 ^ ~x5))));
  assign n4569 = (~x2 | x3 | x4 | ~x0 | x1) & ((~x4 ^ x5) | ((~x0 | ~x1 | x2 | x3) & (x0 | (x1 ^ x3))));
  assign n4570 = n4571 & (n2500 | ((x0 | ~x1 | ~x2 | ~x6) & (x6 | (x0 ? (x1 ^ ~x2) : (x1 | x2)))));
  assign n4571 = ~n4573 & (~x3 | ((~n598 | ~n4572) & (~n642 | ~n1546)));
  assign n4572 = ~x7 & ~x6 & x4 & x5;
  assign n4573 = x6 & ((~x0 & x1 & ~x2 & ~x3) | (x3 & x4 & x0 & ~x1));
  assign n4574 = ~n4576 & ~n4577 & ~n4578 & (n662 | n4575);
  assign n4575 = (x0 | ((x1 | ~x3 | ~x4 | x5) & (~x1 | ~x2 | x3 | (~x4 ^ x5)))) & (x1 | ((x2 | ~x3 | x4 | ~x5) & (~x0 | ((~x4 | x5 | x2 | x3) & (x4 | ((~x3 | ~x5) & (x2 | (~x3 & ~x5))))))));
  assign n4576 = ~x5 & ((n838 & n1021) | (n2237 & n2747 & ~n4109));
  assign n4577 = ~x6 & n664 & ((n1701 & n665) | (x2 & ~n2241));
  assign n4578 = ~n571 & ((x0 & ~x1 & x2 & ~x5 & x7) | (~x0 & ((~x1 & x2 & x5 & x7) | (x1 & ~x2 & ~x5 & ~x7))));
  assign z402 = (~x7 & ~n4580) | (~x5 & ~n4582) | (x7 & ~n4584) | (x5 & ~n4583);
  assign n4580 = (x1 | n4581) & (n2730 | ((~x2 | x5 | ~x0 | x1) & (x0 | (x1 ? (x2 | x5) : (~x2 | ~x5)))));
  assign n4581 = ((~x0 ^ x5) | ((~x3 | ~x4 | ~x6) & (~x2 | x3 | x4 | x6))) & (x2 | x3 | ((x5 | ~x6 | x0 | x4) & (~x0 | ~x5 | (x4 ^ x6))));
  assign n4582 = x4 ? (~x7 | ((x1 | x2 | x3) & (x0 | (x1 & ~x2)))) : ((~x0 | x1 | ~x7 | (~x2 ^ x3)) & (x7 | ((x0 | (~x2 & (x1 | ~x3))) & (x2 | ((~x1 | x3) & (~x0 | (~x1 & x3)))))));
  assign n4583 = (~x2 | ((x4 | ~x7 | x0 | x3) & (~x4 | x7 | ~x0 | x1))) & (~x3 | ((x4 | ~x7 | x0 | ~x1) & (~x4 | x7 | ~x0 | x1))) & (x4 | ~x7 | ((x1 | x2) & (~x0 | (x1 & (x2 | x3))))) & (x7 | ((~x1 | x2 | x3 | ~x4) & (x0 | ((x2 | x3 | ~x4) & (~x1 | (~x4 & (x2 | x3)))))));
  assign n4584 = (n1041 | n2107) & (x3 | n4585);
  assign n4585 = (x0 | ~x1 | x2 | (x4 ? (x5 | x6) : (~x5 | ~x6))) & (~x2 | ((x0 | ((x5 | ~x6 | ~x1 | x4) & (x1 | ~x4 | ~x5 | x6))) & (~x0 | x1 | ~x4 | x5 | x6)));
  assign z403 = n4588 | ~n4589 | n4594 | (x6 ? ~n4587 : ~n4593);
  assign n4587 = (~x5 | ((~x0 | ~x1 | x2 | x3 | x7) & (x0 | ((~x3 | x7) & (x1 | x3 | ~x7))))) & (~x0 | x5 | ((x1 | ((~x3 | x7) & (~x2 | x3 | ~x7))) & (x2 | (x1 ? (x3 | ~x7) : ~x3))));
  assign n4588 = ~n692 & (x0 ? (~x1 & (x2 ? (x5 ^ x6) : (~x5 & ~x6))) : ((x1 & (x2 ? x5 : (~x5 & x6))) | (x2 & x5 & x6) | (~x1 & (x2 ? (~x5 & ~x6) : x5))));
  assign n4589 = (n4590 | n4591) & (~x7 | ~n1812 | n4592);
  assign n4590 = (x2 | x4 | x5 | x6) & (~x2 | ~x4 | ~x5 | ~x6);
  assign n4591 = (~x3 | x7 | ~x0 | x1) & (x3 | ~x7 | x0 | ~x1);
  assign n4592 = (x0 | ~x1 | x4 | x5 | ~x6) & (x1 | x6 | (x0 ? (~x4 ^ ~x5) : (x4 | ~x5)));
  assign n4593 = (~x3 | x5 | x7 | x0 | x1 | ~x2) & (~x5 | (x0 ? (x1 ? (x2 | x3) : (~x3 | x7)) : ((~x1 | ((~x3 | x7) & (~x2 | x3 | ~x7))) & (x2 | (x1 ? ~x3 : (x3 | ~x7))))));
  assign n4594 = ~x2 & ((~x3 & ~n4595) | (~x7 & n1317 & ~n4596));
  assign n4595 = (x4 | ((x0 | ~x1 | x5 | x6 | x7) & (~x0 | x1 | ~x5 | (~x6 & ~x7)))) & (x0 | ~x1 | ~x4 | (x5 ? x6 : (~x6 | ~x7)));
  assign n4596 = (x1 | x6 | (x4 ^ ~x5)) & (x5 | ~x6 | ~x1 | x4);
  assign z404 = n4599 | n4602 | n4603 | ~n4605 | (n1599 & ~n4598);
  assign n4598 = (x0 | ~x2 | x3 | ~x4 | x5 | x6) & (~x0 | (x2 ? ((x3 | x4 | x6) & (~x5 | ~x6 | ~x3 | ~x4)) : (~x3 | x6 | (~x4 & ~x5))));
  assign n4599 = ~x7 & ((n1421 & ~n4601) | (~x5 & ~n4600));
  assign n4600 = x1 ? (x6 | ((x3 | ~x4 | x0 | ~x2) & (~x3 | x4 | ~x0 | x2))) : (~x6 | ((~x2 | x3 | x4) & (x2 | ~x3 | ~x4) & (~x0 | (x4 ? x2 : x3))));
  assign n4601 = (x3 | x4 | ~x6 | (~x0 & ~x2)) & (x2 | ((~x3 | ~x6) & (x0 | x4 | x6)));
  assign n4602 = n1343 & ((~x0 & x1 & ~x2 & ~x4 & x6) | (~x1 & ((~x2 & ~x4 & ~x6) | (x0 & x2 & x4 & x6))));
  assign n4603 = ~n4604 & (x1 ? (x6 ^ ~x7) : (~x6 & x7));
  assign n4604 = (x3 | (x0 ? x2 : x4)) & (x0 | x2 | (x4 ? ~x3 : ~x5));
  assign n4605 = ~n4606 & (~n1400 | n989) & (~n750 | ~n1249);
  assign n4606 = x2 & ((~x1 & x6 & (x3 ^ x4)) | (~x0 & (x1 ? (x3 & ~x6) : (x4 & x6))));
  assign z405 = ~n4616 | ~n4615 | n4614 | n4613 | n4608 | n4611;
  assign n4608 = x7 & ((x3 & ~n4609) | (~x6 & n732 & ~n4610));
  assign n4609 = (~x1 | ((x4 | x5 | x6 | ~x0 | x2) & (~x4 | ~x5 | ~x6 | x0 | ~x2))) & (~x0 | x1 | ~x6 | (x2 ? (~x4 | ~x5) : (x4 | x5)));
  assign n4610 = (x4 | ~x5 | ~x1 | x2) & (~x2 | ~x4 | x5);
  assign n4611 = ~x7 & ((n750 & n1773) | (~x1 & ~n4612));
  assign n4612 = (x0 | x2 | x4 | (x3 ? (~x5 | x6) : (x5 | ~x6))) & (~x4 | ((~x2 | x3 | x5 | ~x6) & (~x0 | ~x5 | (x2 ? (~x3 | x6) : (x3 | ~x6)))));
  assign n4613 = x0 & ~x1 & (x3 ? (x2 ? (~x4 & ~x7) : (x4 & x7)) : (~x4 & x7));
  assign n4614 = ~x0 & ((x2 & ~x3 & ~x4 & x7) | (~x2 & x4 & (~x3 ^ x7)));
  assign n4615 = (x2 | ~n1122 | ~x0 | ~x1) & (x0 | ((~x1 | x2 | ~n1144) & (~x2 | ~n2527)));
  assign n4616 = (x0 & x1) | (~n4182 & (x1 | n4617) & (~n1153 | ~n1812));
  assign n4617 = (x4 | ~x5 | x7 | x0 | x2 | x3) & (~x0 | ~x4 | x5 | (x2 ? (~x3 | x7) : (x3 | ~x7)));
  assign z406 = n4619 | n4620 | ~n4621 | n4623 | (n2127 & ~n4624);
  assign n4619 = x2 & ((x3 & ((~x0 & x5 & (x1 ^ x4)) | (x4 & ~x5 & x0 & ~x1))) | (x0 & ~x1 & ~x4 & (~x3 | x5)));
  assign n4620 = ~x5 & ((~x0 & x2 & ~x3 & x4 & ~x6) | (~x2 & ((~x3 & x4 & x6) | (x0 & x3 & ~x4 & ~x6))));
  assign n4621 = (x2 | x3 | ~x4 | ~x5) & (x0 | ((~x2 | (x3 ? (~x4 | x5) : x4)) & (~x3 | ((~x5 | n4622) & (x2 | x4 | x5)))));
  assign n4622 = x1 ? (~x4 | ~x6 | (~x2 ^ x7)) : (x4 | x6 | (x2 ^ x7));
  assign n4623 = n985 & ((~x0 & x1 & x2 & x4 & ~x6) | (~x1 & ((~x4 & x6 & ~x0 & x2) | (x0 & x4 & (x2 ^ x6)))));
  assign n4624 = (x1 | ~x2 | ((x3 | ~x4 | x6 | x7) & (~x6 | ~x7 | ~x3 | x4))) & (x2 | ((~x6 | x7 | ~x3 | x4) & (~x4 | x6 | ~x7 | ~x1 | x3)));
  assign z407 = n4627 | n4629 | n4630 | ~n4631 | (~n906 & ~n4626);
  assign n4626 = (~x4 | ~x5 | ~x6 | x0 | ~x1) & (x4 | ((~x5 | x6 | x0 | x1) & (~x0 | x5 | ~x6 | (x1 ^ ~x2))));
  assign n4627 = ~x6 & ((x4 & n3824 & n2003) | (~x2 & ~n4628));
  assign n4628 = (x0 | ~x1 | x3 | x4 | ~x5 | ~x7) & (~x0 | ~x4 | x5 | (x1 ? (x3 | x7) : (~x3 | ~x7)));
  assign n4629 = ~x1 & ((~x0 & ~x3 & (x4 ? (~x5 & ~x6) : (x5 & x6))) | (x3 & ((x0 & ~x5 & (~x4 ^ x6)) | (x4 & x5 & (~x0 | ~x6)))));
  assign n4630 = ~x6 & ((n1102 & ~n1680) | (~x3 & n1449 & n750));
  assign n4631 = ~n4632 & (~n686 | ~n2609) & (n4633 | (x4 & ~n641));
  assign n4632 = ~x0 & x1 & ((x5 & ~x6 & x3 & x4) | (~x3 & (x4 ? (~x5 & ~x6) : (x5 & x6))));
  assign n4633 = x0 ? (x3 | ~x5 | (x1 & x2)) : (~x3 | x5);
  assign z408 = ~n4637 | (x5 & (x0 ? (n670 & n4635) : ~n4636));
  assign n4635 = x7 & x6 & ~x3 & ~x4;
  assign n4636 = x1 ? (x4 ? (x6 | x7) : (~x6 | (~x2 & ~x3) | ~x7)) : (x4 ? (~x6 | ~x7) : (x6 | x7));
  assign n4637 = ~n1248 & ~n4639 & (x6 ? (x7 ? n4638 : n4640) : (x7 ? n4640 : n4638));
  assign n4638 = (~x1 | x2 | x3 | (x0 ? (~x4 | x5) : (x4 | ~x5))) & (~x0 | x1 | ~x4 | x5 | (~x2 & ~x3));
  assign n4639 = ~n1041 & ((~x2 & ~x3 & ((~x1 & ~x5) | (x0 & x1 & x5))) | (~x0 & ~x5) | (x0 & ~x1 & x5 & (x2 | x3)));
  assign n4640 = x0 ? (x4 | x5 | (x2 ? x1 : (~x1 & ~x3))) : (~x4 | ~x5);
  assign z409 = n2974 | ~n4643 | (~x2 & ~n4642);
  assign n4642 = x0 ? ((x1 | x3 | ~x4 | ~x5 | ~x7) & (~x1 | ~x3 | x4 | x5 | x7)) : (~x1 | x3 | (x4 ? (x5 | ~x7) : (~x5 | x7)));
  assign n4643 = ~n4644 & ~n4645 & (~n730 | ~n563 | n2656);
  assign n4644 = x0 & ((~x1 & ~x2 & ~x3 & ~x5 & x7) | ((~x5 ^ x7) & (~x1 ^ (~x2 & ~x3))));
  assign n4645 = ~x0 & (x1 ? (~x5 & x7 & (x2 | x3)) : (x5 & ~x7));
  assign z410 = n4648 | ~n4649 | (n563 & ~n4647);
  assign n4647 = (x0 | ~x1 | ~x4 | x6 | ~x7) & (x7 | ((x4 | ~x6 | ~x0 | x1) & (x0 | (x1 ? (~x4 ^ ~x6) : (~x4 | x6)))));
  assign n4648 = ~x2 & ((~x6 & ~x7 & ~x1 & x3) | (x1 & (x0 ? (~x3 & ~x6) : (x3 & (x6 ^ x7)))));
  assign n4649 = n4651 & (x2 | ((x4 | n4650) & (~n586 | ~n762)));
  assign n4650 = (~x3 | x5 | x6 | ~x0 | ~x1) & (x0 | x3 | ((~x6 | ~x7 | ~x1 | x5) & (x6 | x7 | x1 | ~x5)));
  assign n4651 = (x0 | (x1 ? (~x2 | (~x6 ^ x7)) : (~x6 | ~x7))) & (x1 | x6 | (x7 ? ~x0 : ~x2));
  assign z411 = (n651 & (n4653 | n4654)) | ~n4655 | (n943 & n1476);
  assign n4653 = ~x7 & (~x1 ^ ~x3);
  assign n4654 = ~x5 & ((x1 & x3 & ~x4 & ~x7) | (~x1 & ~x3 & x4 & x7));
  assign n4655 = (x0 | ~x7) & (x1 | ((x4 | ~x7 | x2 | x3) & (~x0 | ~x2 | x7)));
  assign z412 = ~n1906 | (n1132 & (x0 ? (~x1 & n838) : (x1 & n1690)));
  assign z413 = ~x0 & (n4659 | ~n4660 | (~x5 & n690 & ~n4658));
  assign n4658 = (x6 | ~x7 | x1 | x2) & (~x6 | x7 | ~x1 | ~x2);
  assign n4659 = ~x3 & ~x4 & ~x5 & (x1 ? (x2 & ~x6) : (~x2 & x6));
  assign n4660 = (x1 & x2) | (~x1 & ~x2 & ~x3 & ~x4 & ~x5);
  assign z414 = n4662 | ~n4663;
  assign n4662 = ~x4 & ((x0 & ~x1 & ~x2 & x3 & ~x5) | (~x0 & ~x3 & x5 & (x1 ^ ~x2)));
  assign n4663 = n4664 & ((x0 & (x2 | x3)) | (x1 & (~x2 | (~x3 & ~x4))) | (~x1 & x2 & x3) | (~x3 & ~x4 & ~x0 & ~x2));
  assign n4664 = ~n597 | ((~n598 | n2091) & (~x7 | ~n732 | n4285));
  assign z415 = ~n4669 | (n690 & ~n4668) | (~x4 & (~n4666 | ~n4667));
  assign n4666 = (~x0 | x1 | x2 | x3 | x5 | x6) & (x0 | ((~x1 | x2 | x3 | ~x5 | x6) & (x1 | x5 | (x2 ? (~x3 | ~x6) : (~x3 ^ x6)))));
  assign n4667 = (x0 | ~x1 | x3 | (x2 ^ x5)) & (x1 | ((x3 | ~x5 | x0 | x2) & (~x3 | (x0 ? (~x2 ^ x5) : (~x2 | ~x5)))));
  assign n4668 = (x5 | ~x6 | x7 | ~x0 | x1 | x2) & (x0 | ((x1 | x2 | x5 | x6 | ~x7) & (~x1 | ~x6 | (x2 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n4669 = (x0 | ~x2 | ((~x3 | ~x4) & (~x1 | (~x3 & ~x4)))) & (x1 | ((x3 | ~x4 | x0 | x2) & (~x0 | (x2 ? x3 : (~x3 | ~x4)))));
  assign z416 = n4677 | n4676 | n4675 | n4674 | n4671 | n4673;
  assign n4671 = ~x2 & ((~x3 & ~n4672) | (n686 & n1743));
  assign n4672 = (x0 | ~x1 | x4 | ~x5 | ~x6 | ~x7) & (x1 | ((x0 | x4 | x5 | x6 | ~x7) & (~x0 | ((~x6 | ~x7 | x4 | x5) & (x6 | x7 | ~x4 | ~x5)))));
  assign n4673 = x4 & ((~x0 & x1 & ~x3) | (~x1 & ((x0 & ((x3 & x5) | (~x2 & ~x3 & ~x5))) | (x3 & (x5 ? ~x2 : (~x0 | x2))))));
  assign n4674 = ~x5 & n1123 & ((~x1 & x3 & x6) | (~x6 & (x1 ^ (x2 & ~x3))));
  assign n4675 = ~x1 & ~x4 & ((x3 & x5) | (x0 & (x2 ? (~x3 & ~x5) : x5)));
  assign n4676 = (x0 ? (~x2 & ~x5) : (x2 & x5)) & (x1 ? (~x3 & ~x4) : (x3 & x4));
  assign n4677 = ~n906 & n2327 & n664 & ~x5 & x6;
  assign z417 = n4679 | ~n4682 | (n1120 & ~n4681);
  assign n4679 = ~x2 & ((n1489 & n686) | (x0 & ~n4680));
  assign n4680 = (x5 | ~x6 | ~x7 | x1 | ~x3 | ~x4) & (x3 | ((x1 | x4 | x5 | ~x6 | ~x7) & (~x1 | (~x4 ^ x5))));
  assign n4681 = (~x0 | x1 | x2 | ~x4 | x7) & (x0 | ~x1 | (~x4 ^ x7));
  assign n4682 = ((x0 & x1) | (x4 ? (x5 | x6) : ~x5)) & (x1 | ((~x0 | ~x2 | ~x4 | x5) & (x0 | x4 | ~x6)));
  assign z418 = ~n4686 | (n949 & ~n4685) | (~x2 & ~n4684);
  assign n4684 = (~x0 | x1 | x3 | x5 | ~x6 | ~x7) & (~x5 | ((x0 | ~x1 | ~x3 | ~x6 | x7) & (~x0 | ((~x1 | x3) & (~x6 | ~x7 | x1 | ~x3)))));
  assign n4685 = (~x4 | ~x5 | ~x7 | ~x0 | x1) & (x0 | ~x1 | x7 | (~x4 ^ ~x5));
  assign n4686 = (~x5 | ((x1 | (x6 & (~x0 | (~x2 & x7)))) & (x0 | (x6 & (~x1 | ~x2 | x7))))) & (x0 | x5 | ~x6 | (x1 & ~x7));
  assign z419 = ~n4689 | (n651 & ~n4688);
  assign n4688 = (x4 | x5 | x6 | ~x1 | ~x3) & (x1 | x3 | ~x4 | ~x7 | (~x5 ^ x6));
  assign n4689 = ~n4691 & n4692 & (~n534 | ~n1967) & (n662 | n4690);
  assign n4690 = (x2 | x3 | x4 | ~x0 | x1) & (x0 | ~x1 | (~x2 & ~x3 & ~x4));
  assign n4691 = ~x1 & (x0 ? (~x6 & (x2 | x3)) : x6);
  assign n4692 = ~x1 | x2 | x3 | (x0 ? x6 : (x4 | ~x6));
  assign z429 = ~x2 & (n4694 | ~n4696 | (~x1 & ~n4695));
  assign n4694 = ~x1 & (x0 ? ((x3 & (~x4 | (~x5 & ~x6))) | (x5 & x6 & ~x3 & x4)) : (~x3 & (x6 ? (~x4 | ~x5) : (x4 | x5))));
  assign n4695 = (~x0 | ~x4 | ((x6 | ~x7 | x3 | ~x5) & (~x3 | x5 | ~x6 | x7))) & (x0 | x3 | x4 | x5 | x6 | ~x7);
  assign n4696 = ~n664 | (x3 ? (x4 | (x5 & ~n540)) : (~x4 & (~x5 | ~n537)));
  assign z430 = ~n4698 | (~x1 & ~n4700) | (x3 & ~n4701);
  assign n4698 = ~n527 & n4699 & (~n664 | (~n1812 & ~n4020));
  assign n4699 = (~n1812 | ~n598 | ~n762) & (~n1365 | ~n650 | ~n924);
  assign n4700 = (x0 | x3 | ~x4 | (x2 ? (x5 | x6) : (~x5 | ~x6))) & (~x0 | ~x2 | ~x3 | x4 | ~x5 | x6);
  assign n4701 = x2 ? (x7 | ((x5 | ~n4702) & (x4 | ~x5 | ~n3391))) : (~x7 | ((~x4 | x5 | ~n3391) & (~x5 | ~n4702)));
  assign n4702 = ~x6 & ~x4 & ~x0 & x1;
  assign z431 = ~n4709 | (x0 ? ~n4706 : (~n4704 | ~n4708));
  assign n4704 = (~n811 | ~n1231) & (~x2 | n4705);
  assign n4705 = (~x1 | ~x3 | ~x4 | ~x5 | ~x6 | x7) & (x5 | (x1 ? (x4 | (x3 ? (x6 | ~x7) : (~x6 | x7))) : (~x4 | (x3 ? (x6 | x7) : (~x6 | ~x7)))));
  assign n4706 = x1 ? (~n563 | ~n1846) : (~n4707 & (~n4020 | ~n2503));
  assign n4707 = x2 & ((~x3 & x4 & ~x5 & ~x6 & ~x7) | (x3 & ~x4 & x5 & x6 & x7));
  assign n4708 = (~x5 | ((x1 | x2 | x3 | ~x4 | ~x6) & (~x1 | ~x3 | (x2 ? (~x4 | x6) : (x4 | ~x6))))) & (~x1 | ~x2 | x4 | x5 | (~x3 ^ ~x6));
  assign n4709 = x3 ? ((~x4 | (x0 ? (x1 | (~x2 & ~x5)) : ((x2 | x5) & (~x1 | (x2 & x5))))) & (x0 | x4 | (x1 & (~x2 | ~x5)))) : ((~x0 | x4 | (x1 ? (x2 | x5) : ~x2)) & (x0 | x1 | ~x2 | ~x4 | ~x5));
  assign z432 = (~x0 & (n4711 | (x7 & ~n4712))) | ~n4714 | (x0 & x7 & ~n4713);
  assign n4711 = ~n1323 & ((~x1 & x2 & x4 & ~x5 & x7) | (~x4 & ((x5 & ~x7 & ~x1 & ~x2) | (x1 & x7 & (x2 ^ x5)))));
  assign n4712 = (x1 | x2 | x3 | x4 | x5 | x6) & (~x4 | ~x5 | ~x6 | ~x1 | ~x2 | ~x3);
  assign n4713 = (x4 | ~x5 | x6 | ~x1 | x2 | x3) & (x1 | (x2 ? ((x3 | ~x4 | x5 | x6) & (~x5 | ~x6 | ~x3 | x4)) : (~x4 | (x3 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n4714 = n3730 & ~n4715 & n4716 & ~n4718 & (~x5 | n4717);
  assign n4715 = ~x5 & n598 & (x2 ? (x3 & ~n783) : (~x3 & n2237));
  assign n4716 = (x3 | ~x4 | x5 | ~x0 | ~x1 | x2) & (x1 | (x2 ? ((x4 | x5 | x0 | x3) & (~x0 | ~x4 | (~x3 ^ x5))) : (~x3 | ((~x4 | ~x5) & (x0 | x4 | x5)))));
  assign n4717 = x0 ? ((~x1 | x2 | x3 | x4 | ~x6) & (x1 | ~x2 | ~x3 | ~x4 | x6)) : (x1 | x2 | x3 | (x4 ^ x6));
  assign n4718 = ~n785 & ((x3 & ~x4 & x6 & n664) | (~x3 & (x4 ? (x6 ? n738 : n664) : (~x6 & n738))));
  assign z433 = ~n4725 | (x4 ? (x2 ? ~n4723 : ~n4724) : ~n4720);
  assign n4720 = (x0 | ~x2 | ~n4721) & (x2 | n4722);
  assign n4721 = (x3 ^ x6) & (x1 ? (~x5 & x7) : (x5 & ~x7));
  assign n4722 = (~x6 | ((x0 | ~x1 | x3 | ~x5 | ~x7) & (x7 | ((~x0 | x1 | (~x3 ^ ~x5)) & (x0 | ~x1 | x3 | x5))))) & (x0 | x6 | ((x1 | x3 | x5 | ~x7) & (~x1 | ~x3 | (x5 ^ x7))));
  assign n4723 = (x0 | ~x1 | ~x5 | (x3 ? (~x6 | ~x7) : (x6 | x7))) & (x1 | ((x0 | ~x3 | x5 | x6 | ~x7) & (x3 | ((~x6 | ~x7 | x0 | x5) & (~x0 | x6 | (~x5 ^ x7))))));
  assign n4724 = (x0 | ~x1 | ~x3 | ~x5 | ~x6 | x7) & (~x0 | x1 | ((x3 | ~x5 | x6 | ~x7) & (~x3 | ~x6 | (~x5 ^ x7))));
  assign n4725 = ~n4726 & ~n4727 & ~n4729 & n4730 & (x1 | n4728);
  assign n4726 = n664 & (x4 ? ((x5 & ~x6 & ~x2 & x3) | (~x5 & x6 & x2 & ~x3)) : (x2 ? (x3 ? (~x5 & x6) : (x5 & ~x6)) : (x3 ? (x5 & x6) : (~x5 & ~x6))));
  assign n4727 = ~n846 & ((x0 & ((~x2 & ~x3 & ~x4) | (~x1 & x2 & x3 & x4))) | (~x2 & ((~x1 & ~x3 & x4) | (~x0 & ((~x3 & x4) | (~x1 & x3 & ~x4))))));
  assign n4728 = (~x0 | ((~x5 | x6 | x2 | ~x3) & (~x2 | x3 | x5 | ~x6))) & (x0 | ~x2 | ~x3 | x5 | ~x6) & (x3 | ((~x2 | x4 | ~x5 | x6) & (x0 | ((~x2 | ~x5 | x6) & (x5 | ~x6 | x2 | x4)))));
  assign n4729 = ~n806 & (x0 ? ((~x1 & x2 & x3 & x6) | (x1 & ~x2 & ~x3 & ~x6)) : (~x1 & ~x2 & (x3 ^ x6)));
  assign n4730 = x0 ? ((~x1 | x2 | x3 | ~x4 | ~x5) & (x1 | ~x2 | ~x3 | x4 | x5)) : (~x3 | ~x4 | (x1 ? (~x2 | x5) : (x2 | ~x5)));
  assign z434 = n4732 | ~n4735 | (x6 ? (x7 ? ~n4740 : ~n4739) : (x7 ? ~n4739 : ~n4740));
  assign n4732 = ~x0 & (x1 ? ~n4734 : ~n4733);
  assign n4733 = (x2 | x3 | ~x5 | (x4 ? (x6 | x7) : (~x6 | ~x7))) & (x5 | ((x2 | x3 | x4 | x6 | ~x7) & (~x2 | ~x3 | (x4 ? (x6 | ~x7) : (~x6 | x7)))));
  assign n4734 = (~x2 | x3 | x4 | ~x5 | x6 | x7) & (x2 | ((~x3 | x4 | ~x5 | x6 | ~x7) & (x3 | ~x6 | (x4 ? (~x5 | x7) : (x5 | ~x7)))));
  assign n4735 = (~n738 | n4738) & (x5 | n4736) & (~x5 | n4737);
  assign n4736 = (x0 | ~x1 | ~x4 | (~x3 ^ x6)) & (x4 | (x3 ? ((x2 | ~x6 | x0 | x1) & (~x0 | x6 | (x1 & x2))) : ((x1 ^ ~x2) | (x0 ^ x6))));
  assign n4737 = ((~x3 ^ x6) | ((x0 | (x1 ? (~x2 | x4) : ~x4)) & (~x0 | x1 | x2 | x4))) & (x0 | x1 | x2 | x3 | x4 | x6) & (~x0 | ~x4 | ((~x3 | ~x6 | x1 | ~x2) & (~x1 | x2 | x3 | x6)));
  assign n4738 = (~x6 | ((x2 | ((~x5 | ~x7 | ~x3 | x4) & (x3 | ~x4 | x5 | x7))) & (~x2 | x3 | x4 | ~x5 | x7))) & (~x2 | ~x4 | ~x5 | x6 | (x3 ^ ~x7));
  assign n4739 = (x3 | ((~x2 | ~x4 | ~x5 | x0 | ~x1) & (~x0 | ((~x4 | x5 | x1 | ~x2) & (x2 | (x1 ? (~x4 ^ x5) : (~x4 | ~x5))))))) & (x0 | ~x3 | (x1 ? (x4 | x5) : ((x4 | ~x5) & (x2 | ~x4 | x5))));
  assign n4740 = x0 ? (x1 | ((~x3 | ((~x4 | x5) & (~x2 | x4 | ~x5))) & (x2 | (x3 ? ~x4 : (x4 | x5))))) : ((~x4 | ~x5 | ~x1 | ~x3) & (x3 | ((x1 | ~x4 | x5) & (x4 | (x1 ? (~x2 ^ x5) : (~x2 | ~x5))))));
  assign z435 = ~n4744 | ~n4748 | (~x5 & ~n4742) | (~n824 & ~n4743);
  assign n4742 = x0 ? ((x2 | ~x3 | x4 | x7) & (x1 | ((~x3 | ~x4 | ~x7) & (~x2 | ((~x4 | ~x7) & (x3 | x4 | x7)))))) : ((~x1 | ~x2 | x3 | x4 | ~x7) & (x2 | ((~x4 | ~x7 | x1 | x3) & (~x1 | (x3 ? (x4 | ~x7) : (~x4 | x7))))));
  assign n4743 = (~x0 | x2 | x3 | (~x1 ^ x4)) & (~x3 | x4 | x1 | ~x2) & (x0 | (~x2 & ~x3) | (x1 ^ x4));
  assign n4744 = ~n4747 & (n1041 | n4745) & (n800 | n4746);
  assign n4745 = (~x3 | x5 | ~x7 | x0 | x1 | ~x2) & (~x5 | (~x2 ^ x3) | (x0 ? (x1 | ~x7) : (~x1 | x7)));
  assign n4746 = (~x0 | ~x1 | x2 | x3 | ~x4) & (x0 | ~x3 | (x1 ? (~x2 | x4) : (x2 | ~x4)));
  assign n4747 = ~x1 & x5 & ~x7 & (x0 ? (~x2 & ~x4) : (x2 & x4));
  assign n4748 = (n783 | n4749) & (x0 | (~n4751 & (x1 | n4750)));
  assign n4749 = (x0 | ~x1 | x2 | x3 | ~x5 | ~x7) & (x1 | ((x3 | ~x5 | x7 | x0 | x2) & (~x0 | ((x5 | ~x7 | x2 | x3) & (~x2 | ~x5 | x7)))));
  assign n4750 = (x2 | x4 | ~x5 | (x3 ? (x6 | x7) : (~x6 | ~x7))) & (x5 | ((x2 | x3 | x4 | ~x6 | x7) & (~x2 | ~x4 | (x3 ? (~x6 | x7) : (x6 | ~x7)))));
  assign n4751 = n539 & ((~x3 & ~x4 & ~x5 & x6 & x7) | (~x6 & ((x3 & ~x4 & x5 & x7) | (~x3 & ~x7 & (x4 ^ ~x5)))));
  assign z436 = n4753 | n4757 | n4758 | ~n4760 | (~x1 & ~n4756);
  assign n4753 = ~x2 & (x6 ? (n690 & ~n4754) : ~n4755);
  assign n4754 = (~x5 | x7 | ~x0 | x1) & (x5 | ~x7 | x0 | ~x1);
  assign n4755 = (x3 | ((x4 | (x0 ? (x1 ? (x5 | x7) : (~x5 | ~x7)) : (x1 ? ~x5 : (x5 | ~x7)))) & (x0 | ~x4 | ((x1 | ~x5 | ~x7) & (x5 | (~x1 & x7)))))) & (x0 | x1 | ~x3 | x7 | (~x4 ^ ~x5));
  assign n4756 = (x2 | ((~x5 | x6 | ~x7 | x0 | ~x3) & (~x0 | x3 | (x5 ? (x6 | x7) : (~x6 | ~x7))))) & (x0 | ~x2 | ~x6 | (x3 ? (x5 | ~x7) : (~x5 | x7)));
  assign n4757 = x5 & (x0 ? (x1 ? (~x2 & ~x3) : (x2 & x6)) : ((x2 & x3 & ~x6) | (~x1 & (x2 ^ x6))));
  assign n4758 = ~n4759 & x6 & n616;
  assign n4759 = (~x1 | ~x3 | x4 | ~x5 | ~x7) & (x1 | ((x5 | ~x7 | x3 | ~x4) & (~x3 | x7 | (~x4 ^ x5))));
  assign n4760 = ~n4761 & ~n4762 & n4763 & (n824 | n1116 | n3068);
  assign n4761 = ~n2181 & (x2 ? (n597 & n738) : (n664 & n1701));
  assign n4762 = (x2 ^ x3) & ((x5 & x6 & ~x0 & x1) | (~x5 & ~x6 & x0 & ~x1));
  assign n4763 = ~x3 | ((x5 | x6 | ~n924) & (x7 | ~n750 | ~x5 | ~x6));
  assign z437 = ~n4766 | ~n4768 | (~n662 & ~n4765);
  assign n4765 = x0 ? (x1 | ((x4 | (x5 ? x2 : x3)) & (x2 | (x5 ? ~x3 : ~x4)))) : ((~x3 | x4 | x1 | ~x2) & (~x4 | (x1 ? (x2 ? (~x3 | ~x5) : (x3 | x5)) : (~x2 | x3))));
  assign n4766 = (~n1163 | ~n2477) & (x2 | n4767);
  assign n4767 = x0 ? (x6 | (x3 ? (x4 | x5) : ((~x4 | ~x5) & (~x1 | (~x4 & ~x5))))) : ((~x3 | (x1 ? (x5 | ~x6) : (~x4 | x6))) & (~x6 | ((x3 | x4 | x5) & (~x1 | (x4 & (x3 | ~x5))))));
  assign n4768 = (n620 | n4771) & (~n2512 | n4769) & (~x2 | n4770);
  assign n4769 = (~x5 | x6 | ~x7 | x0 | x2 | ~x3) & (~x6 | (x0 ? (~x3 | x5 | (x2 ^ ~x7)) : (x3 | ~x5 | (x2 ^ x7))));
  assign n4770 = (x1 | ((~x4 | ~x6 | x0 | ~x3) & (x3 | (x0 ? (~x6 | (~x4 & ~x5)) : (x4 | x6))))) & (x0 | ~x1 | ~x3 | x6 | (x4 & x5));
  assign n4771 = x3 ? ((x0 | ~x1 | x2 | ~x4 | ~x5) & (x1 | ((x4 | x5 | x0 | x2) & (~x0 | ~x2 | (~x4 & ~x5))))) : ((~x0 | ~x1 | x2 | x4 | x5) & (x0 | (x1 ? (~x2 | (x4 & x5)) : (x2 | ~x4))));
  assign z438 = ~n4774 | (~x0 & ((n1386 & n686) | (x5 & ~n4773)));
  assign n4773 = ((~x3 ^ x6) | ((x1 | x4 | ~x7) & (~x4 | x7 | ~x1 | ~x2))) & (x4 | ((x2 | x3 | ~x6 | ~x7) & (x1 | x7 | ((x3 | x6) & (x2 | ~x3 | ~x6)))));
  assign n4774 = ~n4775 & ~n4777 & ~n4779 & (x7 ? n4780 : n4778);
  assign n4775 = x0 & ((~x1 & ~n4776) | (n1082 & n698));
  assign n4776 = (x2 | x7 | ((x3 | ~x4 | ~x5 | ~x6) & (~x3 | x4 | x5 | x6))) & (x4 | x5 | ~x7 | ((~x3 | ~x6) & (~x2 | x3 | x6)));
  assign n4777 = ~x1 & ((x0 & ~x2 & ~x3 & ~x4 & x7) | (x4 & (x0 ? ((x3 & x7) | (x2 & ~x3 & ~x7)) : (x3 ^ x7))));
  assign n4778 = x1 ? ((~x4 | x5 | x0 | ~x3) & (x2 | ((~x4 | ~x5 | x0 | x3) & (~x0 | x4 | (~x3 ^ x5))))) : (~x2 | x4 | (x0 ? (~x3 ^ x5) : (x3 | x5)));
  assign n4779 = x1 & ((~x0 & x2 & ~x3 & ~x4 & x7) | (~x7 & ((~x3 & x4 & x0 & ~x2) | (~x0 & ~x4 & (~x2 | x3)))));
  assign n4780 = (x1 | ((x4 | x5 | x0 | ~x3) & (~x0 | ((~x3 | x4 | ~x5) & (~x4 | x5 | x2 | x3))))) & (x0 | ~x1 | ~x4 | (x3 ^ x5));
  assign z439 = ~n2516 | ~n3830 | ~n3831 | n3835 | (x6 & n3834);
  assign z440 = n3840 | n4786 | (~x1 & ~n4785) | (~x0 & ~n4783);
  assign n4783 = (x7 | n4784) & (x3 | x6 | ~x7 | ~n539 | n868);
  assign n4784 = (~x4 | ((~x1 | x2 | x3 | ~x5) & (x1 | x5 | (x2 ? (~x3 | ~x6) : (x3 | x6))))) & (~x1 | x3 | x4 | (x2 ? (~x5 | x6) : x5));
  assign n4785 = (~x7 & ((~x0 & (x2 ? (x3 & x6) : (~x3 & ~x6))) | (~x2 & ~x3 & x5 & ~x6) | (x0 & x2 & ~x5))) | (~x0 & (x5 ^ x6)) | (x6 & ((~x2 & ~x3 & ~x5) | (x0 & x5 & (~x2 | x7)))) | (x0 & ~x5 & ~x6 & (x3 | x7));
  assign n4786 = x6 & n738 & n2573 & (x3 ? (x4 & ~x7) : ~x4);
  assign z441 = n4788 | n4791 | ~n4792 | (~x0 & ~n4790);
  assign n4788 = ~x5 & ((n923 & n543 & n534) | (~x7 & ~n4789));
  assign n4789 = (x3 | ~x4 | x6 | x0 | ~x1 | ~x2) & (~x3 | ((x0 | x1 | ~x2 | x4 | ~x6) & (~x0 | x2 | (x1 ? (x4 | x6) : (~x4 | ~x6)))));
  assign n4790 = (~x6 | ((~x4 | x7 | ~x2 | x3) & (x1 | ((x3 | ~x7) & (x2 | ~x3 | x7))))) & (~x1 | x6 | ((~x4 | ~x7 | (~x2 ^ ~x3)) & (x2 | ~x3 | (x4 & x7))));
  assign n4791 = ~n692 & ((~x1 & ~x2 & x6) | (~x0 & (x1 ? (~x6 & (x2 ^ x4)) : (~x4 & x6))));
  assign n4792 = (n4010 | n4794) & (~n1132 | n3429) & (n662 | n4793);
  assign n4793 = (~x0 | (x1 ? (x2 | x3) : ~x2)) & (~x1 | x2 | x3 | x4 | x5) & (x1 | ~x2 | ~x3 | ~x4);
  assign n4794 = (x0 | ~x1 | ~x2) & (~x0 | x1 | x2 | x4);
  assign z442 = ~n4798 | (x7 & (x0 ? ~n4796 : (x1 & ~n4797)));
  assign n4796 = (~x1 | x2 | x3 | x4 | x5 | x6) & (x1 | ((~x5 | ~x6 | ~x3 | ~x4) & (~x2 | (~x3 ^ ~x6))));
  assign n4797 = (x2 | x3 | x4 | ~x5 | x6) & (~x2 | ~x4 | (x3 ^ x6));
  assign n4798 = n4800 & ~n4803 & (x7 ? n4804 : (x0 | n4799));
  assign n4799 = (x5 | ((~x4 | x6 | ~x1 | x3) & (x4 | ~x6 | x1 | ~x3))) & (x2 | (x3 ? (~x6 | (x1 & ~x4)) : (~x4 | x6))) & (x1 | x3 | x4 | x6 | (~x2 & ~x5));
  assign n4800 = ~n4802 & (n1323 | n4801) & (~n814 | ~n534 | ~n691);
  assign n4801 = x7 ? ((x0 | ~x1 | ~x2 | ~x4) & (~x0 | ((x1 | ~x2) & (~x1 | x2 | x4 | x5)))) : ((x1 | x2 | ~x4 | ~x5) & (x0 | (x4 ? x2 : x1)));
  assign n4802 = x4 & ((~x2 & ~x3 & x7 & x0 & x1) | (~x0 & ~x1 & x2 & (~x3 ^ x7)));
  assign n4803 = ~x4 & ((~x0 & x1 & x2 & (~x3 ^ x7)) | (~x2 & ((x3 & ~x7 & ~x0 & x1) | (x0 & ~x1 & (x3 ^ x7)))));
  assign n4804 = (~x3 | x4 | ~x5 | x0 | x1 | ~x2) & (x2 | x3 | ((~x0 | (x1 ? (x4 | ~x5) : (~x4 | x5))) & (x4 | x5 | x0 | ~x1)));
  assign z443 = ~n2991 | n4807 | (n2328 & n4015) | (x3 & ~n4806);
  assign n4806 = (x4 | x5 | x6 | ~x0 | ~x1 | x2) & (x1 | ~x4 | ((~x0 | (x2 ? (x5 | ~x6) : (~x5 | x6))) & (x5 | ~x6 | x0 | x2)));
  assign n4807 = x3 & ((n1546 & n1846) | (n2127 & ~n4808));
  assign n4808 = (~x1 | x2 | x4 | ~x6 | x7) & (x1 | ~x2 | ~x4 | x6 | ~x7);
  assign z444 = (x2 & ~n4810) | (~x1 & ~n4811) | (~x2 & ~n4814) | (x1 & ~n4813);
  assign n4810 = (x1 | (x3 ? (x4 | (~x0 & x5)) : (~x4 | ~x5))) & (x0 | (x1 ? (~x3 ^ ~x4) : (x3 | ~x4)));
  assign n4811 = (x6 | n4812) & (~x0 | ~n1812 | ~n678);
  assign n4812 = (~x4 | ~x5 | ~x7 | x0 | x2 | x3) & (~x3 | ((x4 | ~x5 | x7 | x0 | ~x2) & (~x0 | x5 | (x2 ? (~x4 | x7) : (x4 | ~x7)))));
  assign n4813 = x0 ? (~n665 | ~n686) : (~n4707 & (~n1172 | ~n3453));
  assign n4814 = x1 ? ((~x0 | ((x3 | ~x5 | ~x6) & (x5 | x6 | ~x3 | x4))) & (~x4 | ~x5 | x0 | ~x3) & (x3 | ((x0 | (~x5 ^ x6)) & (x4 | ~x5 | ~x6) & (~x4 | (x5 & x6))))) : ((x0 | ((~x5 | ~x6 | x3 | ~x4) & (~x3 | x5 | x6))) & (x4 | x5 | ~x0 | x3) & (~x3 | ((~x0 | (~x5 ^ x6)) & (~x4 | x5 | x6) & (x4 | (~x5 & ~x6)))));
  assign z445 = ~n4821 | (x0 ? ~n4818 : (x1 ? ~n4816 : ~n4817));
  assign n4816 = (~x5 | ((~x2 | ~x3 | x4 | ~x6 | x7) & (x2 | ((~x6 | x7 | x3 | ~x4) & (~x3 | x4 | x6 | ~x7))))) & (~x2 | x3 | x5 | (x4 ? (x6 | x7) : (~x6 | ~x7)));
  assign n4817 = (~x5 | x6 | x7 | x2 | x3 | ~x4) & (x4 | ((x2 | ~x3 | x5 | ~x6 | ~x7) & (~x2 | x6 | (x3 ? (~x5 | x7) : (x5 | ~x7)))));
  assign n4818 = (x2 | n4819) & (x1 | ~x2 | n4820);
  assign n4819 = x1 ? ((~x3 | x4 | x5 | ~x6 | x7) & (~x5 | x6 | ~x7 | x3 | ~x4)) : ((~x3 | x4 | (x5 ? (~x6 | ~x7) : (x6 | x7))) & (x3 | ~x4 | x5 | ~x6 | ~x7));
  assign n4820 = (x3 | x4 | ~x5 | x6 | ~x7) & (~x4 | ((~x3 | (x5 ? (~x6 | ~x7) : (x6 | x7))) & (~x6 | x7 | x3 | x5)));
  assign n4821 = ~n4823 & n4824 & ~n4826 & (x2 | (n4822 & n4825));
  assign n4822 = (~x3 | ((x0 | ~x1 | x4 | ~x5 | ~x6) & (x6 | ((~x0 | (x1 ? (x4 | x5) : (~x4 | ~x5))) & (~x4 | x5 | x0 | x1))))) & (x0 | x3 | ((~x1 | ~x4 | x6) & (~x5 | ~x6 | x1 | x4)));
  assign n4823 = ~n783 & ((x0 & x1 & ~x2 & ~x3 & x5) | (~x0 & ((~x3 & x5 & ~x1 & x2) | (x1 & (x2 ? (x3 & x5) : (~x3 & ~x5))))));
  assign n4824 = (x1 | ((x3 | ~x4 | ~x5 | ~x0 | x2) & (~x3 | ((~x4 | ~x5 | x0 | ~x2) & (~x0 | (x2 ? (x4 | ~x5) : (~x4 | x5))))))) & (x0 | ~x2 | x4 | ((~x3 | x5) & (~x1 | x3 | ~x5)));
  assign n4825 = (x4 | x5 | ~x0 | x3) & (x0 | ((~x4 | x5 | ~x1 | ~x3) & (x1 | (x3 ? (x4 | ~x5) : (~x4 | x5)))));
  assign n4826 = n538 & (n4827 | (~x3 & (x0 ? ~n1716 : n2237)));
  assign n4827 = x6 & ~x5 & ~x4 & x0 & x3;
  assign z446 = n4829 | ~n4833 | ~n4836 | ~n4839 | (n738 & ~n4832);
  assign n4829 = ~x0 & (x1 ? ~n4830 : ~n4831);
  assign n4830 = (x7 | ((x2 | ~x3 | x4 | ~x5 | x6) & (~x2 | x3 | x5 | (~x4 ^ x6)))) & (~x4 | ~x7 | ((~x5 | x6 | ~x2 | x3) & (x2 | ~x3 | (~x5 ^ ~x6))));
  assign n4831 = (x2 | ~x3 | x4 | ~x5 | ~x6 | ~x7) & (~x2 | (x4 ? (~x6 | ~x7) : (x6 | x7)) | (x3 ^ x5));
  assign n4832 = x3 ? (x2 ? (x6 | (x4 ? (x5 | x7) : (~x5 | ~x7))) : (~x6 | (x4 ? (x5 | ~x7) : (~x5 | x7)))) : (~x4 | ((x5 | ~x6 | x7) & (x6 | ~x7 | x2 | ~x5)));
  assign n4833 = ~n4834 & ~n4835 & (n850 | (~n720 & (x0 | n2276)));
  assign n4834 = ~n1041 & ((~x0 & x1 & ~x2 & ~x3 & x5) | (~x1 & (x0 ? (x2 ? (x3 & x5) : (~x3 & ~x5)) : (x2 & (x3 ^ x5)))));
  assign n4835 = ~n1323 & ((x2 & x4 & x5 & ~x0 & x1) | (x0 & ~x1 & (x2 ? (~x4 & ~x5) : (x4 & x5))));
  assign n4836 = (~n1205 | n4837) & (n906 | n4838);
  assign n4837 = x1 ? ((~x2 | x3 | x4 | ~x5) & (x2 | ~x3 | x5)) : (~x3 | ~x4 | (~x2 ^ x5));
  assign n4838 = (x0 | x1 | x2 | x4 | x5 | ~x6) & (~x0 | ((~x1 | x2 | x4 | x5 | ~x6) & (x1 | ((x5 | x6 | x2 | x4) & (~x5 | ~x6 | ~x2 | ~x4)))));
  assign n4839 = (x6 | n4840) & (n800 | n4841);
  assign n4840 = (x4 | (x0 ? (x2 | ~x3 | (x1 ^ ~x5)) : (x3 | (x1 ? x5 : (~x2 | ~x5))))) & (x1 | x5 | ((~x0 | ~x2 | x3 | ~x4) & (x0 | x2 | ~x3)));
  assign n4841 = (~x3 | x4 | ~x6 | x0 | ~x1 | ~x2) & (x3 | ((x0 | ~x1 | x2 | ~x4 | ~x6) & (x6 | ((~x0 | (x1 ? (x2 | ~x4) : (~x2 | x4))) & (x0 | x1 | x2 | ~x4)))));
  assign z447 = n4846 | ~n4848 | (x7 ? (~n4844 | ~n4847) : ~n4843);
  assign n4843 = ((x0 ? (x1 | ~x2) : (~x1 | x2)) | ((~x4 | ~x6) & (~x3 | x4 | x6))) & (~x3 | ((x1 | ~x6 | (x2 ^ x4)) & (x0 | ((x1 | x2 | ~x4 | x6) & (x4 | ~x6 | ~x1 | ~x2)))));
  assign n4844 = (~x5 | n4845) & (n571 | ((x2 | ~x5 | x0 | ~x1) & (~x0 | x1 | (~x2 ^ ~x5))));
  assign n4845 = (~x0 | x1 | x2 | x3 | ~x4 | ~x6) & (x0 | ((~x1 | x2 | x3 | x4 | ~x6) & (x1 | ~x2 | ~x3 | ~x4 | x6)));
  assign n4846 = ~n662 & ((~x0 & ~x1 & x2 & x3 & ~x4) | (~x3 & (x0 ? (x1 ? (~x2 & x4) : (x2 & ~x4)) : (x4 & (x1 ^ ~x2)))));
  assign n4847 = (x6 | ((x3 | x4 | ((~x1 | x2) & (x0 | (~x1 & x2)))) & (~x4 | ((x1 | x2 | ~x3) & (x0 | ~x2 | (x1 ^ x3)))))) & (x1 | x3 | x4 | ~x6 | (~x0 ^ x2));
  assign n4848 = (n783 | n4849) & (x7 | (x0 ? n4850 : n4851));
  assign n4849 = x2 ? ((x5 | ~x7 | x1 | ~x3) & (x0 | ((x5 | x7 | x1 | x3) & (~x1 | ~x5 | (x3 ^ x7))))) : ((x7 | ((x3 | ~x5 | x0 | x1) & (~x0 | (x1 ? (x3 | ~x5) : x5)))) & (x0 | ~x3 | ~x7 | (~x1 ^ x5)));
  assign n4850 = (x1 | ((~x2 | ~x3 | ~x4 | x5 | x6) & (~x5 | ~x6 | x3 | x4))) & (x2 | ((x1 | ~x3 | ~x4 | ~x5 | x6) & (x5 | ~x6 | ~x1 | x4)));
  assign n4851 = ((x2 ^ x5) | ((x4 | ~x6 | x1 | x3) & (~x4 | x6 | ~x1 | ~x3))) & (~x1 | x3 | x4 | (x2 ? (x5 | ~x6) : (~x5 | x6)));
  assign z448 = n4853 | ~n4858 | (~n662 & ~n4856) | (~x1 & ~n4857);
  assign n4853 = x5 & (x3 ? ~n4854 : ~n4855);
  assign n4854 = x6 ? (x7 | ((x0 | ~x4 | (x1 & ~x2)) & (x1 | x4 | (~x0 & ~x2)))) : (~x7 | (x0 ? (x1 | (~x2 ^ ~x4)) : (~x4 | (~x1 & x2))));
  assign n4855 = (x0 | ~x1 | x2 | ~x4 | ~x6 | x7) & (x1 | ~x2 | ((~x0 | (x4 ? (~x6 | x7) : (x6 | ~x7))) & (x6 | ~x7 | x0 | ~x4)));
  assign n4856 = (x1 | ((~x2 | (x0 ? (x3 | ~x5) : (x4 | (x3 ^ x5)))) & (~x0 | x5 | (x4 ? ~x3 : x2)))) & (~x4 | ~x5 | x0 | x3) & (~x1 | ((~x4 | ~x5 | x2 | x3) & (x0 | x5 | ((~x3 | ~x4) & (x2 | x3 | x4)))));
  assign n4857 = x4 ? (x0 ? (x2 | (x3 ? (~x5 | ~x7) : x7)) : (x5 | ((~x2 | x3 | x7) & (~x3 | ~x7)))) : ((~x0 | ~x2 | x5 | (~x3 ^ ~x7)) & (~x5 | ((x2 | x3 | ~x7) & (x0 | ((x3 | ~x7) & (x2 | ~x3 | x7))))));
  assign n4858 = ~n4859 & (x5 | (n4860 & (~n1887 | (~n2347 & ~n1308))));
  assign n4859 = n4431 & ((~x0 & (x3 ? ((x5 & ~x7) | (~x2 & ~x5 & x7)) : ((x5 & x7) | (x2 & ~x5 & ~x7)))) | (~x2 & ~x3 & ((x5 & x7) | (x0 & ~x5 & ~x7))));
  assign n4860 = (x0 | n4862) & (n1306 | n3574) & (n620 | n4861);
  assign n4861 = (~x0 | x1 | ~x2 | x3 | ~x4) & (x0 | ((~x3 | x4 | x1 | ~x2) & (~x1 | x2 | x3 | ~x4)));
  assign n4862 = (x4 | ~x6 | x7 | x1 | x3) & (~x1 | ~x2 | ~x3 | ~x4 | x6 | ~x7);
  assign z449 = ~n4868 | (x0 ? ~n4864 : (x5 ? ~n4867 : ~n4866));
  assign n4864 = x1 ? (~n563 | ~n1163) : n4865;
  assign n4865 = x4 ? ((x6 | ~x7 | ~x2 | x5) & (x2 | (x3 ? (x5 ? (~x6 | ~x7) : (x6 | x7)) : (~x5 | x7)))) : (x2 ? ((~x5 | x6 | x7) & (~x6 | ~x7 | x3 | x5)) : ((x6 | x7 | x3 | x5) & (~x7 | (x3 ? (~x5 ^ x6) : (~x5 | ~x6)))));
  assign n4866 = (x3 | ((x6 | ~x7 | ~x1 | x2) & (~x4 | ~x6 | x1 | ~x2))) & (~x4 | ((~x6 | x7 | x1 | ~x2) & (~x7 | ((x1 | x2 | ~x3 | ~x6) & (~x1 | (x2 ? (~x3 | ~x6) : x6)))))) & (x1 | ~x2 | x4 | x6 | (~x3 & x7));
  assign n4867 = (~x2 | (x1 ? (~x3 | (x4 ? (x6 | ~x7) : (~x6 | x7))) : ((~x4 | x6 | x7) & (~x6 | ~x7 | x3 | x4)))) & (x1 | x2 | ((x4 | ~x6 | x7) & (~x3 | ~x4 | x6)));
  assign n4868 = ~n4870 & ~n4871 & n4872 & (n620 | n4869);
  assign n4869 = x0 ? ((~x1 | x2 | x4 | x5) & (x1 | (x2 ? (~x4 | ~x5) : (~x3 ^ ~x4)))) : ((x4 | ((x1 | (~x2 ^ ~x5)) & (~x2 | x5 | (~x1 & x3)))) & (~x1 | x2 | ~x5 | (x3 & ~x4)));
  assign n4870 = ~n571 & ((x0 & ~x1 & x2 & n691) | (~x0 & (x1 ? (x2 ? n723 : n691) : (~x2 & n723))));
  assign n4871 = ~n1862 & (x0 ? (x1 ? (~x2 & ~x3) : (x2 & x3)) : (x1 ? (x2 ^ x3) : (~x2 & ~x3)));
  assign n4872 = (x1 | n4873) & (~n540 | n2286 | x0 | ~x1);
  assign n4873 = (~x4 | ~x6 | ~x7 | x0 | ~x2 | ~x3) & (~x0 | x2 | ((~x6 | ~x7 | x3 | ~x4) & (x6 | x7 | ~x3 | x4)));
  assign z450 = n4875 | ~n4879 | (~x0 & ~n4878);
  assign n4875 = ~x1 & (x6 ? ~n4877 : ~n4876);
  assign n4876 = x7 ? ((x0 | x4 | (x2 ? x5 : (x3 | ~x5))) & (x3 | x5 | (~x2 & (~x0 | ~x4)))) : ((~x0 | ((x2 | ~x5) & (~x4 | x5 | ~x2 | ~x3))) & (~x5 | ((x2 | ~x3 | ~x4) & (x0 | ~x2 | x3 | x4))));
  assign n4877 = (x3 | ((x0 | ~x7 | (x2 ^ x5)) & (x4 | ((~x2 | x5 | x7) & (~x0 | (x5 ^ x7)))))) & (~x4 | ((x5 | x7 | x2 | ~x3) & (~x0 | ((~x5 | x7 | ~x2 | ~x3) & (x2 | ((x5 | x7) & (~x3 | ~x5 | ~x7)))))));
  assign n4878 = x1 ? ((x2 | x3 | (x4 ? (~x5 | x7) : (x5 | ~x7))) & (~x3 | ((x5 | ~x7 | x2 | ~x4) & (~x2 | ((~x5 | ~x7) & (~x4 | x5 | x7)))))) : (~x3 | ~x4 | (x2 ? (~x5 ^ x7) : (~x5 | ~x7)));
  assign n4879 = ~n4883 & ~n4884 & (~x1 | (n4881 & (x7 | n4880)));
  assign n4880 = (x2 | x3 | x4 | (x5 ^ x6)) & (x0 | ((~x5 | ~x6 | x3 | x4) & (x6 | (x3 ? (~x4 | (x2 ^ x5)) : (x4 | x5)))));
  assign n4881 = ~n4882 & (~n2317 | ~n565) & (x0 | ~n665 | ~n1172);
  assign n4882 = ~x3 & x7 & (~x0 ^ ~x2) & (x5 ^ x6);
  assign n4883 = ~n1099 & (((x2 ^ x7) & ((~x1 & x5) | (~x0 & x1 & ~x5))) | (~x2 & ~x5 & ~x7 & (x0 ^ ~x1)));
  assign n4884 = n738 & (x2 ? (n683 | (x3 & n1156)) : (x3 & n1897));
  assign z451 = n4886 | ~n4889 | n4895 | ~n4896 | (~x0 & ~n4894);
  assign n4886 = ~x1 & (x0 ? ~n4888 : ~n4887);
  assign n4887 = x3 ? (~x5 | ((x4 | x6 | x7) & (~x2 | (x4 ? (~x6 | x7) : x6)))) : (x5 | ((~x4 | ~x6 | ~x7) & (x2 | x7 | (~x4 ^ x6))));
  assign n4888 = (x4 | ((x2 | x3 | x5 | x6 | ~x7) & (x7 | ((x5 | x6 | x2 | ~x3) & (~x2 | (x3 ? (~x5 | x6) : (x5 | ~x6))))))) & (x3 | ~x4 | x5 | ~x6 | (x2 ^ x7));
  assign n4889 = (n627 | n4893) & (~n664 | n4891) & (~n4890 | n4892);
  assign n4890 = x0 & x6;
  assign n4891 = (x3 | ((x6 | x7 | ~x4 | x5) & (~x5 | ~x6 | ~x7 | x2 | x4))) & (x2 | ~x3 | ~x5 | (x4 ? (~x6 | ~x7) : (~x6 ^ x7)));
  assign n4892 = (x2 | x3 | x4 | x7) & (x1 | ((x2 | ~x3 | ~x4 | ~x7) & (~x2 | (x3 ? (~x4 | x7) : (x4 | ~x7)))));
  assign n4893 = (~x0 | x1 | x2 | x3 | ~x6 | ~x7) & (x6 | ((~x0 | x1 | (x2 ? (x3 | x7) : (~x3 | ~x7))) & (~x2 | ~x3 | x7 | x0 | ~x1)));
  assign n4894 = (x1 | ((~x6 | ~x7 | x3 | x4) & (~x4 | x6 | ~x2 | ~x3))) & (~x6 | x7 | (x2 ? (x3 | x4) : (~x3 | ~x4))) & (~x1 | (~x3 ^ ~x4) | ((~x6 | x7) & (x2 | x6 | ~x7)));
  assign n4895 = ~n2500 & ((~x0 & ~x1 & x2 & x6 & x7) | (~x6 & ((~x0 & (~x7 | (x1 & ~x2))) | (x1 & ~x2 & ~x7) | (~x1 & ((x2 & ~x7) | (x0 & ~x2 & x7))))));
  assign n4896 = (~x0 | x1 | x2 | ~x3 | ~x6 | x7) & (~x7 | (x0 ? ((~x3 | x6 | x1 | ~x2) & (~x1 | x2 | x3 | ~x6)) : ((x1 | x2 | ~x3 | x6) & (~x1 | ~x2 | (~x3 ^ x6)))));
  assign z452 = ~n4902 | (x4 ? ~n4900 : (x0 ? ~n4899 : ~n4898));
  assign n4898 = (x1 | x2 | x3 | ~x5 | x6 | x7) & (~x6 | ((x1 | x3 | x5 | x7) & (~x1 | ~x2 | (x3 ? (x5 | x7) : (~x5 | ~x7)))));
  assign n4899 = (~x5 | ~x6 | ~x7 | x1 | ~x2 | ~x3) & (x2 | x5 | ((~x1 | (x3 ? (x6 | ~x7) : (~x6 | x7))) & (x6 | x7 | x1 | ~x3)));
  assign n4900 = x5 ? ((n620 | n3066) & (~n1546 | ~n3109)) : n4901;
  assign n4901 = ((x6 ^ x7) | ((~x0 | ~x1 | x2 | x3) & (x0 | ~x2 | (x1 ^ x3)))) & (x2 | x6 | ~x7 | (x0 ? (x1 | ~x3) : (~x1 | x3)));
  assign n4902 = ~n4904 & ~n4905 & (~n1176 | ~n2692) & (x2 | n4903);
  assign n4903 = (x1 | (x0 ? ((x3 | ~x5 | x7) & (x5 | ~x7 | ~x3 | x4)) : (x3 | ~x7 | (~x4 ^ x5)))) & (x0 | ~x1 | x4 | ~x7 | (x3 ^ x5));
  assign n4904 = ~n592 & ((~x0 & x1 & ~x2 & ~x3 & x5) | (~x1 & ((x3 & ~x5 & ~x0 & x2) | (x0 & ~x2 & (x3 ^ ~x5)))));
  assign n4905 = ~n927 & ((x0 & ((x1 & ~x2 & ~x3 & x5) | (~x1 & x2 & ~x5))) | (x3 & ((~x1 & x2 & x5) | (~x0 & (x5 ? ~x1 : ~x2)))) | (~x0 & x2 & (x5 | (x1 & ~x3))));
  assign z453 = ~n4912 | (x1 ? ~n4907 : (x2 ? ~n4910 : ~n4911));
  assign n4907 = (x2 | n4908) & (x0 | ~x2 | n4909);
  assign n4908 = (x5 | ((x0 | ~x3 | ~x4 | x6 | ~x7) & (x7 | ((~x0 | x4 | (x3 ^ x6)) & (x0 | x3 | ~x4 | ~x6))))) & (~x0 | x3 | ~x5 | ~x7 | (x4 ^ x6));
  assign n4909 = x3 ? ((~x4 | ~x5 | ~x6 | ~x7) & (x4 | x5 | x6 | x7)) : (x4 | ~x6 | (~x5 ^ x7));
  assign n4910 = x0 ? ((x3 | ~x4 | x5 | x6 | ~x7) & (~x3 | x4 | ~x5 | ~x6 | x7)) : ((x3 | x4 | x5 | x6 | x7) & (~x4 | ((~x6 | ~x7 | x3 | ~x5) & (~x3 | x6 | (~x5 ^ x7)))));
  assign n4911 = (x0 | x3 | x4 | ~x5 | x6 | x7) & (x5 | ((x6 | ~x7 | x0 | x3) & (~x3 | ((~x6 | ~x7 | x0 | x4) & (~x0 | x7 | (x4 ^ x6))))));
  assign n4912 = ~n4913 & n4914 & n4916 & (n1716 | n2671);
  assign n4913 = ~n912 & ((~x0 & x1 & ~x2 & (x3 ^ ~x4)) | (~x1 & ((~x3 & x4 & ~x0 & ~x2) | (x0 & x2 & (x3 ^ x4)))));
  assign n4914 = ~n4915 & (~n535 | ~n1546);
  assign n4915 = ~x0 & (x1 ? ((~x2 & x3 & ~x4 & ~x5) | (x4 & x5 & x2 & ~x3)) : (x3 & (x2 ? (~x4 & ~x5) : x5)));
  assign n4916 = (x4 | n4917) & (~n738 | ((~x2 | ~x3 | ~x4 | ~x5) & (x3 | (x4 ? x2 : x5))));
  assign n4917 = (x0 | x3 | ((x1 | x2 | x5 | ~x6) & (~x5 | x6 | ~x1 | ~x2))) & (~x3 | x5 | x6 | ~x0 | ~x1 | x2);
  assign z454 = ~n4919 | ~n4927 | (~n1041 & ~n4926) | (~x1 & ~n4925);
  assign n4919 = ~n4923 & ~n4924 & (n4920 | n4921) & (n620 | n4922);
  assign n4920 = (~x2 | x3 | x6 | x7) & (x2 | ~x3 | ~x6 | ~x7);
  assign n4921 = (~x0 | x1 | ~x4 | ~x5) & (x0 | ~x1 | x4 | x5);
  assign n4922 = ((x1 ^ x3) | ((~x4 | ~x5 | x0 | ~x2) & (x4 | x5 | ~x0 | x2))) & (x1 | ~x3 | (x0 ? (x2 ? (x4 | ~x5) : ~x4) : (x2 | x4))) & (~x1 | x3 | ((x2 | ~x4 | (x0 & ~x5)) & (x0 | x4 | (~x2 & ~x5))));
  assign n4923 = n1021 & ((x5 & ~x6 & ~x2 & ~x4) | (x2 & (x4 ? x6 : (~x5 & ~x6))));
  assign n4924 = (x1 ? n540 : n537) & (n1415 | (n616 & n1343));
  assign n4925 = (x5 | ((x0 | ~x2 | x3 | x6 | x7) & (~x0 | ((~x2 | x3 | ~x6 | ~x7) & (x6 | x7 | x2 | ~x3))))) & (x0 | x2 | ~x5 | (x3 ? (~x6 | ~x7) : (x6 | x7)));
  assign n4926 = ((x5 ^ x7) | ((x0 | x2 | (x1 ^ x3)) & (~x2 | x3 | ~x0 | x1))) & (x3 | ((x0 | x1 | ~x2 | x5 | ~x7) & (~x0 | x2 | (x1 ? (x5 | ~x7) : (~x5 | x7))))) & (x0 | ~x2 | ~x3 | (x1 ? (x5 | ~x7) : x7));
  assign n4927 = x0 | ((~n565 | ~n1602) & n4928 & (x2 | n4929));
  assign n4928 = x1 ? ((x2 | x3 | x4 | x5 | x6) & (~x2 | ((x3 | ~x4 | ~x6) & (~x5 | x6 | ~x3 | x4)))) : ((~x2 | x3 | x4 | ~x5 | x6) & (~x4 | x5 | ~x6 | x2 | ~x3));
  assign n4929 = (~x1 | x3 | x4 | ~x5 | x6 | x7) & ((x3 ? (x6 | x7) : (~x6 | ~x7)) | (x1 ? (~x4 | ~x5) : (x4 | x5)));
  assign z455 = ~n4936 | (x0 ? ~n4933 : (x6 ? ~n4931 : ~n4932));
  assign n4931 = x2 ? ((x4 | x5 | x7 | ~x1 | x3) & (~x4 | ~x5 | ~x7 | x1 | ~x3)) : (x7 ? (x1 ? (x3 ? (~x4 | x5) : ~x5) : (x3 ? (x4 | ~x5) : (~x4 | x5))) : (x1 ? (x4 | ~x5) : (~x3 | (~x4 ^ ~x5))));
  assign n4932 = (~x4 | ((x3 | (x2 ^ x7) | (x1 ^ x5)) & (x1 | ~x3 | ~x5 | (x2 ^ ~x7)))) & (~x2 | x4 | ((x5 | x7 | x1 | ~x3) & (~x1 | (x3 ? (~x5 | x7) : (x5 | ~x7)))));
  assign n4933 = (x2 | n4934) & (x1 | ~x2 | n4935);
  assign n4934 = (~x5 | ~x6 | ~x7 | x1 | ~x3 | ~x4) & ((x4 ? (~x6 | x7) : (x6 ^ x7)) | (x1 ? (x3 | ~x5) : x5));
  assign n4935 = (x3 | x4 | ~x5 | ~x6 | x7) & (x6 | ((x3 | x4 | ~x5 | ~x7) & (~x3 | x5 | (~x4 ^ x7))));
  assign n4936 = n4937 & ~n4939 & ~n4940 & ~n4941 & (x0 | n4942);
  assign n4937 = (n927 | n4938) & (~n650 | ~n691 | ~n694);
  assign n4938 = x0 ? ((x1 | ~x2 | ~x3 | ~x5) & (~x1 | x2 | x3 | x5)) : ((x1 | x2 | x3 | ~x5) & (~x3 | x5 | ~x1 | ~x2));
  assign n4939 = ~n824 & ((x0 & ~x1 & x2 & ~x3 & x4) | (~x0 & ((x1 & ~x2 & x3 & x4) | (~x3 & ~x4 & ~x1 & x2))));
  assign n4940 = ~n1241 & ((x0 & ~x1 & x2 & n1156) | (~x0 & (x1 ? (x2 & n2205) : (~x2 & n1156))));
  assign n4941 = ~n592 & ((x0 & ~x1 & ~x2 & x5) | (~x0 & ~x5 & (x1 ? (~x2 & ~x3) : (x2 & x3))));
  assign n4942 = (~x2 | ~x3 | x4 | ~x5 | ~x7) & ((x2 ? (x3 | ~x4) : (~x3 | x4)) | (x1 ? (x5 | ~x7) : (~x5 | x7)));
  assign z456 = ~n4949 | (x2 ? ~n4946 : (x3 ? ~n4945 : ~n4944));
  assign n4944 = x4 ? ((x7 | ((x0 | (x1 ? (x5 | ~x6) : (~x5 | x6))) & (~x5 | ~x6 | ~x0 | x1))) & (~x0 | x6 | ~x7 | (x1 & ~x5))) : ((x5 | ~x6 | x7 | ~x0 | ~x1) & (x0 | ((~x1 | x6 | (x5 ^ x7)) & (~x5 | ~x6 | x7))));
  assign n4945 = (x0 | ~x1 | ~x4 | ~x5 | ~x6 | x7) & (~x7 | ((x0 | ~x1 | (x4 ? (x5 | ~x6) : (~x5 | x6))) & (x1 | (~x5 ^ ~x6) | (x0 ^ x4))));
  assign n4946 = ~n4948 & (~x4 | n4947) & (x4 | ~x5 | ~n544 | ~n958);
  assign n4947 = (~x5 | x6 | x7 | ~x0 | x1 | ~x3) & (x0 | ((~x1 | ~x3 | x5 | x6 | x7) & (~x6 | (~x3 ^ x7) | (x1 ^ x5))));
  assign n4948 = ~n692 & ((~x0 & x1 & ~x4 & x5 & ~x6) | (~x1 & ~x5 & (x0 ? (x4 ^ x6) : (~x4 & ~x6))));
  assign n4949 = ~n4951 & n4952 & (x3 | n4950);
  assign n4950 = (~x2 | ((x0 | ~x1 | x5 | (~x4 & ~x6)) & (x1 | ~x4 | ~x5 | (~x0 & x6)))) & (x1 | x2 | ((~x4 | x5 | ~x6) & (~x0 | ((x5 | ~x6) & (x4 | ~x5 | x6)))));
  assign n4951 = ~n846 & ((~x0 & x3 & (x1 ^ x4)) | (~x3 & ((x1 & ~x2 & x4) | (x0 & (x1 ? ~x2 : (x2 & ~x4))))));
  assign n4952 = ~n4953 & (~n650 | ~n1120 | ~n534) & (~n3291 | ~n1743);
  assign n4953 = ~x1 & ((~x4 & x5 & ~x6 & ~x0 & ~x3) | (x3 & ((~x5 & x6 & ~x0 & ~x4) | (x0 & (x4 ? (~x5 & x6) : (x5 & ~x6))))));
  assign z457 = ~n4968 | ~n4964 | n4962 | n4960 | n4955 | n4958;
  assign n4955 = ~x1 & ((~x0 & ~n4956) | (~x5 & n610 & ~n4957));
  assign n4956 = (x3 | ((x2 | x4 | ~x5 | x6 | x7) & (~x2 | ~x6 | ~x7 | (~x4 ^ x5)))) & (x2 | ~x3 | ~x4 | x7 | (~x5 ^ ~x6));
  assign n4957 = (x6 | ~x7 | x2 | ~x4) & (~x2 | x4 | (~x6 ^ ~x7));
  assign n4958 = ~n620 & ~n4959;
  assign n4959 = x1 ? ((x3 | ~x4 | ~x5 | ~x0 | x2) & (x0 | x4 | (x2 ? ~x5 : (x3 | x5)))) : ((x4 | x5 | x0 | ~x2) & (~x4 | ((x3 | ~x5 | x0 | x2) & (~x0 | x5 | (~x2 & ~x3)))));
  assign n4960 = ~n4961 & x1 & x4;
  assign n4961 = (x5 | ~x6 | x7 | ~x0 | x2 | x3) & (x0 | ((x2 | x3 | x5 | x6 | x7) & (~x2 | ~x3 | ~x7 | (~x5 ^ ~x6))));
  assign n4962 = x6 & ~n4963;
  assign n4963 = (x2 | (~x0 ^ x4) | (x1 ? (x3 | ~x5) : x5)) & (x1 | ~x2 | ~x5 | (x0 ? (x3 | x4) : ~x4));
  assign n4964 = n4965 & (~n1887 | ((~x4 | ~x5 | ~x6 | ~x7) & (x4 | x7 | (~x5 ^ ~x6))));
  assign n4965 = (x0 | n4967) & (n4966 | (x4 ? (~x5 | ~x7) : (x5 | x7)));
  assign n4966 = (~x0 | x1 | ~x2 | ~x3 | x6) & (x0 | ~x1 | ~x6 | (~x2 ^ x3));
  assign n4967 = (~x5 | ~x6 | ~x7 | x1 | x2 | x4) & (x6 | (~x1 ^ ~x5) | (x2 ? (~x4 | x7) : (x4 | ~x7)));
  assign n4968 = (n1215 | n4971) & (x6 | n4969) & (n2348 | n4970);
  assign n4969 = x0 ? (x2 | ((~x1 | x4 | x5) & (~x4 | ~x5 | x1 | x3))) : (x1 | x4 | ~x5 | (~x2 & ~x3));
  assign n4970 = (~x4 | x6 | x2 | ~x3) & (~x2 | (x3 ? (x4 | ~x6) : (~x4 | x6)));
  assign n4971 = x0 ? (x4 | (x1 ? (x2 | x3) : (~x2 | ~x3))) : (~x4 | (x1 ? x2 : (~x2 | ~x3)));
  assign z458 = ~n4975 | ~n4979 | (x0 & ~n4973);
  assign n4973 = (~x1 | x2 | x3 | ~x7 | n912) & (x1 | ((~x3 | n4974) & (x2 | x3 | x7 | n912)));
  assign n4974 = (x2 | x4 | x5 | ~x6 | x7) & (~x2 | ~x4 | ~x5 | x6 | ~x7);
  assign n4975 = ~n4977 & ~n4978 & (~n3726 | ~n750) & (n846 | n4976);
  assign n4976 = x1 ? (x2 | x7 | ((x3 | x4) & (x0 | (x3 & x4)))) : ((~x0 | (x2 ? (~x3 | x7) : ~x7)) & (~x7 | ((x2 | ~x3 | ~x4) & (x3 | x4 | x0 | ~x2))));
  assign n4977 = x2 & ((~x0 & x1 & (x3 ? (x5 & x7) : (~x5 & ~x7))) | (~x1 & ((~x3 & x5 & ~x7) | (~x5 & x7 & (x0 | x3)))));
  assign n4978 = ~x2 & ((x0 & ~x1 & x3 & x5 & ~x7) | (~x0 & ~x3 & x7 & (x1 ^ x5)));
  assign n4979 = (x0 & (x7 | n4980)) | (~n4982 & ~n4983 & (x7 | (n4980 & n4981)));
  assign n4980 = (~x3 | x4 | ~x5 | x0 | x1 | ~x2) & (x5 | ((x0 | x1 | x2 | x3 | ~x4) & (~x1 | ((~x3 | x4 | x0 | ~x2) & (~x0 | x2 | (~x3 ^ x4))))));
  assign n4981 = (x1 | x2 | x3 | (x4 ? (~x5 | x6) : (x5 | ~x6))) & (~x3 | ((~x4 | ~x5 | ~x6 | x1 | ~x2) & (~x1 | x6 | (x2 ? (x4 | ~x5) : (~x4 | x5)))));
  assign n4982 = ~n912 & ((~x1 & ~x2 & x3 & ~x7) | (x1 & (x2 ? (x3 ? (x4 & ~x7) : (~x4 & x7)) : (x3 & x7))));
  assign n4983 = n1599 & ((n665 & n872) | (n1812 & n757));
  assign z459 = ~n4989 | (x7 ? ~n4985 : (n4988 | (~x1 & ~n4987)));
  assign n4985 = (x1 | n4986) & (~n1365 | ~n923 | ~n924);
  assign n4986 = (~x2 | ((~x4 | x5 | ~x6 | x0 | x3) & (~x0 | x6 | (x3 ? (~x4 | x5) : (x4 | ~x5))))) & (x0 | x2 | ~x3 | x4 | (x5 ^ x6));
  assign n4987 = x0 ? (~x6 | ((~x2 | x3 | ~x4 | ~x5) & (x4 | x5 | x2 | ~x3))) : (x6 | ((~x4 | x5 | ~x2 | ~x3) & (x3 | ((x4 | ~x5) & (x2 | ~x4 | x5)))));
  assign n4988 = n758 & ((~x4 & ~x5 & ~x6 & x0 & ~x2) | (~x0 & (x2 ? (~x4 & (x5 ^ ~x6)) : (x4 & (x5 ^ x6)))));
  assign n4989 = ~n4991 & ~n4992 & ~n4993 & n4994 & (x1 | n4990);
  assign n4990 = (~x2 | ((x4 | ((~x6 | ~x7 | x0 | x3) & (~x0 | x6 | (~x3 ^ ~x7)))) & (x0 | ~x3 | ~x4 | (~x6 ^ x7)))) & (x0 | x2 | ((~x6 | x7 | ~x3 | x4) & (x3 | (x4 ? (~x6 | x7) : (x6 | ~x7)))));
  assign n4991 = x0 & ((~x4 & x6 & ~x2 & ~x3) | (~x1 & (x2 ? (x4 & (~x3 ^ x6)) : (~x3 & x6))));
  assign n4992 = ~n662 & ((x2 & ~x3 & ~x4 & ~x0 & x1) | (x0 & ~x2 & x4 & (x1 ^ x3)));
  assign n4993 = ~x0 & (x1 ? ((x4 & ~x6 & x2 & ~x3) | (~x2 & x3 & ~x4 & x6)) : (x3 & (x2 ? (~x4 & ~x6) : (x4 & x6))));
  assign n4994 = x2 ? ((x7 | n4995) & (~x3 | x6 | ~x7 | ~n664)) : ((~x7 | n4995) & (x3 | ~n664 | (~x6 ^ x7)));
  assign n4995 = (x0 | ~x4 | (x1 ? (~x3 | ~x6) : (x3 | x6))) & (~x0 | x1 | ~x3 | x4 | ~x6);
  assign z460 = ~n4999 | (~x1 & (x4 ? ~n4998 : ~n4997));
  assign n4997 = ((x6 ^ x7) | ((~x0 | x2 | ~x3 | ~x5) & (x0 | ~x2 | x3 | x5))) & (~x5 | ~x6 | x7 | x0 | x2 | ~x3) & (x3 | x5 | ((x2 | ~x6 | x7) & (~x0 | ((~x6 | x7) & (~x2 | x6 | ~x7)))));
  assign n4998 = (x0 | x2 | x3 | x5 | x6 | x7) & (~x2 | ((~x5 | x6 | x7 | ~x0 | x3) & (x0 | ~x7 | (x3 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n4999 = ~n5000 & ~n5001 & n5002 & ~n5004 & (x1 | n5005);
  assign n5000 = ~x2 & (((x1 ^ x4) & (x0 ? (~x3 & ~x7) : (x3 ^ x7))) | (x0 & x4 & x7 & (x1 ^ x3)));
  assign n5001 = ~n1007 & ((~x0 & ~x1 & x2 & x4 & ~x7) | (x0 & x7 & (x1 ? (~x2 & ~x4) : (x2 & x4))));
  assign n5002 = ~n664 | (n5003 & (~n563 | ~n1163));
  assign n5003 = (x2 | x3 | ~x4 | x5 | ~x7) & (~x3 | (~x5 ^ ~x7) | (~x2 ^ x4));
  assign n5004 = x2 & ((x3 & ((~x4 & x7 & x0 & ~x1) | (~x0 & (x1 ? (x4 & x7) : (~x4 & ~x7))))) | (~x0 & x1 & ~x3 & (x4 ^ x7)));
  assign n5005 = ((x0 ^ ~x7) | ((~x2 | ~x4 | (x3 ^ x5)) & (x4 | x5 | x2 | ~x3))) & (x3 | x4 | ~x5 | ((x0 | ~x2 | ~x7) & (x7 | (~x0 & x2))));
  assign z461 = n5007 | n5011 | n5014 | (x5 ? ~n5015 : ~n5010);
  assign n5007 = x0 & ((n539 & ~n5009) | (~x1 & ~n5008));
  assign n5008 = x2 ? (~x3 | ((~x6 | x7 | ~x4 | x5) & (x4 | ~x5 | x6 | ~x7))) : (x3 | ((x6 | x7 | x4 | x5) & (~x5 | ((~x6 | ~x7) & (~x4 | x6 | x7)))));
  assign n5009 = (~x3 | x4 | x5 | ~x6 | x7) & (x3 | ((x6 | ~x7 | ~x4 | ~x5) & (x4 | (x5 ? (~x6 | x7) : (x6 | ~x7)))));
  assign n5010 = (x2 | ((~x0 | ((~x3 | x4 | x6) & (x1 | x3 | ~x4))) & (x1 | ~x3 | x4) & (~x1 | ((x3 | x4 | ~x6) & (x0 | ~x4 | (~x3 & ~x6)))))) & (~x4 | x6 | x1 | ~x2) & (x0 | ~x1 | x4 | (x3 ? ~x2 : ~x6));
  assign n5011 = ~x0 & ((x1 & ~n5012) | (n670 & ~n5013));
  assign n5012 = (x2 | x3 | ~x5 | ~x6 | x7) & (~x7 | ((~x2 | ~x3 | ~x4 | x5 | ~x6) & (x2 | x6 | (x3 ? (x4 | ~x5) : x5))));
  assign n5013 = (~x5 | x6 | x7 | ~x3 | x4) & (x3 | ((x4 | x5 | ~x6 | ~x7) & (~x4 | (x5 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n5014 = ~n783 & ((~x3 & ~x5 & ~x1 & x2) | (x5 & ((x2 & ~x3 & ~x0 & x1) | (x0 & ~x2 & (x1 ^ x3)))));
  assign n5015 = ((~x2 ^ x3) | ((x1 | ~x4 | x6) & (x4 | ~x6 | x0 | ~x1))) & (~x3 | x4 | ~x6 | x1 | ~x2) & (x0 | (x1 ? (x2 ? (~x3 | ~x4) : (x3 | x6)) : (x2 ? (~x3 | x4) : (~x3 ^ ~x4))));
  assign z462 = (x2 | n5019 | ~n5020 | ~n5022) & (~x2 | ~n5017 | ~n5023);
  assign n5017 = (~x3 | n5018) & (n850 | ((x0 | x3 | ~x7) & (x1 | ((x3 | ~x7) & (~x0 | ~x3 | x7)))));
  assign n5018 = (x5 | ~x6 | x7 | x0 | ~x1 | ~x4) & (x4 | ~x7 | ((x1 | x5 | x6) & (x0 | ((x5 | x6) & (x1 | ~x5 | ~x6)))));
  assign n5019 = ~n846 & (x0 ? ((~x3 & ~x4 & ~x7) | (~x1 & x3 & x4 & x7)) : (x4 & ((~x3 & ~x7) | (x1 & x3 & x7))));
  assign n5020 = (x7 | n5021) & (x1 | ~x7 | (~n4827 & (x0 | n759)));
  assign n5021 = x3 ? (x4 | ((x0 | ~x5 | x6) & (x5 | ~x6 | ~x0 | ~x1))) : ((x1 ^ ~x6) | (x0 ? (~x4 | ~x5) : (x4 | x5)));
  assign n5022 = (x6 | ((x4 | ((~x1 | x3 | ~x5) & (~x0 | (x1 ? (~x3 | x5) : ~x5)))) & (x3 | ~x4 | ~x5 | (x0 & x1)))) & (x0 | x3 | x4 | ~x5 | ~x6) & (x5 | ((~x4 | ~x6 | ~x0 | x3) & (~x3 | ((x1 | ~x4 | ~x6) & (x0 | (~x6 & (x1 | ~x4)))))));
  assign n5023 = (x3 & ((x5 & ~x6) | (~x4 & (x5 | ~x6)))) | (~x3 & ((~x5 & x6) | (x4 & (~x5 | x6)))) | (x0 & x1) | (~x4 & x5 & ~x6) | (x4 & ~x5 & x6);
  assign z463 = n5025 | ~n5030 | (~n857 & ~n5029) | (~n662 & ~n5028);
  assign n5025 = ~x1 & ((n1317 & ~n5027) | (~x3 & ~n5026));
  assign n5026 = (x0 | ~x2 | x4 | x5 | x6 | ~x7) & (x7 | (x0 ? (x6 | (x2 ? (x4 | x5) : (~x4 | ~x5))) : (~x6 | (x2 ? (~x4 ^ x5) : (~x4 ^ ~x5)))));
  assign n5027 = (~x2 | x4 | ~x5 | ~x6 | x7) & (x2 | ~x7 | (x4 ? (~x5 ^ x6) : (x5 | x6)));
  assign n5028 = (x0 & ((x1 & (x3 | (~x4 & x5))) | (~x3 & ((~x2 & ~x4 & x5) | (~x5 & (x2 | x4)))))) | (~x0 & ((~x1 & ~x5 & (x4 ? x3 : ~x2)) | (x5 & ((~x3 & x4) | (x2 & x3 & ~x4))))) | (x4 & ((x2 & (~x3 | ~x5)) | (x5 & (x3 ? ~x2 : ~x1)))) | (~x2 & ~x4 & ((x3 & ~x5) | (x1 & ~x3 & x5)));
  assign n5029 = x2 ? (x5 | ((~x4 | ~x6 | x7) & (x3 | x4 | x6 | ~x7))) : (~x5 | ((x6 | ~x7 | ~x3 | ~x4) & (x3 | (x4 ? (~x6 | x7) : (x6 | ~x7)))));
  assign n5030 = ~n5032 & (~n1769 | ~n2010) & (x3 ? n5034 : n5031);
  assign n5031 = (x0 | x1 | x6 | ~x7 | (~x2 ^ ~x4)) & (x2 | x4 | ~x6 | x7 | (~x0 & ~x1));
  assign n5032 = ~n5033 & ((n923 & n543) | (n650 & n544));
  assign n5033 = (x0 | ~x1 | ~x2 | ~x5) & (~x0 | ((x2 | x5) & (x1 | ~x2 | ~x5)));
  assign n5034 = (~x0 | x1 | x2 | x4 | x6 | ~x7) & (~x4 | (x0 & x1) | (x2 ? (x6 | ~x7) : (~x6 | x7)));
  assign z464 = n5036 | ~n5041 | (~n620 & ~n5040) | (~n662 & ~n5039);
  assign n5036 = ~x2 & (x3 ? ~n5038 : (n738 & n5037));
  assign n5037 = x5 & (x4 ? ~x6 : (x6 & ~x7));
  assign n5038 = x0 ? ((~x1 | x4 | x5 | x6 | ~x7) & (x1 | ~x4 | ~x5 | ~x6 | x7)) : ((x1 | ~x4 | x5 | ~x6 | ~x7) & (~x1 | ~x5 | x7 | (~x4 ^ x6)));
  assign n5039 = (x1 | ((~x0 | (x2 ? (x4 | ~x5) : x5)) & (~x5 | ((~x2 | x3) & (x0 | x2 | ~x3 | ~x4))))) & (x3 | ~x5 | x0 | ~x2) & (x5 | ((~x1 | ((x0 | ~x3 | ~x4) & (x2 | x3))) & (x2 | x3 | ~x4) & (x0 | ~x3 | (x2 ^ x4))));
  assign n5040 = (x0 | ~x2 | x3 | x5 | (x1 ^ x4)) & (~x5 | ((~x3 | ~x4 | x0 | ~x2) & (x2 | ((x3 | ~x4 | x0 | x1) & (~x0 | x4 | (~x1 ^ x3))))));
  assign n5041 = ~n5046 & ~n5045 & ~n5044 & ~n5043 & ~n3809 & ~n5042;
  assign n5042 = ~n1226 & ((~x3 & (x0 ? (x1 ? (~x2 & x4) : (x2 & ~x4)) : (x1 & ~x4))) | (~x0 & ~x2 & x3 & (~x1 | x4)));
  assign n5043 = ~n630 & ((x2 & x3 & x4 & x0 & ~x1) | (~x0 & ~x4 & ((x2 & x3) | (~x1 & ~x2 & ~x3))));
  assign n5044 = ~n806 & ((~x2 & ~x3 & x6 & n664) | (x2 & x3 & (x6 ? n664 : n738)));
  assign n5045 = n709 & ((~x0 & ~x3 & x4 & n544) | (x0 & (x3 ? (~x4 & n544) : (x4 & n543))));
  assign n5046 = n538 & (x0 ? (n690 & n2503) : (~x6 & ~n2744));
  assign z465 = (~x2 & ~n5052) | (x2 & ~n5048) | (x3 & ~n5056) | (~x3 & ~n5055);
  assign n5048 = (n662 | n5051) & (x0 | n5049) & (n620 | n5050);
  assign n5049 = (~x5 | ~x6 | ~x7 | x1 | ~x3 | ~x4) & (x6 | ((~x3 | ((~x1 | (x4 ? (~x5 | ~x7) : (x5 | x7))) & (x5 | ~x7 | x1 | ~x4))) & (x1 | x3 | (x4 ? (~x5 | x7) : (x5 | ~x7)))));
  assign n5050 = x0 ? (x1 | (x3 ? (~x4 | ~x5) : (~x4 ^ x5))) : ((x4 | ~x5 | x1 | ~x3) & (~x1 | (x3 ? (~x4 | x5) : x4)));
  assign n5051 = (~x3 | x4 | ~x0 | x1) & (x0 | x3 | ~x4 | (x1 ^ x5));
  assign n5052 = x5 ? n5054 : n5053;
  assign n5053 = ((x1 ^ ~x3) | ((x6 | x7 | x0 | x4) & (~x7 | (x0 ? (~x4 ^ ~x6) : (x4 | ~x6))))) & (x7 | (x0 ? (x3 ? (x4 | ~x6) : (~x4 | x6)) : (~x4 | ((x3 | ~x6) & (~x1 | ~x3 | x6))))) & (x0 | ~x4 | ~x7 | (x1 ? (~x3 | ~x6) : (x3 | x6)));
  assign n5054 = x4 ? ((~x0 | x1 | ~x6 | (~x3 ^ ~x7)) & ((x1 ^ ~x3) | (x0 ? (x6 | x7) : (~x6 ^ x7)))) : (((x6 ^ x7) | (x0 ? (x1 | x3) : ~x3)) & (x0 | x7 | (x1 ? x6 : (x3 | ~x6))));
  assign n5055 = ((x4 ^ x6) | ((~x0 | x2 | (x1 ^ x5)) & (x0 | x1 | ~x2 | ~x5))) & (x0 | ~x1 | ((~x5 | ~x6 | x2 | x4) & (x5 | x6 | ~x2 | ~x4))) & (x1 | (x4 ? (~x5 | x6) : (x5 | ~x6)) | (x0 ^ x2));
  assign n5056 = (x1 | ((x4 | ~x5 | x6 | ~x0 | x2) & (~x4 | ((~x5 | x6 | x0 | ~x2) & (x5 | (x0 ? (~x2 ^ ~x6) : (x2 | ~x6))))))) & (x0 | ((~x1 | x2 | ~x4 | ~x5 | ~x6) & (x4 | ((~x2 | x5 | ~x6) & (~x1 | (x2 ? ~x6 : (x5 | x6)))))));
  assign z466 = n5058 | ~n5062 | ~n5066 | (~n662 & ~n5061);
  assign n5058 = ~x2 & ((n1421 & ~n5060) | (~x5 & ~n5059));
  assign n5059 = (~x1 | ((x0 | x3 | ~x4 | ~x6 | x7) & (~x0 | ~x3 | x4 | x6 | ~x7))) & (~x0 | x1 | ~x3 | ~x4 | (~x6 ^ x7));
  assign n5060 = (~x0 | x3 | ~x4 | ~x6 | x7) & (x0 | ((x3 | x4 | x6 | ~x7) & (~x6 | x7 | ~x3 | ~x4)));
  assign n5061 = ((x4 ^ x5) | ((~x0 | ~x1 | x2 | x3) & (x0 | ~x2 | (x1 ^ x3)))) & (x1 | ((~x0 | ((x3 | ~x4 | x5) & (x4 | ~x5 | ~x2 | ~x3))) & (~x4 | x5 | x2 | x3) & (x0 | ~x3 | (x2 ? (~x4 | x5) : (x4 | ~x5))))) & (x0 | ~x1 | ((x2 | ~x3 | ~x4 | x5) & (x3 | x4 | ~x5)));
  assign n5062 = ~n5063 & n5065 & (n806 | n2653) & (x1 | n5064);
  assign n5063 = ~n868 & ((~x0 & x1 & ~x2 & (x3 ^ ~x7)) | (~x1 & ((~x3 & x7 & ~x0 & ~x2) | (x0 & (x2 ? (~x3 & x7) : (x3 & ~x7))))));
  assign n5064 = x0 ? ((x2 | x3 | ~x4 | x6 | ~x7) & (~x2 | ~x3 | x4 | ~x6 | x7)) : (~x3 | ((x6 | ~x7 | ~x2 | ~x4) & (~x6 | x7 | x2 | x4)));
  assign n5065 = (~n943 | ~n2477) & (~n750 | (~n1308 & ~n1979));
  assign n5066 = (x1 | n5067) & (n627 | n5068);
  assign n5067 = ((~x5 ^ x7) | ((~x3 | x4 | x0 | ~x2) & (~x0 | (x2 ? (~x3 | ~x4) : (x3 | x4))))) & (x2 | ~x3 | ~x7 | (x0 ? (x4 | ~x5) : (~x4 | x5)));
  assign n5068 = (x3 | ~x6 | x7 | ~x0 | x1 | ~x2) & (x0 | x2 | ((~x6 | x7 | x1 | x3) & (~x1 | (x3 ? (~x6 | x7) : (x6 | ~x7)))));
  assign z467 = n5070 | ~n5073 | (n738 & ~n5078) | (x3 & ~n5077);
  assign n5070 = ~x0 & ((n537 & ~n5072) | (~x6 & ~n5071));
  assign n5071 = (x3 | ((x1 | x2 | x4 | ~x5 | ~x7) & (~x1 | ((x5 | ~x7 | x2 | ~x4) & (~x2 | x7 | (x4 & ~x5)))))) & (x1 | ~x3 | x7 | (x4 ? (~x2 & ~x5) : x2));
  assign n5072 = (~x5 | ((x1 | x2 | ~x3 | ~x4) & (~x1 | x3 | (x2 & ~x4)))) & (x4 | ((~x1 | x2 | ~x3 | x5) & (x1 | (x2 ? ~x3 : (x3 | x5)))));
  assign n5073 = (x3 | n5076) & (n620 | n5075) & (n627 | n5074);
  assign n5074 = (x3 | (x0 ? ((~x1 | x2 | ~x6 | ~x7) & (x6 | x7 | x1 | ~x2)) : ((x2 | x6 | x7) & (~x6 | ~x7 | x1 | ~x2)))) & (x0 | ~x1 | ((x2 | x6 | x7) & (~x6 | ~x7 | ~x2 | ~x3)));
  assign n5075 = x5 ? ((x1 | ~x3 | (x0 ? (~x2 ^ x4) : (x2 ^ x4))) & (x2 | x3 | x4 | ~x0 | ~x1) & (x0 | ((~x2 | x3 | x4) & (~x1 | (x2 ? x4 : (x3 | ~x4)))))) : ((x1 | (x0 ? (x2 ? (x3 | ~x4) : x4) : (x2 ? (~x3 | x4) : (x3 | ~x4)))) & (x2 | ~x3 | (x0 ? x4 : (~x1 | ~x4))));
  assign n5076 = x6 ? ((x0 | x1 | x2 | ~x4 | ~x5) & ((~x2 ^ ~x4) | (x0 ? (x1 | ~x5) : (~x1 | x5)))) : (x0 ? (x2 | ((~x4 | ~x5) & (~x1 | x4 | x5))) : (x1 | ~x2 | (~x4 ^ ~x5)));
  assign n5077 = (x0 | ~x1 | ~x2 | x4 | x5 | x6) & (~x4 | ((x1 | x5 | (x0 ? (~x2 ^ ~x6) : (x2 | ~x6))) & (x0 | ~x1 | ~x5 | (~x2 ^ x6))));
  assign n5078 = (x5 | ((x3 | x4 | ~x6 | ~x7) & (x2 | ((x4 | ~x6 | ~x7) & (x6 | x7 | x3 | ~x4))))) & (~x3 | ((x6 | x7 | ~x2 | x4) & (~x5 | ~x6 | ~x7 | (x2 & ~x4))));
  assign z468 = ~n5082 | ~n5084 | (x4 ? ~n5081 : (~x3 & ~n5080));
  assign n5080 = (~x2 | x5 | x7 | x0 | ~x1) & (x2 | ((x5 | x7 | ~x0 | x1) & (x0 | (x1 ? (~x5 ^ x7) : (~x5 | ~x7)))));
  assign n5081 = ((~x5 ^ x7) | ((x0 | ~x1 | x3) & (x1 | x2 | ~x3))) & (~x3 | ~x7 | ((~x0 | x1 | x5) & (x0 | ~x1 | ~x2 | ~x5)));
  assign n5082 = (~x0 | ~n539 | n2744) & (~n538 | (n2744 & (x7 | n5083)));
  assign n5083 = (x0 | x3 | ~x4 | ~x5 | x6) & (~x0 | ~x6 | (x3 ? (~x4 | ~x5) : (x4 | x5)));
  assign n5084 = ~n5085 & (n806 | n5088) & (n800 | n5089);
  assign n5085 = ~x2 & ((n738 & ~n5087) | (~x0 & ~n5086));
  assign n5086 = (((~x5 | ~x7 | x3 | ~x4) & (~x3 | x4 | x5 | x7)) | (x1 ^ x6)) & (x5 | ~x6 | x7 | x1 | x3) & (~x1 | ~x3 | ~x4 | ~x5 | x6 | ~x7);
  assign n5087 = x3 ? ((x5 | x6 | x7) & (~x4 | ~x5 | ~x6 | ~x7)) : (~x7 | ((x5 | ~x6) & (~x4 | ~x5 | x6)));
  assign n5088 = ((x1 ^ x6) | (x0 ? (x2 | x3) : ~x3)) & (~x2 | ((x3 | x6 | x0 | ~x1) & (x1 | (~x3 ^ x6))));
  assign n5089 = (x0 | (x1 ? ((~x3 | x4 | x6) & (~x2 | (x3 ? x6 : (x4 | ~x6)))) : ((~x2 | ~x3 | ~x6) & (x3 | x4 | x6)))) & (~x0 | ~x1 | x2 | x3 | x6) & (x1 | x4 | ((~x3 | ~x6) & (~x2 | x3 | x6)));
  assign z469 = n5091 | n5095 | n5099 | ~n5100 | (~x3 & ~n5098);
  assign n5091 = x4 & ((~x0 & ~n5092) | (~n620 & ~n5093) | (x0 & ~n5094));
  assign n5092 = x7 ? ((x6 | (x2 ^ x5) | (x1 ^ x3)) & (x2 | ~x5 | ~x6 | (~x1 & x3))) : ((~x1 | x2 | x3 | ~x5 | x6) & (x5 | ~x6 | ~x2 | ~x3));
  assign n5093 = x0 ? ((~x1 | x2 | x3 | ~x5) & (x1 | ~x2 | x5)) : ((~x2 | x3 | x5) & (x1 | ~x3 | (x2 ^ x5)));
  assign n5094 = (x5 | ~x6 | x7 | ~x1 | x2 | x3) & (x1 | ~x7 | ((~x5 | x6 | ~x2 | ~x3) & (x2 | ((~x3 | x5 | x6) & (~x5 | ~x6)))));
  assign n5095 = ~x4 & ((~n1215 & ~n1606) | (~x7 & ~n5097) | (x7 & ~n5096));
  assign n5096 = (~x0 | x1 | ~x3 | (x2 ? (x5 | ~x6) : (~x5 | x6))) & (x3 | ((x0 | ((~x2 | x5 | ~x6) & (x1 | x2 | ~x5 | x6))) & (~x0 | x1 | x2 | ~x5 | ~x6)));
  assign n5097 = (x1 | ((~x0 | ~x2 | ((x5 | x6) & (x3 | ~x5 | ~x6))) & (x2 | ~x5 | ~x6 | (x0 & ~x3)))) & (x0 | ((~x5 | ~x6 | x2 | ~x3) & (x6 | ((x5 | (~x2 ^ x3)) & (~x1 | ((~x3 | x5) & (x2 | x3 | ~x5)))))));
  assign n5098 = (~x0 | x1 | x5 | ~x6 | (~x2 ^ x4)) & (~x1 | ((x4 | ~x5 | ~x6 | ~x0 | x2) & (x0 | ((x2 | ~x4 | x5 | x6) & (~x5 | ~x6 | ~x2 | x4)))));
  assign n5099 = ~n857 & ((x5 & ~n4970) | (~x2 & ~x4 & ~x5 & ~n1185));
  assign n5100 = ~n5101 & (~n965 | ~n694) & (~n1546 | ~n1112);
  assign n5101 = ~x0 & ~x1 & ((x5 & x6 & x2 & ~x4) | (~x2 & (x4 ? (x5 & ~x6) : (~x5 & x6))));
  assign z470 = ~n5105 | ~n5110 | (~n846 & ~n5103) | (n664 & ~n5104);
  assign n5103 = x2 ? ((x1 | ((~x0 | (x3 ? (~x4 | x7) : (x4 | ~x7))) & (~x4 | x7 | x0 | x3))) & (x0 | ~x3 | x7 | (~x1 & x4))) : ((~x0 | ~x1 | x3 | x4 | x7) & (x0 | ~x3 | ~x7 | (x1 ^ x4)));
  assign n5104 = (~x2 | x3 | x4 | x5 | x6 | ~x7) & (x2 | ((~x3 | ~x6 | (x4 ? (x5 | x7) : (~x5 | ~x7))) & (x3 | ~x4 | ~x5 | x6 | x7)));
  assign n5105 = ~n5107 & ~n5108 & n5109 & (n912 | n5106);
  assign n5106 = (x2 | ((x7 | ((~x3 | ~x4 | ~x0 | x1) & (x0 | (x1 ? (~x3 | x4) : x3)))) & (~x0 | x3 | ~x7 | (~x1 & x4)))) & (x0 | ~x2 | ~x3 | ~x7 | (x1 & ~x4));
  assign n5107 = ~x1 & ((x0 & x2 & x3 & ~x5 & x7) | (~x0 & ((~x2 & x3 & x5 & ~x7) | (~x5 & x7 & x2 & ~x3))));
  assign n5108 = ~n1099 & ((~x0 & x1 & x2 & ~x5 & x7) | (x0 & ((~x2 & ~x5 & ~x7) | (~x1 & x5 & (x2 ^ x7)))));
  assign n5109 = (x2 | n824 | ~n2328) & (~n2205 | ((~n814 | ~n924) & (~x2 | ~n2328)));
  assign n5110 = x1 | (n5111 & ~n5112 & (x5 | n3446 | n1311));
  assign n5111 = (x0 | ((x2 | x3 | x4 | ~x5 | ~x7) & (~x2 | ~x3 | ~x4 | x5 | x7))) & (x3 | x4 | x7 | ((~x2 | ~x5) & (~x0 | x2 | x5)));
  assign n5112 = n2573 & (x0 ? (x3 & ~n1307) : (~x3 & n1844));
  assign z471 = ~n5116 | (~x0 & (x6 ? ~n5114 : ~n5115));
  assign n5114 = (x2 | ((x5 | ~x7 | x1 | ~x4) & (~x1 | ~x3 | (x4 ? (x5 | x7) : ~x5)))) & (x1 | ((x3 | ~x4 | x5 | x7) & (~x2 | x4 | ~x5 | (~x3 & x7))));
  assign n5115 = (~x1 | ((x2 | x3 | ~x4 | x5) & (~x2 | ~x3 | x4 | ~x5 | ~x7))) & (x2 | ((x3 | ~x4 | x5 | ~x7) & (x4 | ~x5 | x7 | x1 | ~x3)));
  assign n5116 = n5118 & (x1 ? n5123 : (n5122 & (~x0 | n5117)));
  assign n5117 = x2 ? ((x3 | ~x4 | x5 | ~x6 | ~x7) & (~x3 | x4 | ~x5 | x6 | x7)) : ((~x3 | ~x5 | ~x6 | (~x4 ^ ~x7)) & (x6 | (x3 ^ x7) | (~x4 ^ x5)));
  assign n5118 = n5121 & (n2500 | n5119) & (n1041 | n5120);
  assign n5119 = x0 ? (x6 | ((x2 | x7) & (x1 | (x2 & x7)))) : ((~x1 | x6 | ~x7) & (~x6 | (x1 & (x2 | x7))));
  assign n5120 = (~x0 | x1 | ~x2 | x3 | x5 | x7) & (x0 | ~x7 | ((x1 | x2 | ~x3 | ~x5) & (x3 | x5 | ~x1 | ~x2)));
  assign n5121 = (x0 | ~x1 | ~x2 | x7 | (~x3 ^ ~x6)) & (~x7 | ((~x2 | x3 | x6 | x0 | x1) & (~x0 | ((~x3 | x6 | x1 | ~x2) & (~x1 | x2 | x3 | ~x6)))));
  assign n5122 = (~x6 | (x0 ? (x3 ? (~x4 | x7) : (x4 | ~x7)) : ((~x4 | ~x7 | ~x2 | ~x3) & (x2 | x3 | x4 | x7)))) & (x0 | x6 | (x3 ? (~x4 | x7) : (x4 | (x2 ^ ~x7))));
  assign n5123 = (x4 | ~x6 | x7 | ~x0 | x2 | x3) & (x0 | ((x2 | x3 | x4 | x6) & (~x6 | ~x7 | ~x3 | ~x4)));
  assign z472 = n5128 | ~n5129 | n5132 | (~x2 & (~n5125 | ~n5131));
  assign n5125 = x4 ? n5126 : (x5 | n5127);
  assign n5126 = x3 ? (~x5 | x7 | ((x1 | ~x6) & (x0 | ~x1 | x6))) : (x5 | ((~x0 | x7 | (~x1 ^ x6)) & (~x7 | (x1 ^ x6))));
  assign n5127 = (~x0 | x6 | (x1 ? (~x3 | ~x7) : (x3 | x7))) & (x3 | ~x6 | ((~x1 | x7) & (x0 | x1 | ~x7)));
  assign n5128 = ~n927 & (x1 ? (~x2 & x5 & (~x0 | ~x3)) : ((x3 & ~x5) | (x2 & (x3 | ~x5))));
  assign n5129 = ~n5130 & (~n750 | ~n1144) & (~n534 | ~n2542);
  assign n5130 = ~x0 & x1 & x2 & ((x4 & ~x7) | (x3 & ~x4 & x7));
  assign n5131 = (x0 | ((~x5 | ~x7 | x1 | x4) & (~x1 | x5 | ((~x4 | x7) & (~x3 | x4 | ~x7))))) & (x1 | ~x5 | (x3 ? (x4 | ~x7) : (~x4 | x7)));
  assign n5132 = n601 & (((~x4 ^ x7) & (x6 ? n664 : ~x1)) | (~x4 & x7 & (x6 ? ~x1 : n664)));
  assign z473 = (x5 & ~n5134) | (~x5 & ~n5136) | (~x2 & ~n5139) | (x2 & ~n5140);
  assign n5134 = (~x4 | n5135) & (x3 | x4 | ~n543 | ~n924);
  assign n5135 = x7 ? (x0 ? ((~x3 | x6 | x1 | ~x2) & (~x1 | x2 | x3 | ~x6)) : ((x1 | x2 | x3 | ~x6) & (~x3 | x6 | ~x1 | ~x2))) : ((x0 & x1) | (x2 ? (x3 | ~x6) : (~x3 | x6)));
  assign n5136 = (x4 | n5138) & (n857 | n5137) & (~x4 | ~n544 | ~n947);
  assign n5137 = (~x4 | ~x6 | ~x7 | ~x2 | x3) & (x2 | x6 | (x3 ? (~x4 | ~x7) : (x4 | x7)));
  assign n5138 = x0 ? (~x1 | x2 | x7 | (~x3 ^ ~x6)) : (x1 | ~x7 | ((x3 | x6) & (~x2 | ~x3 | ~x6)));
  assign n5139 = (~x5 | ~x6 | x3 | x4) & (x5 | ((x0 | ((~x3 | ~x6) & (x1 | ~x4 | x6))) & (x3 | ~x4 | x6) & (~x3 | (x6 ? x1 : x4))));
  assign n5140 = (x4 & (x0 | x1) & (~x5 | (x3 & ~x6))) | (~x5 & (x3 | ~x6)) | (x0 & x1) | (~x3 & x5 & x6);
  assign z474 = (~x0 & (~n5143 | (~x4 & ~n5142))) | ~n5145;
  assign n5142 = (~x1 | ~x2 | ~x3 | x5 | ~x6 | ~x7) & (x2 | ((x5 | ~x6 | ~x7 | x1 | ~x3) & (x3 | ((x6 | ~x7 | x1 | x5) & (~x1 | (x5 ? (x6 | x7) : (~x6 | ~x7)))))));
  assign n5143 = (~n1902 | n910 | x3 | x4) & (~x4 | (n5144 & (~x3 | ~n1901 | n910)));
  assign n5144 = ((~x1 ^ ~x2) | ((x6 | x7 | x3 | x5) & (~x6 | ~x7 | ~x3 | ~x5))) & (x2 | ~x3 | ~x5 | x6 | x7) & (~x1 | ((x2 | ~x3 | ((x6 | x7) & (x5 | ~x6 | ~x7))) & (~x5 | ((~x3 | x6 | x7) & (x2 | x3 | ~x6 | ~x7)))));
  assign n5145 = ~n5146 & n5150 & (n620 | n5149) & (x1 | n5148);
  assign n5146 = x0 & ((~x1 & ~n5147) | (n1082 & n559));
  assign n5147 = (x2 | ((~x3 | ((~x6 | ~x7 | x4 | ~x5) & (~x4 | x6 | x7))) & (x6 | x7 | ~x4 | ~x5) & (x3 | x4 | x5 | (x6 ^ x7)))) & (~x3 | ~x4 | ((~x5 | x6 | x7) & (~x6 | ~x7 | (~x2 & x5))));
  assign n5148 = (x4 | ~x5 | x6 | x0 | x2 | x3) & (~x0 | ((x2 | x3 | ~x4 | ~x5 | ~x6) & (~x2 | x4 | (x3 ? ~x6 : (~x5 | x6)))));
  assign n5149 = (~x0 | ((x3 | ~x4 | x1 | ~x2) & (~x1 | x2 | ~x3 | x4 | x5))) & (x3 | ~x4 | ((~x5 | (x1 ^ ~x2)) & (x0 | (~x1 & x2)))) & (x0 | ~x3 | x4 | x5 | (x1 & ~x2));
  assign n5150 = (n5151 | (~x4 ^ x5)) & (n2322 | ((x0 | x4 | (~x1 & ~x5)) & (x1 | x5 | (~x0 ^ x4))));
  assign n5151 = (~x0 | x2 | x3 | x6) & (x0 | ~x2 | ~x3 | ~x6);
  assign z475 = ~n5157 | (x1 ? ~n5155 : (x0 ? ~n5154 : ~n5153));
  assign n5153 = (x5 | ((~x6 | ((x2 | (x3 ? (x4 | ~x7) : (~x4 | x7))) & (x4 | ~x7 | ~x2 | x3))) & (x2 | ~x3 | x6 | (~x4 ^ ~x7)))) & (~x2 | ~x3 | ~x5 | (x4 ? (~x6 ^ x7) : (x6 | x7)));
  assign n5154 = x2 ? ((x3 | x4 | ~x5 | x6 | ~x7) & (~x3 | ~x4 | x5 | ~x6 | x7)) : (~x3 | ~x5 | (x4 ? (x6 ^ x7) : (~x6 ^ x7)));
  assign n5155 = (~n2317 | ~n587) & (x5 | n5156);
  assign n5156 = (x3 | ((x7 | ((x4 | x6 | ~x0 | x2) & (x0 | ~x2 | (~x4 ^ ~x6)))) & (~x0 | x2 | ~x7 | (~x4 ^ x6)))) & (x0 | ~x2 | ~x7 | ((~x4 | x6) & (~x3 | x4 | ~x6)));
  assign n5157 = (x5 | n5160) & (n592 | n5159) & (~x5 | n5158);
  assign n5158 = (x0 | ~x1 | x2 | x3 | x7) & (x1 | ((~x3 | x4 | ~x7 | x0 | ~x2) & (~x0 | x3 | (x2 ? (~x4 | x7) : ~x7))));
  assign n5159 = ((~x2 ^ x3) | (x0 ? (x1 | x5) : ~x5)) & (x2 | ~x3 | x0 | ~x1) & (~x5 | (x0 ? (x1 ? (x2 | x3) : (~x2 | ~x3)) : (x1 ^ x3)));
  assign n5160 = (x1 | (((x4 ^ x7) | (x0 ? (x2 | x3) : ~x2)) & (x4 | ~x7 | (x0 ? (~x2 | ~x3) : (x2 | x3))))) & (~x3 | x4 | x7 | ~x0 | ~x1 | x2) & (x0 | ((x4 | x7 | ~x2 | ~x3) & (~x1 | x3 | (x2 ? (x4 | ~x7) : x7))));
  assign z476 = n5163 | ~n5165 | ~n5169 | (x0 & ~n5162);
  assign n5162 = (~x1 | x2 | x3 | ~x4 | ~x5 | x6) & (x1 | ((x2 | ~x5 | ~x6 | (~x3 & ~x4)) & (x5 | ((~x4 | x6 | x2 | ~x3) & (~x2 | (x3 ? (~x4 | ~x6) : (x4 | x6)))))));
  assign n5163 = x3 & ((n750 & n678) | (~x6 & n2512 & ~n5164));
  assign n5164 = (x0 | ~x2 | ~x5 | ~x7) & (x7 | (x0 ? (~x2 ^ ~x5) : (~x2 | x5)));
  assign n5165 = ~n5166 & ~n5168 & (n912 | n3377) & (x0 | n5167);
  assign n5166 = ~x1 & ((~x3 & x5 & ~x0 & x2) | (x0 & ((~x4 & x5 & ~x2 & ~x3) | (x2 & ~x5 & (x3 ^ x4)))));
  assign n5167 = x1 ? ((x2 | x3 | x5 | x6) & (~x2 | x4 | (x3 ? (~x5 | x6) : (x5 | ~x6)))) : ((x2 | x3 | x5 | ~x6) & (~x3 | ((x2 | ~x4 | ~x5 | x6) & (~x2 | ((~x5 | ~x6) & (~x4 | x5 | x6))))));
  assign n5168 = ~x0 & x1 & x3 & (x2 ? (x4 & x5) : ~x5);
  assign n5169 = (~x5 | ((x7 | n5170) & (x3 | ~x7 | n5171))) & (x5 | ~x7 | n5170) & (x3 | (~n5172 & (x5 | x7 | n5171)));
  assign n5170 = (x0 | ~x1 | ~x2 | x4 | (x3 ^ x6)) & (~x4 | (x0 ? ((x3 | ~x6 | ~x1 | x2) & (~x3 | x6 | x1 | ~x2)) : (x1 | x2 | (x3 ^ x6))));
  assign n5171 = (~x0 | x1 | (x2 ? (x4 | ~x6) : (~x4 | x6))) & (x0 | ~x1 | x2 | ~x4 | ~x6);
  assign n5172 = x7 & n1123 & ((x1 & ~x2 & x5 & x6) | (~x1 & ~x5 & (~x2 ^ x6)));
  assign z477 = n5174 | ~n5178 | (x2 & ~n5177);
  assign n5174 = ~x1 & (x0 ? ~n5176 : ~n5175);
  assign n5175 = x2 ? (~x7 | ((x4 | ~x5 | x6) & (x3 | x5 | (~x4 ^ x6)))) : ((x5 | ~x6 | x7 | x3 | ~x4) & (~x5 | (x3 ? (x4 ? (x6 | x7) : ~x6) : (x4 | x7))));
  assign n5176 = x2 ? (~x4 | ((x6 | x7 | x3 | x5) & (~x6 | ~x7 | ~x3 | ~x5))) : (x4 | ~x5 | ~x6 | (~x3 & x7));
  assign n5177 = (x1 | ((x7 | ((x0 | (x3 ? (x4 | ~x6) : x6)) & (x3 | x4 | x6) & (~x0 | ~x3 | ~x4 | ~x6))) & (~x0 | ~x7 | (x3 ? (~x4 | x6) : (x4 | ~x6))))) & (x0 | ~x1 | ((x6 | x7 | ~x3 | ~x4) & (x3 | ((~x6 | x7) & (x4 | x6 | ~x7)))));
  assign n5178 = ~n5180 & n5182 & (~n664 | n5179) & (~n549 | n5181);
  assign n5179 = (~x6 | (x2 ? (~x7 | (~x4 ^ x5)) : (x7 | (x3 ? (~x4 | ~x5) : (x4 | x5))))) & (~x5 | x6 | ((x2 | x4 | (~x3 & x7)) & (~x2 | ~x3 | ~x4 | ~x7)));
  assign n5180 = ~n2500 & (x1 ? ((~x2 & ~x6 & ~x7) | (x6 & x7 & ~x0 & x2)) : ((~x6 & ((x2 & x7) | (x0 & (x2 | x7)))) | (~x2 & x6 & (~x0 | ~x7))));
  assign n5181 = (x0 | x1 | ~x3 | ~x4 | ~x6) & (x3 | ((~x1 | ~x4 | ~x6) & (x0 | (x1 ^ x6))));
  assign n5182 = n5184 & (n5183 | ((~x4 | x5 | x2 | x3) & (x4 | ~x5 | ~x2 | ~x3)));
  assign n5183 = (x0 | ~x1 | x6 | x7) & (~x0 | x1 | (~x6 ^ x7));
  assign n5184 = (~x3 | ~x4 | ((x2 | ~x6 | ~x0 | x1) & (x0 | (x1 ? (x2 | x6) : (~x2 | ~x6))))) & (~x0 | x2 | x3 | x4 | (x1 ^ x6));
  assign z478 = ~n5190 | (x0 ? (n5189 | (~x2 & ~n5188)) : ~n5186);
  assign n5186 = (x2 | n5187) & (n918 | ((~x1 | ~x2 | x4 | x6) & (x1 | ~x4 | (x2 ^ x6))));
  assign n5187 = x3 ? ((~x4 | ((~x6 | ~x7 | x1 | x5) & (x6 | x7 | ~x1 | ~x5))) & (~x1 | x4 | x5 | (~x6 ^ x7))) : (x4 | (~x5 ^ x6) | (x1 ^ x7));
  assign n5188 = (x6 | ((x1 | x3 | x4 | ~x5 | x7) & (~x1 | x5 | (x3 ? (x4 | ~x7) : (~x4 | x7))))) & (x1 | ~x5 | ~x6 | (x3 ? (~x4 ^ ~x7) : (x4 | ~x7)));
  assign n5189 = x4 & n538 & (x3 ? (x5 & n543) : (~x5 & ~n620));
  assign n5190 = ~n5192 & n5194 & (x1 ? (x0 | n5193) : n5191);
  assign n5191 = x4 ? ((~x2 | ((~x5 | x7 | x0 | ~x3) & (~x0 | (x3 ? (x5 | ~x7) : (~x5 | x7))))) & (x0 | x2 | ~x7 | (x3 ^ x5))) : (x2 ? (x0 ? (~x3 | (x5 ^ x7)) : (x3 | (~x5 ^ x7))) : ((~x5 | ~x7 | x0 | x3) & (~x0 | x5 | (~x3 ^ ~x7))));
  assign n5192 = ~x2 & ((~x0 & x1 & ~x3 & x4 & x7) | (~x7 & ((x0 & (x1 ? (~x3 & ~x4) : (x3 & x4))) | (x3 & ~x4 & ~x0 & ~x1))));
  assign n5193 = (x5 | (~x3 ^ ~x4) | (x2 ^ x7)) & (~x3 | ~x5 | (x2 ? (~x4 | x7) : (x4 ^ x7)));
  assign n5194 = (~x3 | x4 | ~x7 | x0 | ~x2) & (x3 | ((~x4 | x7 | x0 | ~x2) & (~x0 | ~x7 | ((x2 | ~x4) & (x1 | ~x2 | x4)))));
  assign z479 = n5196 | n5200 | ~n5203 | (x1 ? ~n5202 : ~n5199);
  assign n5196 = ~x2 & (x5 ? ~n5197 : ~n5198);
  assign n5197 = (x1 | ((~x4 | ~x6 | ~x7 | x0 | ~x3) & (x7 | ((~x4 | x6 | ~x0 | x3) & ((~x4 ^ ~x6) | (x0 ^ x3)))))) & (x0 | ~x1 | (x4 ? (x6 | (~x3 ^ x7)) : (~x6 | ~x7)));
  assign n5198 = (~x0 | ~x1 | ~x3 | x4 | ~x6 | x7) & (x3 | ((~x0 | ~x4 | (x1 ? (x6 | x7) : (~x6 | ~x7))) & (x4 | ((x1 | x6 | ~x7) & (~x6 | x7 | x0 | ~x1)))));
  assign n5199 = x4 ? (x6 | (x0 ? ((~x3 | ~x5) & (~x2 | x3 | x5)) : ((x3 | ~x5) & (x2 | ~x3 | x5)))) : (x3 ? (x0 ? (x5 | x6) : (~x5 | (x2 & x6))) : ((~x0 | x2 | (~x5 ^ x6)) & (~x2 | (x0 ? (~x5 | ~x6) : (x5 | x6)))));
  assign n5200 = x2 & ((n738 & ~n4319) | (~x0 & ~n5201));
  assign n5201 = x7 ? ((~x4 | x5 | x6 | x1 | x3) & (~x1 | ~x3 | x4 | ~x5 | ~x6)) : ((x3 ? (x5 | x6) : (~x5 | ~x6)) | (~x1 ^ x4));
  assign n5202 = ((~x3 ^ x5) | ((~x0 | x2 | x4 | x6) & (x0 | ~x4 | ~x6))) & (x0 | x5 | ((x2 | x3 | x4 | x6) & (~x2 | (x3 ? ~x4 : (x4 | ~x6)))));
  assign n5203 = (x0 | ~x1 | x6 | (x2 ? (x3 | ~x5) : (~x3 | x5))) & (~x6 | (x0 ? ((~x1 | x2 | x3 | ~x5) & (x1 | ~x3 | x5)) : (x1 | ((x3 | x5) & (~x2 | ~x3 | ~x5)))));
  assign z480 = ~n5210 | (x7 ? ~n5207 : (n5206 | (~x4 & ~n5205)));
  assign n5205 = (~x2 | ((x0 | ~x1 | x6) & (~x3 | x5 | ~x6 | ~x0 | x1))) & (x0 | ~x1 | ((~x3 | x5 | x6) & (~x5 | ~x6 | x2 | x3))) & (x1 | x6 | ((x2 | x3 | ~x5) & (~x0 | ((x3 | ~x5) & (x2 | (x3 & ~x5))))));
  assign n5206 = x4 & n664 & ((~x2 & ((~x5 & x6) | (x3 & x5 & ~x6))) | (x6 & ((x2 & x3 & x5) | (~x3 & ~x5))));
  assign n5207 = (~n1205 | n5209) & (n783 | n5208);
  assign n5208 = (~x0 | x1 | x2 | x3 | ~x5) & (x0 | ~x1 | x5 | (~x2 ^ x3));
  assign n5209 = (x1 | x2 | x3 | x4 | ~x5) & (~x1 | ~x4 | ((~x3 | ~x5) & (x2 | x3 | x5) & (~x2 | (~x3 & ~x5))));
  assign n5210 = x6 ? ((x7 | n5212) & (x4 | (x7 ? n5213 : n5211))) : ((~x7 | n5212) & (~x4 | (x7 ? n5211 : n5213)));
  assign n5211 = (~x0 | x3 | (x1 ? (x2 | ~x5) : (~x2 | x5))) & (x1 | ((x2 | ~x3 | x5) & (x0 | (x2 ? (~x3 | ~x5) : x5))));
  assign n5212 = x1 ? ((x0 | ((~x3 | x4 | ~x5) & (~x2 | ((x4 | ~x5) & (~x3 | ~x4 | x5))))) & (x2 | x4 | x5 | (~x0 & x3))) : ((x4 | x5 | x0 | ~x2) & (~x4 | ((~x5 | (x2 & x3)) & (~x0 | (~x5 & (x2 | x3))))));
  assign n5213 = (~x2 & ((~x1 & ~x3 & x5) | (x0 & (x3 ? x5 : ~x1)))) | (x1 & (x2 | x3 | (~x0 & ~x5)));
  assign z481 = ~n5220 | (~n846 & ~n5218) | (~x1 & (~n5215 | ~n5219));
  assign n5215 = x3 ? n5217 : n5216;
  assign n5216 = (~x7 | ((x0 | x2 | x4 | x5 | x6) & ((~x5 ^ x6) | (x0 ? (x2 | x4) : ~x2)))) & (~x0 | ~x4 | ~x5 | ~x6 | (x2 & x7));
  assign n5217 = (x0 | x2 | x4 | ~x5 | ~x6 | x7) & (~x2 | ~x7 | ((x0 | ((x5 | ~x6) & (x4 | ~x5 | x6))) & (~x4 | ((x5 | ~x6) & (~x0 | ~x5 | x6)))));
  assign n5218 = (x1 | ~x3 | ((~x4 | x7 | x0 | x2) & (~x0 | (x2 ? x7 : (x4 | ~x7))))) & (x0 | ((~x2 | x3 | x7) & (~x1 | ((~x2 | x4 | x7) & (~x4 | ~x7 | x2 | x3)))));
  assign n5219 = (~x0 | ((x7 | ((~x2 | x3 | x4 | ~x5) & (x2 | (x3 ^ x5)))) & (~x2 | x5 | ~x7 | (x3 & x4)))) & (~x4 | x5 | ~x7 | x2 | ~x3) & (x0 | ((~x3 | (x2 ? ((~x4 | ~x5 | ~x7) & (x5 | x7)) : (x5 | ~x7))) & (x2 | ((~x4 | x5 | ~x7) & (x3 | ~x5 | x7)))));
  assign n5220 = ~x1 | ((~n559 | ~n1415) & n5221 & (~x7 | n5222));
  assign n5221 = (x2 | ((x7 | ((x5 | (x0 ? (~x3 ^ x4) : (x3 | x4))) & (x0 | ~x5 | (~x3 & ~x4)))) & (x0 | ~x7 | (x3 ? x5 : (x4 | ~x5))))) & (x0 | ~x2 | x5 | (x3 ? (~x4 | x7) : ~x7));
  assign n5222 = (x0 | ~x2 | ~x4 | ~x5 | x6) & ((x0 ? (x2 | x3) : (~x2 | ~x3)) | (~x5 ^ x6));
  assign z482 = ~n5226 | (~x2 & (x4 ? ~n5225 : ~n5224));
  assign n5224 = (x5 | ((x0 | x1 | x3 | ~x6 | ~x7) & (x7 | ((x0 | x1 | ~x3 | x6) & (~x1 | (x0 ? (~x3 ^ x6) : (x3 | x6))))))) & (x0 | x1 | ~x5 | (x3 ? (~x6 | x7) : x6));
  assign n5225 = (x0 | ~x1 | ~x3 | ~x5 | ~x6 | x7) & (~x0 | x1 | x6 | (x3 ? (~x5 | ~x7) : x5));
  assign n5226 = (n662 | n5230) & (x2 ? (n5228 & n5231) : n5227);
  assign n5227 = x0 ? ((~x1 | x3 | x4 | ~x6 | ~x7) & (x1 | ~x3 | ~x4 | x6 | x7)) : ((x1 | ~x3 | ~x4 | ~x6 | x7) & (x6 | ((~x1 | (~x3 & (x4 | ~x7))) & (~x3 | ~x7) & (x1 | x3 | ~x4))));
  assign n5228 = (x1 | n5229) & (~n2756 | (~n2467 & (x3 | n846)));
  assign n5229 = (x0 | ~x3 | ~x4 | ~x5 | x6) & (~x0 | ((x3 | ~x4 | x5 | x6 | x7) & (~x3 | x4 | ~x5 | ~x6 | ~x7)));
  assign n5230 = (x2 | ((~x0 | ((x3 | ~x4 | ~x5) & (x1 | x4))) & (~x1 | x3 | (~x4 & (x0 | ~x5))))) & (x0 | ~x2 | ~x3 | (x1 ^ (x4 & x5)));
  assign n5231 = (x0 | ((~x1 | x4 | (x3 ? ~x6 : (x6 | ~x7))) & (x3 | ~x6 | (x1 & x7)))) & (x1 | ((x3 | ~x4 | ~x6 | x7) & (~x0 | ((~x3 | ~x6 | (~x4 & x7)) & (x6 | ((x4 | ~x7) & (x3 | (x4 & ~x7))))))));
  assign z483 = ~n5239 | (x2 ? (~n5233 | ~n5238) : (~n5235 | ~n5237));
  assign n5233 = (x1 | n5234) & (~x3 | ~x4 | ~n2488 | x0 | ~x1);
  assign n5234 = x0 ? (x6 | ((~x5 | ~x7 | ~x3 | x4) & (x3 | ~x4 | x5 | x7))) : (~x6 | ((~x5 | x7 | ~x3 | ~x4) & (x3 | (x4 ? (~x5 | ~x7) : (x5 | x7)))));
  assign n5235 = ~n5236 & (n1107 | ((x4 | ~x6 | x0 | x1) & (~x0 | x6 | (x1 ^ ~x4))));
  assign n5236 = x5 & n664 & (n4635 | (x3 & x4 & ~n662));
  assign n5237 = ((x5 ^ x7) | ((~x3 | x4 | x0 | x1) & (~x0 | x3 | (~x1 ^ x4)))) & (~x0 | x1 | ~x3 | ~x4 | ~x5 | x7) & (x0 | x5 | ((x1 | x3 | x4 | ~x7) & (~x4 | x7 | ~x1 | ~x3)));
  assign n5238 = (x0 | ~x1 | ~x4 | (x3 ? (~x5 | ~x7) : (~x5 ^ x7))) & (x1 | ((~x0 | ~x3 | x4 | x5 | ~x7) & (x0 | ((~x5 | x7 | x3 | x4) & (x5 | ~x7 | ~x3 | ~x4)))));
  assign n5239 = x1 ? ((x2 | ((x3 | ~x4 | ~x7) & (x0 | x4 | x7))) & (x0 | x4 | ((~x3 | x7) & (~x2 | x3 | ~x7)))) : (x7 ? (x0 ? (x2 ? (x3 | ~x4) : x4) : (~x3 | (~x2 ^ x4))) : (x0 ? (~x2 | (~x3 ^ ~x4)) : (x3 | ~x4)));
  assign z484 = n5241 | ~n5242 | ~n5244 | (x1 ? ~n5249 : ~n5248);
  assign n5241 = x2 & ((~x1 & (x0 ? (~x4 & (x3 ^ x5)) : (x4 & ~x5))) | (~x0 & ((~x3 & x4 & ~x5) | (~x4 & x5 & x1 & x3))));
  assign n5242 = ~n5243 & (n2322 | ((~n738 | ~n2743) & (~n1123 | n3713)));
  assign n5243 = ~x2 & ((x0 & ~x4 & (x1 ? (~x3 & ~x5) : x5)) | (x4 & ((x1 & ~x3 & x5) | (~x0 & (x1 ? (x3 & ~x5) : x5)))));
  assign n5244 = x0 ? (x4 | n5247) : (~n5246 & (~x2 | n5245));
  assign n5245 = (x5 | ~x6 | ~x7 | ~x1 | ~x3 | x4) & (x1 | ~x4 | ~x5 | x7 | (~x3 ^ x6));
  assign n5246 = n563 & ((~x1 & ~x4 & ~x6 & ~n800) | (x1 & ~n1465));
  assign n5247 = (x1 | ~x2 | ~x3 | ~x5 | ~x6 | x7) & (x2 | ((x1 | x3 | x5 | x6 | ~x7) & (~x1 | x7 | (x3 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n5248 = x4 ? ((x0 | ~x2 | x3 | ~x5 | x6) & (~x3 | ((~x0 | (x2 ? (~x5 | ~x6) : (x5 | x6))) & (x5 | ~x6 | x0 | x2)))) : ((~x0 | ((x3 | x5 | ~x6) & (~x5 | x6 | ~x2 | ~x3))) & (x0 | ~x3 | (x2 ? (~x5 | ~x6) : (x5 | x6))) & (x2 | x3 | x5 | ~x6));
  assign n5249 = (~x0 | x2 | ~x3 | x4 | x5 | x6) & (x0 | (x2 ? ((~x5 | ~x6 | x3 | x4) & (x5 | x6 | ~x3 | ~x4)) : ((~x5 | x6 | ~x3 | ~x4) & (x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))))));
  assign z485 = n5251 | ~n5254 | n5260 | ~n5261 | (~x2 & ~n5259);
  assign n5251 = ~x4 & ((n738 & n1136 & ~n5253) | (x1 & ~n5252));
  assign n5252 = (x0 | x3 | x6 | ((x5 | ~x7) & (~x2 | ~x5 | x7))) & (x2 | ((~x5 | ~x6 | ~x7 | x0 | x3) & (~x0 | x7 | (x3 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n5253 = (~x5 | ~x7) & (x2 | x5 | x7);
  assign n5254 = ~n5256 & ~n5257 & ~n5258 & (n868 | n5255);
  assign n5255 = (x0 | ~x1 | x2 | x3 | ~x6) & (~x0 | x1 | (x2 ? (x3 | x6) : (~x3 | ~x6)));
  assign n5256 = ~x2 & (x0 ? (~x5 & (x1 ? (~x3 & x6) : (x3 & ~x6))) : (x3 & x5 & (~x1 ^ ~x6)));
  assign n5257 = (x3 ^ x6) & ((x0 & ~x1 & x2 & x5) | (~x0 & ~x5 & (x1 ^ ~x2)));
  assign n5258 = n2238 & n610 & (n644 | (~x1 & ~x7 & ~n785));
  assign n5259 = x0 ? (x4 | ((x1 | x3 | ~x5 | ~x6) & (x5 | x6 | ~x1 | ~x3))) : (~x4 | ((x1 | x3 | x5 | x6) & (~x1 | (x3 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n5260 = n616 & ((x4 & x5 & x6 & x1 & x3) | (~x1 & (x3 ? (x4 ? (~x5 & x6) : (x5 & ~x6)) : (x5 & (x4 ^ x6)))));
  assign n5261 = x2 ? (x7 ? n5262 : n5263) : (x7 ? n5263 : n5262);
  assign n5262 = (~x4 | x5 | ~x6 | ~x0 | x1 | ~x3) & (x0 | (x1 ? ((x3 | ~x4 | x5 | x6) & (~x5 | ~x6 | ~x3 | x4)) : (x4 | (x3 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n5263 = (x4 | ~x5 | ~x6 | ~x0 | x1 | ~x3) & (x0 | ((~x3 | ((x5 | ~x6 | ~x1 | x4) & (x1 | ~x4 | ~x5 | x6))) & (x1 | x3 | (x4 ? (~x5 | ~x6) : (x5 | x6)))));
  assign z486 = ~n5265 | (~x3 & ~n5271) | (~x0 & ~n5272);
  assign n5265 = ~n5266 & n5270 & (~x3 | n5269) & (n662 | n5268);
  assign n5266 = ~x2 & ((n837 & n958) | (x3 & ~n5267));
  assign n5267 = (~x0 | ((~x1 | x4 | x5 | ~x6 | x7) & (~x5 | x6 | ~x7 | x1 | ~x4))) & (x0 | ~x1 | ~x4 | x5 | x6 | ~x7);
  assign n5268 = (~x3 | ~x4 | ~x5 | x0 | x1) & (x3 | (x0 ? (x4 ? (x5 | (x1 ^ ~x2)) : ((x2 | ~x5) & (x1 | (x2 & ~x5)))) : (x4 | ((~x2 | x5) & (~x1 | (~x2 & x5))))));
  assign n5269 = (x1 | ((~x0 | ((~x5 | x6 | ~x2 | ~x4) & (x4 | x5 | ~x6))) & (x5 | x6 | x0 | ~x4))) & (x0 | ~x4 | x6 | (x5 ? ~x1 : ~x2));
  assign n5270 = (~n1812 | ~n598 | ~n1163) & (n627 | n620 | ~n1021);
  assign n5271 = x4 ? (~x6 | ((x0 | (~x1 & x5)) & (~x1 | x2 | ~x5) & (x1 | (x5 ? ~x0 : x2)))) : (x0 ? (x5 | x6 | (x1 ^ ~x2)) : (~x5 | ~x6 | (x1 & x2)));
  assign n5272 = (~x3 | x4 | x6 | ~x7) & (x7 | ((~x1 | ((~x3 | x4 | ~x6) & (x5 | x6 | x3 | ~x4))) & (~x3 | x4 | x5 | ~x6) & (x1 | x3 | ~x5 | (x4 ^ x6))));
  assign z487 = n5277 | n5278 | ~n5279 | ~n5282 | (~x7 & ~n5274);
  assign n5274 = (n1041 | n5276) & (~x0 | ~n538 | ~n1179) & (x0 | n5275);
  assign n5275 = (x5 | ((x3 | x4 | ~x6 | x1 | x2) & (~x1 | ((x2 | x3 | ~x4 | x6) & (x4 | ~x6 | ~x2 | ~x3))))) & (x1 | ~x5 | (x4 ? (~x6 | (x2 & x3)) : x6));
  assign n5276 = (~x0 | x1 | x2 | ~x3 | ~x5) & (x0 | ~x1 | x5 | (~x2 ^ x3));
  assign n5277 = ~n857 & ((x2 & x3 & ~x4 & x5 & ~x7) | (~x2 & ~x3 & (x4 ? (x5 & x7) : (~x5 & ~x7))));
  assign n5278 = ~n2465 & ((x4 & x5 & x7 & n664) | (~x4 & (x5 ? (~x7 & n664) : (x7 & n738))));
  assign n5279 = (x5 | (x7 ? (~n545 | n2113) : n5280)) & n5281 & (~x5 | ~x7 | n5280);
  assign n5280 = (~x0 | ~x1 | x2 | x3 | ~x4) & (x1 | (~x2 & ~x3) | (x0 ^ x4));
  assign n5281 = (~n1415 | ~n745) & (~n753 | ~n1546);
  assign n5282 = ~x7 | (n5283 & (x2 | n5284));
  assign n5283 = (~x3 | ~x4 | ~x5 | x0 | ~x1 | ~x2) & (x5 | ((x1 | x2 | x3 | ~x4) & (~x0 | x4 | (x1 ? (x2 | x3) : (~x2 | ~x3)))));
  assign n5284 = (~x0 | ~x1 | ~x3 | x4 | x5 | x6) & (x0 | x3 | (x1 ? (x4 ? (x5 | ~x6) : (~x5 | x6)) : (~x5 | (~x4 ^ x6))));
  assign z488 = n5287 | n5291 | ~n5292 | (~x6 & (~n5286 | ~n5290));
  assign n5286 = (x5 | ((~x0 | ((~x3 | x7 | x1 | ~x2) & (~x1 | x2 | x3))) & (x1 | x2 | ~x3 | ~x7) & (~x1 | x3 | ((x2 | ~x7) & (x0 | ~x2 | x7))))) & (x0 | ~x5 | (~x2 ^ x7) | (x1 ^ x3));
  assign n5287 = ~x2 & ((~n620 & ~n5288) | (~x4 & ~n5289));
  assign n5288 = (x0 | ~x1 | x3 | ~x4 | ~x5) & (~x0 | x4 | (x1 ? (~x3 | x5) : (x3 | ~x5)));
  assign n5289 = (~x0 | ((x1 | x3 | ~x5 | ~x6 | ~x7) & (~x1 | ~x3 | x5 | x6 | x7))) & (x0 | ~x1 | x3 | x5 | ~x6);
  assign n5290 = (x1 | (x2 ? (x5 | ~x7) : (~x5 | x7))) & (x0 | ~x1 | (x2 ? (~x5 | ~x7) : (x5 | x7)));
  assign n5291 = n2327 & n540 & ((~x3 & x5 & x0 & ~x1) | (~x0 & x3 & (x1 ^ x5)));
  assign n5292 = ~n5293 & (~n2825 | n5294);
  assign n5293 = x6 & ((~x1 & x2 & ~x5) | (~x0 & (x1 ? (x5 & (x2 | x7)) : ~x5)));
  assign n5294 = (~x0 | x5 | (x1 ^ ~x3)) & (x0 | ~x1 | ~x3 | ~x5 | x7);
  assign z489 = ~n5298 | (~x7 & (n5297 | (~x5 & ~n5296)));
  assign n5296 = (~x2 | x6 | ((x0 | ~x3 | (~x1 ^ x4)) & (x3 | ~x4 | ~x0 | x1))) & (~x0 | x2 | ~x6 | (x1 ? (~x3 | x4) : (x3 | ~x4)));
  assign n5297 = x5 & n605 & (x0 ? (x2 & n641) : (~x2 & n642));
  assign n5298 = ~n5300 & ~n5301 & ~n5302 & n5303 & (x7 | n5299);
  assign n5299 = (x1 | ((~x3 | ~x4 | ~x6 | x0 | ~x2) & (x4 | ((~x3 | x6 | x0 | ~x2) & (~x0 | x3 | (~x2 ^ x6)))))) & (x0 | x2 | x3 | ((~x4 | x6) & (~x1 | x4 | ~x6)));
  assign n5300 = ~x1 & ((x3 & ((x2 & x6 & x7) | (x0 & (x2 ? x6 : (~x6 & ~x7))))) | (~x2 & ~x3 & x7 & (~x0 ^ x6)));
  assign n5301 = n975 & ~n1041 & x7 & ~x3 & ~x5;
  assign n5302 = (x2 ^ x3) & ((~x1 & x6 & x7) | (~x0 & (~x6 ^ x7)));
  assign n5303 = ~x6 | ((~x7 | ~n923 | ~n924) & (~x1 | n1606));
  assign z490 = ~n5310 | ~n5308 | n5305 | n5307;
  assign n5305 = x4 & ((n1343 & n540 & n1546) | (~x3 & ~n5306));
  assign n5306 = (x0 | ~x1 | x2 | x5 | x6 | ~x7) & (~x6 | ((x0 | ~x1 | x2 | x5 | x7) & (~x0 | x1 | (x2 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n5307 = ~x1 & ((~x4 & ((x3 & ~x7 & ~x0 & x2) | (x0 & ~x3 & (x2 ^ x7)))) | (~x0 & x3 & x4 & (x2 ^ ~x7)));
  assign n5308 = (x2 | (x0 ? (x1 ? (x3 | ~x7) : (~x3 | x7)) : (x1 ? (~x3 | x7) : (x3 | ~x7)))) & n5309 & (~x2 | ((x0 | x3 | x7) & (~x3 | ~x7 | ~x0 | x1)));
  assign n5309 = (~x7 | ~n664 | n2286) & (x5 | ~n1035 | (~x2 ^ x7));
  assign n5310 = x5 ? n5311 : (~n650 | n5312);
  assign n5311 = (x3 | ~x4 | ~x7 | ~x0 | x1 | ~x2) & (x0 | ((x1 | x2 | ~x3 | x4 | x7) & (~x1 | ((~x4 | x7 | x2 | x3) & (x4 | ~x7 | ~x2 | ~x3)))));
  assign n5312 = (~x0 | ~x1 | x2 | x6 | ~x7) & (x0 | ((x1 | x2 | ~x6 | x7) & (~x1 | ~x2 | (~x6 ^ ~x7))));
  assign z491 = n5314 | (n538 & ~n5318) | (~x0 & ~n5316) | (x0 & ~n5317);
  assign n5314 = ~x2 & ((~x4 & ~n5315) | (n568 & n586));
  assign n5315 = (~x3 | ((x0 | x1 | x5 | x6 | x7) & (~x0 | ~x6 | (x1 ? (x5 | x7) : (~x5 | ~x7))))) & (x0 | x3 | ~x7 | (x1 ? (~x5 | ~x6) : (x5 | x6)));
  assign n5316 = (~x1 | ((~x2 | x3) & (~x4 | ~x5 | ~x6 | x2 | ~x3))) & (x3 | ((x1 | x2 | (~x5 & ~x6)) & (~x4 | x5 | x6) & (~x2 | (~x4 & (~x5 | ~x6))))) & (~x2 | ~x3 | x4 | (x1 & (x5 | x6)));
  assign n5317 = (x2 | ((~x1 | (x3 & (x4 | x5 | x6))) & (x1 | ~x3 | ~x4) & (x3 | (x4 ? x5 : (~x5 | ~x6))))) & (x1 | x3 | (x4 ? (x5 | x6) : ~x2));
  assign n5318 = (x0 | x3 | x4 | ~x5 | x6 | ~x7) & (~x4 | ((x0 | ~x3 | x5 | x6 | x7) & (~x0 | ~x6 | (x3 ? (~x5 | ~x7) : (x5 | x7)))));
  assign z492 = n5321 | ~n5323 | n5326 | ~n5327 | (n538 & ~n5320);
  assign n5320 = x3 ? ((x0 | ~x4 | x5 | x6 | x7) & (~x0 | ~x5 | (x4 ? (~x6 | x7) : (x6 | ~x7)))) : (x0 ? (x5 | (x4 ? (~x6 | x7) : (x6 | ~x7))) : (~x5 | (x4 ? (~x6 | ~x7) : (x6 | x7))));
  assign n5321 = ~x2 & (n5322 | (x3 & ~x5 & n598 & ~n1307));
  assign n5322 = ~n1243 & ((~x0 & ~x3 & ~x4 & x6 & x7) | (x0 & ((x3 & ~x4 & x6 & ~x7) | (~x6 & x7 & ~x3 & x4))));
  assign n5323 = ~n5324 & n5325 & (n1475 | n2136) & (~n750 | ~n1112);
  assign n5324 = ~x0 & ((x1 & x2 & x4 & x5) | (~x1 & (x2 ? (~x4 & ~x5) : (x4 & x5))));
  assign n5325 = ~x0 | x2 | ((x1 | x4 | x5) & (~x4 | ~x5 | ~x1 | x3));
  assign n5326 = n651 & ((~n2730 & ~n1243) | (n605 & n983));
  assign n5327 = ~n5328 & (n2354 | n5329);
  assign n5328 = ~x0 & (x1 ? ((x4 & ~x5 & x2 & ~x3) | (~x2 & x3 & ~x4 & x5)) : ((x4 & ~x5 & ~x2 & ~x3) | (~x4 & x5 & x2 & x3)));
  assign n5329 = (x0 | ~x1 | x2 | ~x4 | x6) & (~x0 | x1 | ~x2 | (~x4 ^ x6));
  assign z493 = ~n5334 | ~n5335 | (x4 & ~n5333) | (x1 & ~n5331);
  assign n5331 = (x5 | x7 | n571 | ~x0 | x2) & (x0 | (n5332 & (~x7 | n571 | ~x2 | ~x5)));
  assign n5332 = (x2 | ~x3 | ~x4 | x5 | x6 | ~x7) & (x3 | ~x6 | ((x5 | ~x7 | ~x2 | x4) & (x2 | ((~x5 | ~x7) & (x4 | x5 | x7)))));
  assign n5333 = x0 ? (x1 | ((~x5 | ~x6 | x2 | ~x3) & (~x2 | x6 | (~x3 ^ ~x5)))) : ((~x3 | ((x1 | x2 | x5 | x6) & (~x1 | (x2 ? (x5 | ~x6) : (~x5 | x6))))) & (x1 | x3 | ~x5 | (~x2 ^ x6)));
  assign n5334 = x1 ? ((x3 | ~x5 | ~x6 | ~x0 | x2) & (x0 | (x2 ? (x3 ? (x5 | x6) : (~x5 | ~x6)) : (x5 | (x3 ^ x6))))) : ((~x3 | ~x5 | ~x6 | x0 | ~x2) & ((~x0 ^ ~x3) | (x2 ? (x5 | ~x6) : (~x5 | x6))));
  assign n5335 = (x4 | n5336) & (x1 | (~n5337 & (x7 | n5338)));
  assign n5336 = (x6 | ((~x0 | ((~x3 | x5 | x1 | ~x2) & (x2 | x3 | ~x5))) & (x0 | x1 | ~x2 | (~x3 ^ ~x5)) & (~x1 | ((x2 | ~x3 | x5) & (x3 | ~x5 | x0 | ~x2))))) & (x1 | ~x6 | ((x2 | ((x3 | x5) & (x0 | ~x3 | ~x5))) & (~x0 | (x2 ? (x3 | ~x5) : x5))));
  assign n5337 = ~n783 & ((x0 & ~x2 & ~x3 & ~x5 & x7) | (~x7 & ((x3 & ~x5 & ~x0 & ~x2) | (x2 & (x0 ? (x3 ^ ~x5) : (~x3 & x5))))));
  assign n5338 = (x0 | ~x2 | ~x3 | ~x4 | x5 | x6) & (x2 | ~x5 | ((x4 | ~x6 | x0 | x3) & (~x0 | (x3 ? (x4 | ~x6) : (~x4 | x6)))));
  assign z494 = n5340 | ~n5344 | ~n5346 | (~n620 & ~n5343);
  assign n5340 = ~x0 & ((x7 & ~n5341) | (n540 & ~n5342));
  assign n5341 = (x1 | x2 | x3 | x4 | x5 | x6) & (~x6 | ((x3 | ((~x4 | x5 | ~x1 | ~x2) & (x1 | (x2 ? (x4 | x5) : ~x4)))) & (~x1 | ~x3 | (x2 ? (~x4 | ~x5) : (x4 | x5)))));
  assign n5342 = (~x4 | ~x5 | ~x1 | x3) & (x1 | x4 | ((x3 | ~x5) & (x2 | ~x3 | x5)));
  assign n5343 = x1 ? ((x2 | ((~x3 | x4 | x5) & (~x4 | ~x5 | x0 | x3))) & (x0 | x4 | ((x3 | x5) & (~x2 | ~x3 | ~x5)))) : ((~x5 | (~x0 ^ ~x3) | (x2 ^ x4)) & (~x4 | x5 | (x2 & (~x0 | x3))));
  assign n5344 = (~x6 | n5345) & (n1451 | n1957) & (n1019 | n1252);
  assign n5345 = (x3 | ~x4 | ~x5 | ~x0 | x1 | ~x2) & (x0 | ((x1 | x2 | ~x3 | ~x4 | ~x5) & (~x1 | ((~x4 | x5 | ~x2 | ~x3) & (x3 | x4 | ~x5)))));
  assign n5346 = (~n738 | n5348) & (x6 | n5347);
  assign n5347 = (x0 | ~x1 | ((x2 | ~x4 | (x3 ^ x5)) & (x4 | x5 | ~x2 | ~x3))) & (x1 | (x0 ? (x3 ? (x5 | (x2 ^ x4)) : (x4 | ~x5)) : ((~x4 | x5 | ~x2 | x3) & (x2 | ~x3 | x4 | ~x5))));
  assign n5348 = (~x6 | ~x7 | ((~x2 | ~x3 | x4 | x5) & (x2 | ~x4 | (~x3 & ~x5)))) & (x4 | x6 | x7 | (x3 ^ x5));
  assign z495 = ~n5355 | (x5 ? ~n5352 : (x0 ? ~n5351 : ~n5350));
  assign n5350 = x3 ? (x2 ? ((x6 | ~x7 | ~x1 | x4) & (x1 | ~x4 | (x6 ^ x7))) : ((x4 | ~x6 | ~x7) & (~x1 | ((~x6 | ~x7) & (x4 | x6 | x7))))) : ((x1 | ~x2 | x4 | x6 | ~x7) & (~x4 | (x1 ? (~x2 | (~x6 ^ x7)) : (x2 | (x6 ^ x7)))));
  assign n5351 = (x2 | ((x1 | x3 | x4 | x6 | x7) & (~x4 | (x6 ^ x7) | (~x1 ^ x3)))) & (x1 | x4 | ~x7 | ((x3 | ~x6) & (~x2 | ~x3 | x6)));
  assign n5352 = (x1 | n5353) & (x0 | ~x1 | n5354);
  assign n5353 = (x0 | ((~x2 | x3 | x4 | ~x6 | ~x7) & (x2 | ~x3 | ~x4 | x6 | x7))) & (x2 | x3 | ~x4 | ~x6 | x7) & (~x0 | (x2 ? ((x3 | ~x4 | x6 | x7) & (~x6 | ~x7 | ~x3 | x4)) : ((x6 | ~x7 | x3 | x4) & (~x4 | ~x6 | x7))));
  assign n5354 = (~x6 | ((x2 | ~x3 | x4 | x7) & (~x4 | (x2 ? (~x3 ^ x7) : (x3 | x7))))) & (x4 | x6 | (x2 ? (x3 | x7) : ~x7));
  assign n5355 = ~n5358 & ~n5359 & (x1 ? (x0 | n5357) : n5356);
  assign n5356 = (x5 | ((~x3 | ((x4 | ~x7 | ~x0 | x2) & (x0 | (x2 ? (x4 | ~x7) : (~x4 | x7))))) & (~x0 | x3 | x7 | (~x2 & ~x4)))) & (x0 | ~x5 | (x2 ? (x3 | x7) : (~x3 | ~x7)));
  assign n5357 = (x3 | x4 | x5 | x7) & (~x4 | ((~x5 | ~x7 | x2 | ~x3) & (~x2 | (x3 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n5358 = ~n906 & (x0 ? (x1 ? (~x4 & n1184) : n2895) : (x1 ? (x4 ? n1184 : n2895) : (~x4 & n1184)));
  assign n5359 = ~n1311 & ((x0 & x1 & ~x2 & ~x3 & x5) | (~x1 & ((x3 & x5 & ~x0 & x2) | ((x2 ^ x5) & (x0 ^ ~x3)))));
  assign z496 = ~n5366 | (x5 ? (x1 ? ~n5365 : ~n5364) : ~n5361);
  assign n5361 = (x0 | n5363) & (~n534 | ~n1967) & (n662 | n5362);
  assign n5362 = (x0 | ~x1 | x2 | ~x3 | ~x4) & (x1 | ((~x3 | x4 | x0 | x2) & (~x2 | (x0 ? (~x3 ^ ~x4) : (x3 | ~x4)))));
  assign n5363 = (x4 | (x1 ? ((~x6 | ~x7 | ~x2 | ~x3) & (x2 | x3 | x6 | x7)) : ((x2 | x3 | x6 | ~x7) & (~x6 | x7 | ~x2 | ~x3)))) & (~x3 | ~x4 | ~x6 | x7 | (~x1 ^ ~x2));
  assign n5364 = ((x2 ^ x7) | ((~x0 | (x3 ? (x4 | ~x6) : (~x4 | x6))) & (~x4 | ~x6 | x0 | ~x3))) & (~x4 | ((~x0 | ~x2 | x3 | ~x6 | x7) & (x0 | x2 | ~x3 | x6 | ~x7))) & (x0 | x2 | x3 | x4 | (~x6 ^ x7));
  assign n5365 = (x0 | ~x2 | ~x3 | ~x4 | ~x6 | x7) & (x3 | ((~x4 | ~x6 | ~x7 | ~x0 | x2) & ((~x6 ^ x7) | (x0 ? (x2 | x4) : (~x2 ^ x4)))));
  assign n5366 = (n1323 | n5369) & (x5 | n5368) & (~x5 | n5367);
  assign n5367 = x6 ? ((x0 | ~x1 | x2 | ~x3 | x4) & (x1 | ((~x3 | ~x4 | ~x0 | x2) & (x0 | (x2 ? (~x3 | x4) : (x3 | ~x4)))))) : (((x0 ? (x1 | ~x2) : (~x1 | x2)) | (~x3 ^ ~x4)) & (x0 | ((~x3 | x4 | ~x1 | ~x2) & (x1 | (x2 ? (x3 | ~x4) : (~x3 | x4))))));
  assign n5368 = ((x4 ^ x6) | (~x1 ^ x3) | (~x0 ^ x2)) & ((x0 ? (x1 | ~x2) : (~x1 | x2)) | (x3 ? (x4 | ~x6) : (~x4 | x6))) & (~x0 | x1 | x2 | x3 | x4 | ~x6) & (x0 | ((x1 | x2 | ~x4 | (~x3 ^ x6)) & (~x2 | ((~x4 | x6 | ~x1 | ~x3) & (x4 | ~x6 | x1 | x3)))));
  assign n5369 = (~x4 | ~x5 | ~x7 | x0 | ~x1 | ~x2) & (x4 | (x1 ? (x5 | x7) : (~x5 | ~x7)) | (~x0 ^ x2));
  assign z497 = (~x3 & ~n5371) | (x3 & ~n5372) | ~n5374 | (~n662 & ~n5373);
  assign n5371 = ((~x0 ^ x2) | (x1 ? (x4 ? (x5 | x7) : (~x5 | ~x7)) : (x7 | (~x4 ^ ~x5)))) & (x0 | ~x1 | x2 | x4 | ~x5 | x7) & (~x7 | ((x0 | ~x1 | x2 | ~x4 | ~x5) & (x1 | ((x4 | ~x5 | x0 | x2) & (~x2 | (x0 ? (~x4 ^ ~x5) : (~x4 | x5)))))));
  assign n5372 = ((~x5 ^ x7) | ((~x0 | x1 | ~x2 | ~x4) & (x0 | x4 | (~x1 ^ ~x2)))) & (~x0 | x1 | x2 | x4 | ~x5 | ~x7) & (x0 | ~x4 | ((x5 | x7 | x1 | ~x2) & (~x7 | (x1 ? (x2 ^ x5) : (x2 | ~x5)))));
  assign n5373 = ((x4 ^ x5) | (~x1 ^ x3) | (~x0 ^ x2)) & ((x0 ? (x1 | ~x2) : (~x1 | x2)) | (x3 ? (x4 | ~x5) : (~x4 | x5))) & (~x0 | x1 | x2 | x3 | x4 | ~x5) & (x0 | ((x1 | x2 | ~x4 | (~x3 ^ x5)) & (~x2 | ((~x4 | x5 | ~x1 | ~x3) & (x4 | ~x5 | x1 | x3)))));
  assign n5374 = (x2 & (x1 | n5379)) | (~x2 & ~n5375 & ~n5376 & n5378);
  assign n5375 = n1205 & ((x1 & x4 & ~x7 & (~x3 ^ x5)) | (~x1 & ~x3 & ~x4 & ~x5 & x7));
  assign n5376 = ~n5377 & (n732 | n669);
  assign n5377 = (~x1 | x4 | x5 | x6 | ~x7) & (x1 | ~x6 | x7 | (~x4 & x5));
  assign n5378 = (~n3098 | ~n1743) & (~n586 | (~n3262 & ~n1231));
  assign n5379 = (~x3 | ((x5 | ~x6 | x7 | ~x0 | x4) & (x0 | x6 | ~x7 | (x4 & ~x5)))) & (~x0 | x3 | ~x6 | x7 | (~x4 ^ x5));
  assign z498 = ~n5385 | (~x3 & (~n5382 | (~x0 & ~n5381)));
  assign n5381 = (x2 | x7 | (x1 ? ((x5 | x6) & (x4 | ~x5 | ~x6)) : (~x4 | x6))) & (x1 | ~x2 | ~x6 | ~x7 | (~x4 & x5));
  assign n5382 = n5384 & (n627 | n5383) & (~n534 | (~n3290 & ~n1163));
  assign n5383 = (~x2 | ~x6 | ~x7 | x0 | ~x1) & (~x0 | ((x1 | x6 | x7) & (~x1 | x2 | ~x6 | ~x7)));
  assign n5384 = ((~x4 ^ ~x5) | ((x0 | ~x1 | ~x2 | x6) & (~x0 | (x1 ? (x2 | x6) : (~x2 | ~x6))))) & (x0 | ~x5 | ((~x4 | ~x6 | ~x1 | x2) & (x1 | x4 | (~x2 ^ x6))));
  assign n5385 = (n620 | n5386) & (~x3 | (~n5387 & n5388));
  assign n5386 = x5 ? (x1 ? ((x3 | x4 | ~x0 | x2) & (x0 | (x2 ? (~x3 ^ ~x4) : (~x3 | x4)))) : ((x2 | ~x3 | ~x4) & (x0 | (x2 ? (~x3 | x4) : ~x4)))) : ((x0 | ((x2 | x3 | x4) & (~x1 | (x2 ? (~x3 | x4) : x3)))) & (~x3 | x4 | ~x0 | x2) & (x1 | ((x2 | ~x3 | x4) & (~x4 | ((~x2 | x3) & (~x0 | (~x2 & x3)))))));
  assign n5387 = ~n912 & ((x0 & ~x1 & x2 & ~x4 & x7) | (~x0 & x4 & ~x7 & (~x1 ^ ~x2)));
  assign n5388 = ~n3567 & ~n5389 & n5391 & (~n537 | ~n545 | n5390);
  assign n5389 = ~x1 & ~x4 & ((x2 & ~x6 & ~x7) | (x6 & x7 & ~x0 & ~x2));
  assign n5390 = x1 ? (~x2 ^ ~x5) : (x2 ^ ~x5);
  assign n5391 = (~x0 | x1 | x2 | x4 | ~x5 | ~x6) & (x0 | ~x4 | x5 | x6 | (~x1 ^ ~x2));
  assign z499 = n5394 | ~n5395 | ~n5399 | (~x3 & ~n5393);
  assign n5393 = (x4 | ~x7 | ~n750 | (~x5 ^ ~x6)) & (~n534 | ((~x6 | x7 | ~x4 | x5) & (x4 | (x5 ? (~x6 ^ ~x7) : (x6 | ~x7)))));
  assign n5394 = n664 & ((x5 & ~x6 & ~x7 & ~x3 & ~x4) | (x4 & ((~x3 & (x5 ? (~x6 & x7) : (x6 & ~x7))) | (x3 & x5 & x6 & x7))));
  assign n5395 = ~n3670 & ~n5396 & ~n5397 & (n5398 | (x1 & ~n539));
  assign n5396 = ~x0 & ~x5 & ~x7 & (x1 ? (x3 & ~x4) : (~x3 & x4));
  assign n5397 = ~n800 & ((~x4 & ~n910 & x0 & ~x3) | (~x0 & x1 & x3 & x4));
  assign n5398 = (x0 | x3 | x4 | ~x5 | ~x7) & (~x0 | ((x3 | ~x4 | ~x5 | ~x7) & (~x3 | x4 | x5 | x7)));
  assign n5399 = (n620 | n5400) & (x1 | n5401);
  assign n5400 = (~x3 | x4 | ~x5 | x0 | ~x1) & (x3 | ((~x4 | ~x5 | x0 | x1) & (x5 | (x0 ? (~x4 | (x1 ^ ~x2)) : (x4 | (x1 & x2))))));
  assign n5401 = x0 ? (~x3 | ((~x5 | (x4 ? (~x6 | x7) : (x6 | ~x7))) & (~x4 | x5 | (x6 ^ x7)))) : (x3 ? ((x4 | ~x5 | ~x6 | x7) & (x6 | ~x7 | ~x4 | x5) & ((~x4 ^ ~x5) | (x6 ^ x7))) : ((x4 | ~x5 | x6 | x7) & (~x6 | ~x7 | ~x4 | x5)));
  assign z500 = n5409 | ~n5410 | (x4 ? (n5407 | ~n5408) : ~n5403);
  assign n5403 = ~n5405 & ~n5406 & (x0 | n5404);
  assign n5404 = x5 ? ((x6 | ~x7 | (x1 & (x2 | x3))) & (~x1 | ~x6 | (~x2 & ~x3) | x7)) : (~x6 | x7 | (x1 & (x2 | x3)));
  assign n5405 = n534 & n544 & n708;
  assign n5406 = ~n662 & ((x0 & ~x2 & ~x3 & (~x1 ^ x5)) | ((x2 | x3) & (x0 ? (~x1 & x5) : (x1 & ~x5))));
  assign n5407 = ~n620 & ((x1 & ((~x0 & ~x5) | (~x3 & x5 & x0 & ~x2))) | (x0 & ~x1 & ((~x2 & ~x3 & ~x5) | (x5 & (x2 | x3)))));
  assign n5408 = ~n5405 & (x0 | ((~x1 | ~x5 | ~x6 | ~x7) & (x1 | (x5 ? (x6 | x7) : (~x6 | ~x7)))));
  assign n5409 = n651 & ((x1 & ~x3 & x4 & ~x5 & x6) | (~x1 & ((x5 & ~x6 & ~x3 & x4) | (x3 & ~x5 & (~x4 ^ x6)))));
  assign n5410 = (x6 | ((~x4 | ~x5 | x0 | ~x1) & (x5 | (x0 ? (x4 | (x1 ^ ~x2)) : (x1 | ~x4))))) & (x1 | ~x4 | ~x6 | (x0 ? (~x2 | x5) : ~x5));
  assign z501 = n5412 | n5414 | ~n5416 | (~x2 & ~n5413);
  assign n5412 = x7 & ((~n846 & ~n4690) | (~x0 & ~x1 & n1121));
  assign n5413 = (~x0 | ~x1 | ~x3 | x4 | x5 | x7) & (x3 | ~x5 | (x0 ? (x1 | (x4 ^ x7)) : (~x1 | (~x4 ^ x7))));
  assign n5414 = n540 & n1558 & (n5415 | (~x1 & (n3453 | ~n2113)));
  assign n5415 = ~x4 & ~x3 & x1 & ~x2;
  assign n5416 = n5418 & (n800 | n5417);
  assign n5417 = (x3 | ~x4 | x6 | ~x0 | x1 | x2) & (x0 | ~x6 | (x1 & (x2 | x3 | x4)));
  assign n5418 = ((~x2 & ~x3) | ((~x5 | x7 | x0 | ~x1) & (~x0 | x1 | (x5 ^ x7)))) & (~x0 | ~x1 | x2 | x3 | (x5 ^ x7));
  assign z138 = z004;
  assign z215 = ~n2074 | (~x3 & (x6 ? (~x7 & ~n577) : ~n2073));
  assign z254 = z037;
  assign z339 = z032;
  assign z340 = z033;
  assign z363 = n1673 | ~n1675 | (x5 ? (x7 ? ~n1671 : ~n1672) : (x7 ? ~n1672 : ~n1671));
  assign z364 = n1683 | ~n1686 | ~n1691 | ~n1694 | (~n620 & ~n1685);
  assign z420 = z033;
  assign z421 = z034;
  assign z422 = z034;
  assign z423 = z034;
  assign z424 = z034;
  assign z425 = z034;
  assign z426 = z034;
  assign z427 = z034;
  assign z428 = z034;
  assign z502 = z419;
  assign z503 = z033;
  assign z504 = z034;
  assign z505 = z034;
  assign z506 = z034;
  assign z507 = z034;
  assign z508 = z034;
  assign z509 = z034;
  assign z510 = z034;
  assign z511 = z034;
  assign z512 = z034;
endmodule


