// Benchmark "X_26" written by ABC on Fri Jun 02 03:25:15 2023

module X_76 ( 
    x0, x1, x2, x3, x4, x5,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11  );
  input  x0, x1, x2, x3, x4, x5;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11;
  assign z00 = 1'b0;
  assign z01 = 1'b0;
  assign z02 = 1'b0;
  assign z03 = 1'b0;
  assign z04 = 1'b0;
  assign z05 = 1'b0;
  assign z06 = x0;
  assign z07 = x1;
  assign z08 = x2;
  assign z09 = x3;
  assign z10 = x4;
  assign z11 = x5;
endmodule


