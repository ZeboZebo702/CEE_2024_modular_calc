// Benchmark "X_5" written by ABC on Wed Jun 07 00:27:44 2023

module X_41 ( 
    x0, x1, x2, x3, x4, x5,
    z0, z1, z2, z3, z4, z5, z6, z7  );
  input  x0, x1, x2, x3, x4, x5;
  output z0, z1, z2, z3, z4, z5, z6, z7;
  assign z0 = 1'b0;
  assign z1 = 1'b0;
  assign z2 = x0;
  assign z3 = x1;
  assign z4 = x2;
  assign z5 = x3;
  assign z6 = x4;
  assign z7 = x5;
endmodule


