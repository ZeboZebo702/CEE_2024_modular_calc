module x_100_mod_4051(
    input [100:1] X,
    output [12:1] R
    );

wire [12:1] r1,r2,r3,r4,r5,r6,r7,r8,r9,r10,r11,r12,r13,r14,r15,r16;
/*wire [14:1] R_temp_1;
wire [14:1] R_temp_2;
wire [14:1] R_temp_3;
wire [14:1] R_temp_4;

wire [13:1] R_temp_5;
wire [13:1] R_temp_6;
wire [13:1] R_temp_7;

wire [12:1] R_temp_8;
wire [12:1] R_temp_9;

wire [12:1] R_temp_10;

wire [12:1] R_temp_11;
wire [12:1] R_temp_12;

wire [13:1] R_temp_13;

reg [12:1]  R_temp;
*/
X_2 label2 (.x0(X[12]),.x1(X[11]),.x2(X[10]),.x3(X[9]),.x4(X[8]),.x5(X[7]),
.z00(r1[12]),.z01(r1[11]),.z02(r1[10]),.z03(r1[9]),.z04(r1[8]),.z05(r1[7]),.z06(r1[6]),.z07(r1[5]),.z08(r1[4]),.z09(r1[3]),.z10(r1[2]),.z11(r1[1]));

X_3 label3 (.x0(X[18]),.x1(X[17]),.x2(X[16]),.x3(X[15]),.x4(X[14]),.x5(X[13]),
.z00(r2[12]),.z01(r2[11]),.z02(r2[10]),.z03(r2[9]),.z04(r2[8]),.z05(r2[7]),.z06(r2[6]),.z07(r2[5]),.z08(r2[4]),.z09(r2[3]),.z10(r2[2]),.z11(r2[1]));

X_4 label4 (.x0(X[24]),.x1(X[23]),.x2(X[22]),.x3(X[21]),.x4(X[20]),.x5(X[19]),
.z00(r3[12]),.z01(r3[11]),.z02(r3[10]),.z03(r3[9]),.z04(r3[8]),.z05(r3[7]),.z06(r3[6]),.z07(r3[5]),.z08(r3[4]),.z09(r3[3]),.z10(r3[2]),.z11(r3[1]));

X_5 label5 (.x0(X[30]),.x1(X[29]),.x2(X[28]),.x3(X[27]),.x4(X[26]),.x5(X[25]),
.z00(r4[12]),.z01(r4[11]),.z02(r4[10]),.z03(r4[9]),.z04(r4[8]),.z05(r4[7]),.z06(r4[6]),.z07(r4[5]),.z08(r4[4]),.z09(r4[3]),.z10(r4[2]),.z11(r4[1]));

X_6 label6 (.x0(X[36]),.x1(X[35]),.x2(X[34]),.x3(X[33]),.x4(X[32]),.x5(X[31]),
.z00(r5[12]),.z01(r5[11]),.z02(r5[10]),.z03(r5[9]),.z04(r5[8]),.z05(r5[7]),.z06(r5[6]),.z07(r5[5]),.z08(r5[4]),.z09(r5[3]),.z10(r5[2]),.z11(r5[1]));

X_7 label7 (.x0(X[42]),.x1(X[41]),.x2(X[40]),.x3(X[39]),.x4(X[38]),.x5(X[37]),
.z00(r6[12]),.z01(r6[11]),.z02(r6[10]),.z03(r6[9]),.z04(r6[8]),.z05(r6[7]),.z06(r6[6]),.z07(r6[5]),.z08(r6[4]),.z09(r6[3]),.z10(r6[2]),.z11(r6[1]));

X_8 label8 (.x0(X[48]),.x1(X[47]),.x2(X[46]),.x3(X[45]),.x4(X[44]),.x5(X[43]),
.z00(r7[12]),.z01(r7[11]),.z02(r7[10]),.z03(r7[9]),.z04(r7[8]),.z05(r7[7]),.z06(r7[6]),.z07(r7[5]),.z08(r7[4]),.z09(r7[3]),.z10(r7[2]),.z11(r7[1]));

X_9 label9 (.x0(X[54]),.x1(X[53]),.x2(X[52]),.x3(X[51]),.x4(X[50]),.x5(X[49]),
.z00(r8[12]),.z01(r8[11]),.z02(r8[10]),.z03(r8[9]),.z04(r8[8]),.z05(r8[7]),.z06(r8[6]),.z07(r8[5]),.z08(r8[4]),.z09(r8[3]),.z10(r8[2]),.z11(r8[1]));

X_10 label10 (.x0(X[60]),.x1(X[59]),.x2(X[58]),.x3(X[57]),.x4(X[56]),.x5(X[55]),
.z00(r9[12]),.z01(r9[11]),.z02(r9[10]),.z03(r9[9]),.z04(r9[8]),.z05(r9[7]),.z06(r9[6]),.z07(r9[5]),.z08(r9[4]),.z09(r9[3]),.z10(r9[2]),.z11(r9[1]));

X_11 label11 (.x0(X[66]),.x1(X[65]),.x2(X[64]),.x3(X[63]),.x4(X[62]),.x5(X[61]),
.z00(r10[12]),.z01(r10[11]),.z02(r10[10]),.z03(r10[9]),.z04(r10[8]),.z05(r10[7]),.z06(r10[6]),.z07(r10[5]),.z08(r10[4]),.z09(r10[3]),.z10(r10[2]),.z11(r10[1]));

X_12 label12 (.x0(X[72]),.x1(X[71]),.x2(X[70]),.x3(X[69]),.x4(X[68]),.x5(X[67]),
.z00(r11[12]),.z01(r11[11]),.z02(r11[10]),.z03(r11[9]),.z04(r11[8]),.z05(r11[7]),.z06(r11[6]),.z07(r11[5]),.z08(r11[4]),.z09(r11[3]),.z10(r11[2]),.z11(r11[1]));

X_13 label13 (.x0(X[78]),.x1(X[77]),.x2(X[76]),.x3(X[75]),.x4(X[74]),.x5(X[73]),
.z00(r12[12]),.z01(r12[11]),.z02(r12[10]),.z03(r12[9]),.z04(r12[8]),.z05(r12[7]),.z06(r12[6]),.z07(r12[5]),.z08(r12[4]),.z09(r12[3]),.z10(r12[2]),.z11(r12[1]));

X_14 label14 (.x0(X[84]),.x1(X[83]),.x2(X[82]),.x3(X[81]),.x4(X[80]),.x5(X[79]),
.z00(r13[12]),.z01(r13[11]),.z02(r13[10]),.z03(r13[9]),.z04(r13[8]),.z05(r13[7]),.z06(r13[6]),.z07(r13[5]),.z08(r13[4]),.z09(r13[3]),.z10(r13[2]),.z11(r13[1]));

X_15 label15 (.x0(X[90]),.x1(X[89]),.x2(X[88]),.x3(X[87]),.x4(X[86]),.x5(X[85]),
.z00(r14[12]),.z01(r14[11]),.z02(r14[10]),.z03(r14[9]),.z04(r14[8]),.z05(r14[7]),.z06(r14[6]),.z07(r14[5]),.z08(r14[4]),.z09(r14[3]),.z10(r14[2]),.z11(r14[1]));

X_16 label16 (.x0(X[96]),.x1(X[95]),.x2(X[94]),.x3(X[93]),.x4(X[92]),.x5(X[91]),
.z00(r15[12]),.z01(r15[11]),.z02(r15[10]),.z03(r15[9]),.z04(r15[8]),.z05(r15[7]),.z06(r15[6]),.z07(r15[5]),.z08(r15[4]),.z09(r15[3]),.z10(r15[2]),.z11(r15[1]));

X_17 label17 (.x0(X[100]),.x1(X[99]),.x2(X[98]),.x3(X[97]),
.z00(r16[12]),.z01(r16[11]),.z02(r16[10]),.z03(r16[9]),.z04(r16[8]),.z05(r16[7]),.z06(r16[6]),.z07(r16[5]),.z08(r16[4]),.z09(r16[3]),.z10(r16[2]),.z11(r16[1]));

wire [14:1] R_temp_1;
wire [14:1] R_temp_2;
wire [14:1] R_temp_3;
wire [14:1] R_temp_4;
wire [14:1] R_temp_5;

assign R_temp_1 = r1 + r2 + r3;
assign R_temp_2 = r4 + r5 + r6;
assign R_temp_3 = r7 + r8 + r9;
assign R_temp_4 = r10 + r11 + r12;
assign R_temp_5 = r13 + r14 + r15;

wire [15:1] R_temp_6;
wire [15:1] R_temp_7;

assign R_temp_6 = r16 + R_temp_1 + R_temp_2;
assign R_temp_7 = R_temp_3 + R_temp_4 + R_temp_5;

wire [13:1] R_temp_8;

assign R_temp_8 = R_temp_6 [6:1] + 64* R_temp_6 [12:7] + 45* R_temp_6 [15:13] + 
            R_temp_7 [6:1] + 64* R_temp_7 [12:7] + 45* R_temp_7 [15:13] + X[6:1];


/*assign R_temp_1 = r1 + r2 + r3 + r16;

assign R_temp_2 = r4 + r5 + r6 + r7;

assign R_temp_3 = r8 + r9 + r10 + r11;

assign R_temp_4 = r12 + r13 + r14 + r15;


assign R_temp_5 = R_temp_1 [6:1] + 64 * R_temp_1 [12:7] + 45 * R_temp_1 [14:13] + 64 * R_temp_2 [12:7];

assign R_temp_6 = R_temp_2 [6:1] + 45 * R_temp_2 [14:13] + R_temp_3 [6:1] + 64 * R_temp_3 [12:7];

assign R_temp_7 = R_temp_4 [6:1] + 45 * R_temp_3 [14:13] + 64 * R_temp_4 [12:7] + 45 * R_temp_4 [14:13];


assign R_temp_8 = R_temp_5 [6:1] + 64 * R_temp_5 [12:7] + 45 * R_temp_5 [13];

assign R_temp_9 = R_temp_6 [6:1] + 64 * R_temp_7 [12:7] + 45 * R_temp_6 [13];

assign R_temp_10 = 64 * R_temp_6 [12:7] + R_temp_7 [6:1] + 45 * R_temp_7 [13];


assign R_temp_11 = X[6:1] + R_temp_8 [6:1] + 64 * R_temp_8 [12:7];

assign R_temp_12 = R_temp_9 [6:1] + 64 * R_temp_9 [12:7] + 45 * R_temp_8 [13] + 45 * R_temp_9 [13];


assign R_temp_13 = R_temp_11 [6:1] + R_temp_12 [6:1] + 64 * R_temp_11 [12:7] + 64 * R_temp_12 [12:7];

*/

reg [12:1]  R_temp;

always @(R_temp_8)
begin
  if (R_temp_8 >= 12'b111111010011  )
    R_temp <= R_temp_8 - 12'b111111010011;
  else
    R_temp <= R_temp_8;
end

assign R = R_temp;

endmodule