module x_300_mod_2011(
    input [300:1] X,
    output [11:1] R
    );

wire [11:1] r1,r2,r3,r4,r5,r6,r7,r8,r9,r10,r11,r12,r13,r14,r15,r16,r17,
        r18,r19,r20,r21,r22,r23,r24,r25,r26,r27,r28,r29,r30,r31,r32,r33,
	r34,r35,r36,r37,r38,r39,r40,r41,r42,r43,r44,r45,r46,r47,r48,r49;

X_2 label2 (.x0(X[12]),.x1(X[11]),.x2(X[10]),.x3(X[9]),.x4(X[8]),.x5(X[7]),
.z00(r1[11]),.z01(r1[10]),.z02(r1[9]),.z03(r1[8]),.z04(r1[7]),.z05(r1[6]),.z06(r1[5]),.z07(r1[4]),.z08(r1[3]),.z09(r1[2]),.z10(r1[1]));

X_3 label3 (.x0(X[18]),.x1(X[17]),.x2(X[16]),.x3(X[15]),.x4(X[14]),.x5(X[13]),
.z00(r2[11]),.z01(r2[10]),.z02(r2[9]),.z03(r2[8]),.z04(r2[7]),.z05(r2[6]),.z06(r2[5]),.z07(r2[4]),.z08(r2[3]),.z09(r2[2]),.z10(r2[1]));

X_4 label4 (.x0(X[24]),.x1(X[23]),.x2(X[22]),.x3(X[21]),.x4(X[20]),.x5(X[19]),
.z00(r3[11]),.z01(r3[10]),.z02(r3[9]),.z03(r3[8]),.z04(r3[7]),.z05(r3[6]),.z06(r3[5]),.z07(r3[4]),.z08(r3[3]),.z09(r3[2]),.z10(r3[1]));

X_5 label5 (.x0(X[30]),.x1(X[29]),.x2(X[28]),.x3(X[27]),.x4(X[26]),.x5(X[25]),
.z00(r4[11]),.z01(r4[10]),.z02(r4[9]),.z03(r4[8]),.z04(r4[7]),.z05(r4[6]),.z06(r4[5]),.z07(r4[4]),.z08(r4[3]),.z09(r4[2]),.z10(r4[1]));

X_6 label6 (.x0(X[36]),.x1(X[35]),.x2(X[34]),.x3(X[33]),.x4(X[32]),.x5(X[31]),
.z00(r5[11]),.z01(r5[10]),.z02(r5[9]),.z03(r5[8]),.z04(r5[7]),.z05(r5[6]),.z06(r5[5]),.z07(r5[4]),.z08(r5[3]),.z09(r5[2]),.z10(r5[1]));

X_7 label7 (.x0(X[42]),.x1(X[41]),.x2(X[40]),.x3(X[39]),.x4(X[38]),.x5(X[37]),
.z00(r6[11]),.z01(r6[10]),.z02(r6[9]),.z03(r6[8]),.z04(r6[7]),.z05(r6[6]),.z06(r6[5]),.z07(r6[4]),.z08(r6[3]),.z09(r6[2]),.z10(r6[1]));

X_8 label8 (.x0(X[48]),.x1(X[47]),.x2(X[46]),.x3(X[45]),.x4(X[44]),.x5(X[43]),
.z00(r7[11]),.z01(r7[10]),.z02(r7[9]),.z03(r7[8]),.z04(r7[7]),.z05(r7[6]),.z06(r7[5]),.z07(r7[4]),.z08(r7[3]),.z09(r7[2]),.z10(r7[1]));

X_9 label9 (.x0(X[54]),.x1(X[53]),.x2(X[52]),.x3(X[51]),.x4(X[50]),.x5(X[49]),
.z00(r8[11]),.z01(r8[10]),.z02(r8[9]),.z03(r8[8]),.z04(r8[7]),.z05(r8[6]),.z06(r8[5]),.z07(r8[4]),.z08(r8[3]),.z09(r8[2]),.z10(r8[1]));

X_10 label10 (.x0(X[60]),.x1(X[59]),.x2(X[58]),.x3(X[57]),.x4(X[56]),.x5(X[55]),
.z00(r9[11]),.z01(r9[10]),.z02(r9[9]),.z03(r9[8]),.z04(r9[7]),.z05(r9[6]),.z06(r9[5]),.z07(r9[4]),.z08(r9[3]),.z09(r9[2]),.z10(r9[1]));

X_11 label11 (.x0(X[66]),.x1(X[65]),.x2(X[64]),.x3(X[63]),.x4(X[62]),.x5(X[61]),
.z00(r10[11]),.z01(r10[10]),.z02(r10[9]),.z03(r10[8]),.z04(r10[7]),.z05(r10[6]),.z06(r10[5]),.z07(r10[4]),.z08(r10[3]),.z09(r10[2]),.z10(r10[1]));

X_12 label12 (.x0(X[72]),.x1(X[71]),.x2(X[70]),.x3(X[69]),.x4(X[68]),.x5(X[67]),
.z00(r11[11]),.z01(r11[10]),.z02(r11[9]),.z03(r11[8]),.z04(r11[7]),.z05(r11[6]),.z06(r11[5]),.z07(r11[4]),.z08(r11[3]),.z09(r11[2]),.z10(r11[1]));

X_13 label13 (.x0(X[78]),.x1(X[77]),.x2(X[76]),.x3(X[75]),.x4(X[74]),.x5(X[73]),
.z00(r12[11]),.z01(r12[10]),.z02(r12[9]),.z03(r12[8]),.z04(r12[7]),.z05(r12[6]),.z06(r12[5]),.z07(r12[4]),.z08(r12[3]),.z09(r12[2]),.z10(r12[1]));

X_14 label14 (.x0(X[84]),.x1(X[83]),.x2(X[82]),.x3(X[81]),.x4(X[80]),.x5(X[79]),
.z00(r13[11]),.z01(r13[10]),.z02(r13[9]),.z03(r13[8]),.z04(r13[7]),.z05(r13[6]),.z06(r13[5]),.z07(r13[4]),.z08(r13[3]),.z09(r13[2]),.z10(r13[1]));

X_15 label15 (.x0(X[90]),.x1(X[89]),.x2(X[88]),.x3(X[87]),.x4(X[86]),.x5(X[85]),
.z00(r14[11]),.z01(r14[10]),.z02(r14[9]),.z03(r14[8]),.z04(r14[7]),.z05(r14[6]),.z06(r14[5]),.z07(r14[4]),.z08(r14[3]),.z09(r14[2]),.z10(r14[1]));

X_16 label16 (.x0(X[96]),.x1(X[95]),.x2(X[94]),.x3(X[93]),.x4(X[92]),.x5(X[91]),
.z00(r15[11]),.z01(r15[10]),.z02(r15[9]),.z03(r15[8]),.z04(r15[7]),.z05(r15[6]),.z06(r15[5]),.z07(r15[4]),.z08(r15[3]),.z09(r15[2]),.z10(r15[1]));

X_17 label17 (.x0(X[102]),.x1(X[101]),.x2(X[100]),.x3(X[99]),.x4(X[98]),.x5(X[97]),
.z00(r16[11]),.z01(r16[10]),.z02(r16[9]),.z03(r16[8]),.z04(r16[7]),.z05(r16[6]),.z06(r16[5]),.z07(r16[4]),.z08(r16[3]),.z09(r16[2]),.z10(r16[1]));

X_18 label18 (.x0(X[108]),.x1(X[107]),.x2(X[106]),.x3(X[105]),.x4(X[104]),.x5(X[103]),
.z00(r17[11]),.z01(r17[10]),.z02(r17[9]),.z03(r17[8]),.z04(r17[7]),.z05(r17[6]),.z06(r17[5]),.z07(r17[4]),.z08(r17[3]),.z09(r17[2]),.z10(r17[1]));

X_19 label19 (.x0(X[114]),.x1(X[113]),.x2(X[112]),.x3(X[111]),.x4(X[110]),.x5(X[109]),
.z00(r18[11]),.z01(r18[10]),.z02(r18[9]),.z03(r18[8]),.z04(r18[7]),.z05(r18[6]),.z06(r18[5]),.z07(r18[4]),.z08(r18[3]),.z09(r18[2]),.z10(r18[1]));

X_20 label20 (.x0(X[120]),.x1(X[119]),.x2(X[118]),.x3(X[117]),.x4(X[116]),.x5(X[115]),
.z00(r19[11]),.z01(r19[10]),.z02(r19[9]),.z03(r19[8]),.z04(r19[7]),.z05(r19[6]),.z06(r19[5]),.z07(r19[4]),.z08(r19[3]),.z09(r19[2]),.z10(r19[1]));

X_21 label21 (.x0(X[126]),.x1(X[125]),.x2(X[124]),.x3(X[123]),.x4(X[122]),.x5(X[121]),
.z00(r20[11]),.z01(r20[10]),.z02(r20[9]),.z03(r20[8]),.z04(r20[7]),.z05(r20[6]),.z06(r20[5]),.z07(r20[4]),.z08(r20[3]),.z09(r20[2]),.z10(r20[1]));

X_22 label22 (.x0(X[132]),.x1(X[131]),.x2(X[130]),.x3(X[129]),.x4(X[128]),.x5(X[127]),
.z00(r21[11]),.z01(r21[10]),.z02(r21[9]),.z03(r21[8]),.z04(r21[7]),.z05(r21[6]),.z06(r21[5]),.z07(r21[4]),.z08(r21[3]),.z09(r21[2]),.z10(r21[1]));

X_23 label23 (.x0(X[138]),.x1(X[137]),.x2(X[136]),.x3(X[135]),.x4(X[134]),.x5(X[133]),
.z00(r22[11]),.z01(r22[10]),.z02(r22[9]),.z03(r22[8]),.z04(r22[7]),.z05(r22[6]),.z06(r22[5]),.z07(r22[4]),.z08(r22[3]),.z09(r22[2]),.z10(r22[1]));

X_24 label24 (.x0(X[144]),.x1(X[143]),.x2(X[142]),.x3(X[141]),.x4(X[140]),.x5(X[139]),
.z00(r23[11]),.z01(r23[10]),.z02(r23[9]),.z03(r23[8]),.z04(r23[7]),.z05(r23[6]),.z06(r23[5]),.z07(r23[4]),.z08(r23[3]),.z09(r23[2]),.z10(r23[1]));

X_25 label25 (.x0(X[150]),.x1(X[149]),.x2(X[148]),.x3(X[147]),.x4(X[146]),.x5(X[145]),
.z00(r24[11]),.z01(r24[10]),.z02(r24[9]),.z03(r24[8]),.z04(r24[7]),.z05(r24[6]),.z06(r24[5]),.z07(r24[4]),.z08(r24[3]),.z09(r24[2]),.z10(r24[1]));

X_26 label26 (.x0(X[156]),.x1(X[155]),.x2(X[154]),.x3(X[153]),.x4(X[152]),.x5(X[151]),
.z00(r25[11]),.z01(r25[10]),.z02(r25[9]),.z03(r25[8]),.z04(r25[7]),.z05(r25[6]),.z06(r25[5]),.z07(r25[4]),.z08(r25[3]),.z09(r25[2]),.z10(r25[1]));

X_27 label27 (.x0(X[162]),.x1(X[161]),.x2(X[160]),.x3(X[159]),.x4(X[158]),.x5(X[157]),
.z00(r26[11]),.z01(r26[10]),.z02(r26[9]),.z03(r26[8]),.z04(r26[7]),.z05(r26[6]),.z06(r26[5]),.z07(r26[4]),.z08(r26[3]),.z09(r26[2]),.z10(r26[1]));

X_28 label28 (.x0(X[168]),.x1(X[167]),.x2(X[166]),.x3(X[165]),.x4(X[164]),.x5(X[163]),
.z00(r27[11]),.z01(r27[10]),.z02(r27[9]),.z03(r27[8]),.z04(r27[7]),.z05(r27[6]),.z06(r27[5]),.z07(r27[4]),.z08(r27[3]),.z09(r27[2]),.z10(r27[1]));

X_29 label29 (.x0(X[174]),.x1(X[173]),.x2(X[172]),.x3(X[171]),.x4(X[170]),.x5(X[169]),
.z00(r28[11]),.z01(r28[10]),.z02(r28[9]),.z03(r28[8]),.z04(r28[7]),.z05(r28[6]),.z06(r28[5]),.z07(r28[4]),.z08(r28[3]),.z09(r28[2]),.z10(r28[1]));

X_30 label30 (.x0(X[180]),.x1(X[179]),.x2(X[178]),.x3(X[177]),.x4(X[176]),.x5(X[175]),
.z00(r29[11]),.z01(r29[10]),.z02(r29[9]),.z03(r29[8]),.z04(r29[7]),.z05(r29[6]),.z06(r29[5]),.z07(r29[4]),.z08(r29[3]),.z09(r29[2]),.z10(r29[1]));

X_31 label31 (.x0(X[186]),.x1(X[185]),.x2(X[184]),.x3(X[183]),.x4(X[182]),.x5(X[181]),
.z00(r30[11]),.z01(r30[10]),.z02(r30[9]),.z03(r30[8]),.z04(r30[7]),.z05(r30[6]),.z06(r30[5]),.z07(r30[4]),.z08(r30[3]),.z09(r30[2]),.z10(r30[1]));

X_32 label32 (.x0(X[192]),.x1(X[191]),.x2(X[190]),.x3(X[189]),.x4(X[188]),.x5(X[187]),
.z00(r31[11]),.z01(r31[10]),.z02(r31[9]),.z03(r31[8]),.z04(r31[7]),.z05(r31[6]),.z06(r31[5]),.z07(r31[4]),.z08(r31[3]),.z09(r31[2]),.z10(r31[1]));

X_33 label33 (.x0(X[198]),.x1(X[197]),.x2(X[196]),.x3(X[195]),.x4(X[194]),.x5(X[193]),
.z00(r32[11]),.z01(r32[10]),.z02(r32[9]),.z03(r32[8]),.z04(r32[7]),.z05(r32[6]),.z06(r32[5]),.z07(r32[4]),.z08(r32[3]),.z09(r32[2]),.z10(r32[1]));

X_34 label34 (.x0(X[204]),.x1(X[203]),.x2(X[202]),.x3(X[201]),.x4(X[200]),.x5(X[199]),
.z00(r33[11]),.z01(r33[10]),.z02(r33[9]),.z03(r33[8]),.z04(r33[7]),.z05(r33[6]),.z06(r33[5]),.z07(r33[4]),.z08(r33[3]),.z09(r33[2]),.z10(r33[1]));

X_35 label35 (.x0(X[210]),.x1(X[209]),.x2(X[208]),.x3(X[207]),.x4(X[206]),.x5(X[205]),
.z00(r34[11]),.z01(r34[10]),.z02(r34[9]),.z03(r34[8]),.z04(r34[7]),.z05(r34[6]),.z06(r34[5]),.z07(r34[4]),.z08(r34[3]),.z09(r34[2]),.z10(r34[1]));

X_36 label36 (.x0(X[216]),.x1(X[215]),.x2(X[214]),.x3(X[213]),.x4(X[212]),.x5(X[211]),
.z00(r35[11]),.z01(r35[10]),.z02(r35[9]),.z03(r35[8]),.z04(r35[7]),.z05(r35[6]),.z06(r35[5]),.z07(r35[4]),.z08(r35[3]),.z09(r35[2]),.z10(r35[1]));

X_37 label37 (.x0(X[222]),.x1(X[221]),.x2(X[220]),.x3(X[219]),.x4(X[218]),.x5(X[217]),
.z00(r36[11]),.z01(r36[10]),.z02(r36[9]),.z03(r36[8]),.z04(r36[7]),.z05(r36[6]),.z06(r36[5]),.z07(r36[4]),.z08(r36[3]),.z09(r36[2]),.z10(r36[1]));

X_38 label38 (.x0(X[228]),.x1(X[227]),.x2(X[226]),.x3(X[225]),.x4(X[224]),.x5(X[223]),
.z00(r37[11]),.z01(r37[10]),.z02(r37[9]),.z03(r37[8]),.z04(r37[7]),.z05(r37[6]),.z06(r37[5]),.z07(r37[4]),.z08(r37[3]),.z09(r37[2]),.z10(r37[1]));

X_39 label39 (.x0(X[234]),.x1(X[233]),.x2(X[232]),.x3(X[231]),.x4(X[230]),.x5(X[229]),
.z00(r38[11]),.z01(r38[10]),.z02(r38[9]),.z03(r38[8]),.z04(r38[7]),.z05(r38[6]),.z06(r38[5]),.z07(r38[4]),.z08(r38[3]),.z09(r38[2]),.z10(r38[1]));

X_40 label40 (.x0(X[240]),.x1(X[239]),.x2(X[238]),.x3(X[237]),.x4(X[236]),.x5(X[235]),
.z00(r39[11]),.z01(r39[10]),.z02(r39[9]),.z03(r39[8]),.z04(r39[7]),.z05(r39[6]),.z06(r39[5]),.z07(r39[4]),.z08(r39[3]),.z09(r39[2]),.z10(r39[1]));

X_41 label41 (.x0(X[246]),.x1(X[245]),.x2(X[244]),.x3(X[243]),.x4(X[242]),.x5(X[241]),
.z00(r40[11]),.z01(r40[10]),.z02(r40[9]),.z03(r40[8]),.z04(r40[7]),.z05(r40[6]),.z06(r40[5]),.z07(r40[4]),.z08(r40[3]),.z09(r40[2]),.z10(r40[1]));

X_42 label42 (.x0(X[252]),.x1(X[251]),.x2(X[250]),.x3(X[249]),.x4(X[248]),.x5(X[247]),
.z00(r41[11]),.z01(r41[10]),.z02(r41[9]),.z03(r41[8]),.z04(r41[7]),.z05(r41[6]),.z06(r41[5]),.z07(r41[4]),.z08(r41[3]),.z09(r41[2]),.z10(r41[1]));

X_43 label43 (.x0(X[258]),.x1(X[257]),.x2(X[256]),.x3(X[255]),.x4(X[254]),.x5(X[253]),
.z00(r42[11]),.z01(r42[10]),.z02(r42[9]),.z03(r42[8]),.z04(r42[7]),.z05(r42[6]),.z06(r42[5]),.z07(r42[4]),.z08(r42[3]),.z09(r42[2]),.z10(r42[1]));

X_44 label44 (.x0(X[264]),.x1(X[263]),.x2(X[262]),.x3(X[261]),.x4(X[260]),.x5(X[259]),
.z00(r43[11]),.z01(r43[10]),.z02(r43[9]),.z03(r43[8]),.z04(r43[7]),.z05(r43[6]),.z06(r43[5]),.z07(r43[4]),.z08(r43[3]),.z09(r43[2]),.z10(r43[1]));

X_45 label45 (.x0(X[270]),.x1(X[269]),.x2(X[268]),.x3(X[267]),.x4(X[266]),.x5(X[265]),
.z00(r44[11]),.z01(r44[10]),.z02(r44[9]),.z03(r44[8]),.z04(r44[7]),.z05(r44[6]),.z06(r44[5]),.z07(r44[4]),.z08(r44[3]),.z09(r44[2]),.z10(r44[1]));

X_46 label46 (.x0(X[276]),.x1(X[275]),.x2(X[274]),.x3(X[273]),.x4(X[272]),.x5(X[271]),
.z00(r45[11]),.z01(r45[10]),.z02(r45[9]),.z03(r45[8]),.z04(r45[7]),.z05(r45[6]),.z06(r45[5]),.z07(r45[4]),.z08(r45[3]),.z09(r45[2]),.z10(r45[1]));

X_47 label47 (.x0(X[282]),.x1(X[281]),.x2(X[280]),.x3(X[279]),.x4(X[278]),.x5(X[277]),
.z00(r46[11]),.z01(r46[10]),.z02(r46[9]),.z03(r46[8]),.z04(r46[7]),.z05(r46[6]),.z06(r46[5]),.z07(r46[4]),.z08(r46[3]),.z09(r46[2]),.z10(r46[1]));

X_48 label48 (.x0(X[288]),.x1(X[287]),.x2(X[286]),.x3(X[285]),.x4(X[284]),.x5(X[283]),
.z00(r47[11]),.z01(r47[10]),.z02(r47[9]),.z03(r47[8]),.z04(r47[7]),.z05(r47[6]),.z06(r47[5]),.z07(r47[4]),.z08(r47[3]),.z09(r47[2]),.z10(r47[1]));

X_49 label49 (.x0(X[294]),.x1(X[293]),.x2(X[292]),.x3(X[291]),.x4(X[290]),.x5(X[289]),
.z00(r48[11]),.z01(r48[10]),.z02(r48[9]),.z03(r48[8]),.z04(r48[7]),.z05(r48[6]),.z06(r48[5]),.z07(r48[4]),.z08(r48[3]),.z09(r48[2]),.z10(r48[1]));

X_50 label50 (.x0(X[300]),.x1(X[299]),.x2(X[298]),.x3(X[297]),.x4(X[296]),.x5(X[295]),
.z00(r49[11]),.z01(r49[10]),.z02(r49[9]),.z03(r49[8]),.z04(r49[7]),.z05(r49[6]),.z06(r49[5]),.z07(r49[4]),.z08(r49[3]),.z09(r49[2]),.z10(r49[1]));

wire [13:1] R_temp_1,R_temp_2,R_temp_3,R_temp_4,R_temp_5,R_temp_6,R_temp_7,R_temp_8,R_temp_9,R_temp_10,R_temp_11,
	R_temp_12,R_temp_13,R_temp_14,R_temp_15,R_temp_16;

assign R_temp_1 = r1 + r2 + r3;
assign R_temp_2 = r4 + r5 + r6;
assign R_temp_3 = r7 + r8 + r9;
assign R_temp_4 = r10 + r11 + r12;
assign R_temp_5 = r13 + r14 + r15;
assign R_temp_6 = r16 + r17 + r18;
assign R_temp_7 = r19 + r20 + r21;
assign R_temp_8 = r22 + r23 + r24;
assign R_temp_9 = r25 + r26 + r27;
assign R_temp_10 = r28 + r29 + r30;
assign R_temp_11 = r31 + r32 + r33;
assign R_temp_12 = r34 + r35 + r36;
assign R_temp_13 = r37 + r38 + r39;
assign R_temp_14 = r40 + r41 + r42;
assign R_temp_15 = r43 + r44 + r45;
assign R_temp_16 = r46 + r47 + r48;

wire [14:1] R_temp_17,R_temp_18,R_temp_19,R_temp_20,R_temp_21;

assign R_temp_17 = R_temp_1 + R_temp_2 + R_temp_3;
assign R_temp_18 = R_temp_4 + R_temp_5 + R_temp_6;
assign R_temp_19 = R_temp_7 + R_temp_8 + R_temp_9;
assign R_temp_20 = R_temp_10 + R_temp_11 + R_temp_12;
assign R_temp_21 = R_temp_13 + R_temp_14 + R_temp_15;

wire [15:1] R_temp_22,R_temp_23;

assign R_temp_22 = R_temp_17 + R_temp_18 + R_temp_19;
assign R_temp_23 = R_temp_20 + R_temp_21 + R_temp_16;

wire [13:1] R_temp_24,R_temp_25;

assign R_temp_24 = R_temp_22 [6:1] + 64 * R_temp_22 [11:7] + R_temp_23 [6:1] + 64* R_temp_23 [11:7]; 

assign R_temp_25 = 64 * r49 [11:7] + 37* R_temp_23 [15:12] + X[6:1] + r49 [6:1] +  37 * R_temp_22 [15:12]; 

wire [12:1] R_temp_26;

assign R_temp_26 = R_temp_24 [6:1] + 64 * R_temp_24 [11:7] + 37 * R_temp_24 [13:12] + R_temp_25 [6:1] + 64 * R_temp_25 [11:7] + 37 * R_temp_25 [13:12];

/*
wire [12:1] R_temp_24,R_temp_25,R_temp_26;

assign R_temp_24 = R_temp_22 [6:1] + 64 * R_temp_22 [11:7] + R_temp_23 [6:1];
            
assign R_temp_25 = 64* R_temp_23 [11:7] + r49 [6:1] +  37 * R_temp_22 [15:12]; 

assign R_temp_26 = 64 * r49 [11:7] + 37* R_temp_23 [15:12] + X[6:1]; 

wire [12:1] R_temp_27,R_temp_28;

assign R_temp_27 = R_temp_24 [6:1] + 64 * R_temp_24 [11:7] + 37 * R_temp_24 [12] + 64 * R_temp_26 [11:7];

assign R_temp_28 = R_temp_25 [6:1] + 64 * R_temp_25 [11:7] + 37 * R_temp_25 [12] + R_temp_26 [6:1] + 37 * R_temp_26 [12];

wire [12:1] R_temp_29;

assign R_temp_29 = R_temp_27 [6:1] + 64 * R_temp_27 [11:7] + 37 * R_temp_27 [12] + R_temp_28 [6:1] + 64 * R_temp_28 [11:7] + 37 * R_temp_28 [12];
*/

reg [11:1]  R_temp;

always @(R_temp_26)
begin
  if (R_temp_26 >= 11'b11111011011  )
    R_temp <= R_temp_26 - 11'b11111011011;
  else
    R_temp <= R_temp_26;
end

assign R = R_temp;

endmodule