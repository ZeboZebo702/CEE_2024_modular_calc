// Benchmark "X_15" written by ABC on Wed Jun 07 16:49:06 2023

module X_57 ( 
    x0, x1, x2, x3, x4, x5,
    z0, z1, z2, z3, z4, z5, z6  );
  input  x0, x1, x2, x3, x4, x5;
  output z0, z1, z2, z3, z4, z5, z6;
  assign z0 = 1'b0;
  assign z1 = x0;
  assign z2 = x1;
  assign z3 = x2;
  assign z4 = x3;
  assign z5 = x4;
  assign z6 = x5;
endmodule


