module mult_mod_461_bits(A,B,R
    );

    input [9:1] A;
    input [9:1] B;
    output [9:1] R;
wire [6:1] r1;
wire [9:1] r2;
wire [9:1] r3;
wire [9:1] r4;
wire [9:1] r5;
wire [9:1] r6;
wire [9:1] r7;
wire [9:1] r8;
wire [9:1] r9;

reg [9:1] temp_R;

mult_3x3  label1 (.x0(A[3]),.x1(A[2]),.x2(A[1]),
          .x3(B[3]),.x4(B[2]),.x5(B[1]),
          .z0(r1[6]),.z1(r1[5]),.z2(r1[4]),.z3(r1[3]),.z4(r1[2]),.z5(r1[1]));

mult_3x3_8  label2 (.x0(A[3]),.x1(A[2]),.x2(A[1]),
          .x3(B[6]),.x4(B[5]),.x5(B[4]),
          .z0(r2[9]),.z1(r2[8]),.z2(r2[7]),.z3(r2[6]),.z4(r2[5]),.z5(r2[4]),.z6(r2[3]),.z7(r2[2]),.z8(r2[1]));

mult_3x3_64  label3 (.x0(A[3]),.x1(A[2]),.x2(A[1]),
          .x3(B[9]),.x4(B[8]),.x5(B[7]),
	  .z0(r3[9]),.z1(r3[8]),.z2(r3[7]),.z3(r3[6]),.z4(r3[5]),.z5(r3[4]),.z6(r3[3]),.z7(r3[2]),.z8(r3[1]));


mult_3x3_8  label4 (.x0(A[6]),.x1(A[5]),.x2(A[4]),
          .x3(B[3]),.x4(B[2]),.x5(B[1]),
          .z0(r4[9]),.z1(r4[8]),.z2(r4[7]),.z3(r4[6]),.z4(r4[5]),.z5(r4[4]),.z6(r4[3]),.z7(r4[2]),.z8(r4[1]));

mult_3x3_64  label5 (.x0(A[6]),.x1(A[5]),.x2(A[4]),
          .x3(B[6]),.x4(B[5]),.x5(B[4]),
	  .z0(r5[9]),.z1(r5[8]),.z2(r5[7]),.z3(r5[6]),.z4(r5[5]),.z5(r5[4]),.z6(r5[3]),.z7(r5[2]),.z8(r5[1]));

mult_3x3_51  label6 (.x0(A[6]),.x1(A[5]),.x2(A[4]),
          .x3(B[9]),.x4(B[8]),.x5(B[7]),
	  .z0(r6[9]),.z1(r6[8]),.z2(r6[7]),.z3(r6[6]),.z4(r6[5]),.z5(r6[4]),.z6(r6[3]),.z7(r6[2]),.z8(r6[1]));


mult_3x3_64 label7 (.x0(A[9]),.x1(A[8]),.x2(A[7]),
          .x3(B[3]),.x4(B[2]),.x5(B[1]),
	  .z0(r7[9]),.z1(r7[8]),.z2(r7[7]),.z3(r7[6]),.z4(r7[5]),.z5(r7[4]),.z6(r7[3]),.z7(r7[2]),.z8(r7[1]));

mult_3x3_51  label8 (.x0(A[9]),.x1(A[8]),.x2(A[7]),
          .x3(B[6]),.x4(B[5]),.x5(B[4]),
	  .z0(r8[9]),.z1(r8[8]),.z2(r8[7]),.z3(r8[6]),.z4(r8[5]),.z5(r8[4]),.z6(r8[3]),.z7(r8[2]),.z8(r8[1]));

mult_3x3_408  label9 (.x0(A[9]),.x1(A[8]),.x2(A[7]),
          .x3(B[9]),.x4(B[8]),.x5(B[7]),
	  .z0(r9[9]),.z1(r9[8]),.z2(r9[7]),.z3(r9[6]),.z4(r9[5]),.z5(r9[4]),.z6(r9[3]),.z7(r9[2]),.z8(r9[1]));
/*

wire [11:1] temp_R_1,temp_R_2;

assign temp_R_1 = r2 + r3 + r4 + r5;

assign temp_R_2 = r6 + r7 + r8 + r9;


wire [9:1] r18,r19;


X_5_64  label18 (.x0(temp_R_1[11]),.x1(temp_R_1[10]),.x2(temp_R_1[9]),.x3(temp_R_1[8]),.x4(temp_R_1[7]),
	  .z0(r18[9]),.z1(r18[8]),.z2(r18[7]),.z3(r18[6]),.z4(r18[5]),.z5(r18[4]),.z6(r18[3]),.z7(r18[2]),.z8(r18[1]));

X_5_64  label19 (.x0(temp_R_2[11]),.x1(temp_R_2[10]),.x2(temp_R_2[9]),.x3(temp_R_2[8]),.x4(temp_R_2[7]),
	  .z0(r19[9]),.z1(r19[8]),.z2(r19[7]),.z3(r19[6]),.z4(r19[5]),.z5(r19[4]),.z6(r19[3]),.z7(r19[2]),.z8(r19[1]));


wire [10:1] temp_R_15;

assign temp_R_15 = temp_R_1[6:1] + r18 + r19 + r1 + temp_R_2[6:1];   
*/


wire [12:1] temp_R_1;

assign temp_R_1 = r1 + r2 + r3 + r4 + r5 + r6 + r7 + r8 + r9;


wire [9:1] r18;

X_6_64  label18 (.x0(temp_R_1[12]),.x1(temp_R_1[11]),.x2(temp_R_1[10]),.x3(temp_R_1[9]),.x4(temp_R_1[8]),.x5(temp_R_1[7]),
	  .z0(r18[9]),.z1(r18[8]),.z2(r18[7]),.z3(r18[6]),.z4(r18[5]),.z5(r18[4]),.z6(r18[3]),.z7(r18[2]),.z8(r18[1]));


wire [10:1] temp_R_15;

assign temp_R_15 = temp_R_1 [6:1] + r18;   




/*
assign temp_R_1 = r1 + r2 + r3 + r4 + r5 + r6 + r7 + r8 + r9;

mult_3_8  label10 (.x0(temp_R_1[6]),.x1(temp_R_1[5]),.x2(temp_R_1[4]),
	  .z0(r10[6]),.z1(r10[5]),.z2(r10[4]),.z3(r10[3]),.z4(r10[2]),.z5(r10[1]));

mult_3_64  label11 (.x0(temp_R_1[9]),.x1(temp_R_1[8]),.x2(temp_R_1[7]),
	  .z0(r11[9]),.z1(r11[8]),.z2(r11[7]),.z3(r11[6]),.z4(r11[5]),.z5(r11[4]),.z6(r11[3]),.z7(r11[2]),.z8(r11[1]));

mult_3_9  label12 (.x0(temp_R_1[12]),.x1(temp_R_1[11]),.x2(temp_R_1[10]),
	  .z0(r12[6]),.z1(r12[5]),.z2(r12[4]),.z3(r12[3]),.z4(r12[2]),.z5(r12[1]));


assign temp_R_2 = temp_R_1[3:1] + r10 + r11 + r12;
*/

always @(temp_R_15)
begin
  if (temp_R_15 >= 9'b111001101)
    temp_R <= temp_R_15 - 9'b111001101;
  else
    temp_R <= temp_R_15;
end

assign R = temp_R;

endmodule