module x_200_mod_997_reg(
    input [200:1] X,
    output [10:1] R
    );


assign R = X % 997;

endmodule
