// Benchmark "mult_3_9" written by ABC on Sun Dec 11 02:20:07 2022

module mult_3_9 ( 
    x0, x1, x2,
    z0, z1, z2, z3, z4, z5  );
  input  x0, x1, x2;
  output z0, z1, z2, z3, z4, z5;
  assign z0 = x0;
  assign z1 = x1;
  assign z2 = x2;
  assign z3 = x0;
  assign z4 = x1;
  assign z5 = x2;
endmodule


