module mult_const_128_bit_mod(
     a,
     r
    );

input [8:1] a;
output [258:1] r;

assign r = (a * 258'd428092581552246531046308046973043184312835253714261251748800951846523264768000) % 258'd429937808196868283335300754072064922176252647049236515764959576638965175392000;

endmodule