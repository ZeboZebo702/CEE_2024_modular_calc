// Benchmark "128_128_mod" written by ABC on Thu Dec 01 02:19:59 2022

module const_128_128_mod ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z000, z001, z002, z003, z004, z005, z006, z007, z008, z009, z010, z011,
    z012, z013, z014, z015, z016, z017, z018, z019, z020, z021, z022, z023,
    z024, z025, z026, z027, z028, z029, z030, z031, z032, z033, z034, z035,
    z036, z037, z038, z039, z040, z041, z042, z043, z044, z045, z046, z047,
    z048, z049, z050, z051, z052, z053, z054, z055, z056, z057, z058, z059,
    z060, z061, z062, z063, z064, z065, z066, z067, z068, z069, z070, z071,
    z072, z073, z074, z075, z076, z077, z078, z079, z080, z081, z082, z083,
    z084, z085, z086, z087, z088, z089, z090, z091, z092, z093, z094, z095,
    z096, z097, z098, z099, z100, z101, z102, z103, z104, z105, z106, z107,
    z108, z109, z110, z111, z112, z113, z114, z115, z116, z117, z118, z119,
    z120, z121, z122, z123, z124, z125, z126, z127, z128, z129, z130, z131,
    z132, z133, z134, z135, z136, z137, z138, z139, z140, z141, z142, z143,
    z144, z145, z146, z147, z148, z149, z150, z151, z152, z153, z154, z155,
    z156, z157, z158, z159, z160, z161, z162, z163, z164, z165, z166, z167,
    z168, z169, z170, z171, z172, z173, z174, z175, z176, z177, z178, z179,
    z180, z181, z182, z183, z184, z185, z186, z187, z188, z189, z190, z191,
    z192, z193, z194, z195, z196, z197, z198, z199, z200, z201, z202, z203,
    z204, z205, z206, z207, z208, z209, z210, z211, z212, z213, z214, z215,
    z216, z217, z218, z219, z220, z221, z222, z223, z224, z225, z226, z227,
    z228, z229, z230, z231, z232, z233, z234, z235, z236, z237, z238, z239,
    z240, z241, z242, z243, z244, z245, z246, z247, z248, z249, z250, z251,
    z252, z253, z254, z255, z256, z257  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z000, z001, z002, z003, z004, z005, z006, z007, z008, z009, z010,
    z011, z012, z013, z014, z015, z016, z017, z018, z019, z020, z021, z022,
    z023, z024, z025, z026, z027, z028, z029, z030, z031, z032, z033, z034,
    z035, z036, z037, z038, z039, z040, z041, z042, z043, z044, z045, z046,
    z047, z048, z049, z050, z051, z052, z053, z054, z055, z056, z057, z058,
    z059, z060, z061, z062, z063, z064, z065, z066, z067, z068, z069, z070,
    z071, z072, z073, z074, z075, z076, z077, z078, z079, z080, z081, z082,
    z083, z084, z085, z086, z087, z088, z089, z090, z091, z092, z093, z094,
    z095, z096, z097, z098, z099, z100, z101, z102, z103, z104, z105, z106,
    z107, z108, z109, z110, z111, z112, z113, z114, z115, z116, z117, z118,
    z119, z120, z121, z122, z123, z124, z125, z126, z127, z128, z129, z130,
    z131, z132, z133, z134, z135, z136, z137, z138, z139, z140, z141, z142,
    z143, z144, z145, z146, z147, z148, z149, z150, z151, z152, z153, z154,
    z155, z156, z157, z158, z159, z160, z161, z162, z163, z164, z165, z166,
    z167, z168, z169, z170, z171, z172, z173, z174, z175, z176, z177, z178,
    z179, z180, z181, z182, z183, z184, z185, z186, z187, z188, z189, z190,
    z191, z192, z193, z194, z195, z196, z197, z198, z199, z200, z201, z202,
    z203, z204, z205, z206, z207, z208, z209, z210, z211, z212, z213, z214,
    z215, z216, z217, z218, z219, z220, z221, z222, z223, z224, z225, z226,
    z227, z228, z229, z230, z231, z232, z233, z234, z235, z236, z237, z238,
    z239, z240, z241, z242, z243, z244, z245, z246, z247, z248, z249, z250,
    z251, z252, z253, z254, z255, z256, z257;
  wire n268, n269, n270, n271, n273, n274, n275, n276, n277, n278, n279,
    n281, n282, n283, n284, n285, n286, n287, n288, n290, n291, n292, n293,
    n294, n295, n296, n298, n299, n300, n301, n302, n303, n304, n305, n306,
    n307, n308, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
    n320, n321, n322, n323, n325, n326, n327, n328, n329, n330, n332, n333,
    n334, n335, n336, n337, n338, n339, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n352, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n390, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n410,
    n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
    n423, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n441, n442, n443, n444, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467, n468, n469, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n484, n485, n486,
    n487, n488, n489, n490, n491, n492, n493, n494, n496, n497, n498, n499,
    n500, n501, n502, n503, n504, n505, n506, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n520, n521, n522, n523, n524, n525,
    n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
    n550, n551, n552, n554, n555, n556, n557, n558, n559, n560, n561, n562,
    n563, n564, n566, n567, n568, n569, n570, n571, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n583, n584, n585, n586, n587, n588, n589,
    n590, n591, n592, n594, n595, n596, n597, n598, n600, n601, n602, n603,
    n605, n606, n607, n608, n610, n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
    n631, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
    n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
    n657, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n675, n676, n677, n678, n679, n680, n681, n682,
    n683, n685, n686, n687, n688, n689, n690, n691, n692, n693, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n715, n716, n717, n718, n719, n720, n721,
    n722, n723, n724, n725, n726, n727, n729, n730, n731, n732, n733, n734,
    n735, n736, n737, n738, n739, n740, n741, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754, n755, n756, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
    n799, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
    n812, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
    n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
    n838, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
    n851, n852, n853, n854, n855, n856, n858, n859, n860, n861, n862, n863,
    n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
    n876, n877, n878, n879, n881, n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n895, n896, n897, n898, n899, n900, n901,
    n902, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n915,
    n916, n917, n918, n919, n920, n921, n922, n923, n924, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n935, n936, n937, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n955, n956, n957, n958, n959, n960, n961, n963, n964, n965, n966, n967,
    n968, n969, n970, n971, n973, n974, n975, n976, n977, n978, n979, n980,
    n981, n982, n983, n984, n985, n987, n988, n989, n990, n991, n992, n993,
    n994, n995, n996, n997, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1026, n1027,
    n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
    n1038, n1039, n1040, n1041, n1042, n1044, n1045, n1046, n1047, n1048,
    n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1091,
    n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1115, n1116, n1117, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1132, n1133, n1134,
    n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
    n1145, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1183, n1184, n1185, n1186, n1187, n1188,
    n1189, n1190, n1191, n1192, n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1211,
    n1212, n1213, n1214, n1215, n1217, n1218, n1219, n1220, n1222, n1223,
    n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
    n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1332, n1333, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1373, n1374,
    n1375, n1376, n1377, n1378, n1379, n1381, n1382, n1383, n1384, n1385,
    n1386, n1387, n1388, n1389, n1390, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1400, n1401, n1402, n1403, n1404, n1406, n1407, n1408,
    n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1419, n1420,
    n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1430, n1431,
    n1432, n1433, n1434, n1435, n1436, n1437, n1439, n1440, n1441, n1442,
    n1443, n1444, n1445, n1446, n1447, n1448, n1450, n1451, n1452, n1453,
    n1454, n1455, n1456, n1457, n1458, n1460, n1461, n1462, n1463, n1464,
    n1465, n1466, n1467, n1468, n1469, n1470, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1484, n1485, n1486,
    n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
    n1508, n1509, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
    n1519, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1546, n1547, n1548, n1549, n1550, n1551,
    n1552, n1553, n1554, n1555, n1557, n1558, n1559, n1560, n1561, n1562,
    n1563, n1564, n1565, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1576, n1577, n1578, n1579, n1580, n1581, n1583, n1584, n1585,
    n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
    n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1618,
    n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
    n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1648, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
    n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
    n1672, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
    n1683, n1684, n1685, n1686, n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1703, n1704,
    n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
    n1715, n1716, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
    n1737, n1738, n1739, n1740, n1742, n1743, n1744, n1745, n1746, n1747,
    n1748, n1749, n1750, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
    n1759, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
    n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
    n1781, n1782, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
    n1792, n1793, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
    n1803, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
    n1814, n1815, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
    n1825, n1826, n1827, n1828, n1829, n1831, n1832, n1833, n1834, n1835,
    n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1846,
    n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
    n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1890, n1891,
    n1892, n1893, n1894, n1896, n1897, n1898, n1899, n1901, n1902, n1903,
    n1904, n1905, n1906, n1908, n1909, n1910, n1912, n1913, n1914, n1915,
    n1916, n1917, n1918, n1919, n1921, n1922, n1923, n1924, n1925, n1926,
    n1927, n1928, n1929, n1931, n1932, n1933, n1934, n1936, n1937, n1938,
    n1939, n1940, n1942, n1943, n1944, n1945, n1946, n1948, n1949, n1950,
    n1952, n1953, n1955, n1956, n1957, n1958, n1960, n1961, n1962, n1963,
    n1964, n1965, n1966, n1967, n1968, n1969, n1971, n1972, n1973, n1974,
    n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1983, n1984, n1985,
    n1986, n1987, n1988, n1989, n1990, n1992, n1993, n1994, n1995, n1996,
    n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
    n2007, n2008, n2009, n2010, n2012, n2013, n2014, n2015, n2016, n2017,
    n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2026, n2027, n2028,
    n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2038, n2039,
    n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
    n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2082,
    n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
    n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
    n2104, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
    n2115, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
    n2126, n2127, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
    n2137, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
    n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
    n2159, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
    n2171, n2172, n2173, n2174, n2176, n2177, n2178, n2179, n2180, n2181,
    n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2190, n2191, n2192,
    n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2202, n2203,
    n2204, n2205, n2206, n2207, n2208, n2209, n2211, n2212, n2213, n2214,
    n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2225, n2226,
    n2227, n2228, n2229, n2230, n2231, n2232, n2234, n2235, n2236, n2237,
    n2238, n2239, n2240, n2242, n2243, n2244, n2245, n2246, n2248, n2249,
    n2250, n2251, n2252, n2253, n2254, n2255, n2257, n2258, n2259, n2260,
    n2261, n2262, n2263, n2264, n2265, n2266, n2268, n2269, n2270, n2271,
    n2272, n2273, n2274, n2275, n2276, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
    n2294, n2295, n2296, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
    n2305, n2306, n2307, n2308, n2309, n2310, n2312, n2313, n2314, n2315,
    n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2324, n2325, n2326,
    n2327, n2328, n2329, n2330, n2331, n2332, n2334, n2335, n2336, n2337,
    n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2347, n2348,
    n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2359,
    n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
    n2370, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
    n2381, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2397, n2398, n2399, n2400, n2401, n2402,
    n2403, n2404, n2406, n2407, n2408, n2409, n2410, n2411, n2413, n2414,
    n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2423, n2424, n2425,
    n2426, n2427, n2428, n2429, n2430, n2432, n2433, n2434, n2435, n2436,
    n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2445, n2446, n2447,
    n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
    n2459, n2460, n2462, n2463, n2464, n2465, n2467, n2468, n2469, n2470,
    n2471, n2472, n2473, n2474, n2475, n2477, n2478, n2479, n2480, n2481,
    n2482, n2483, n2484, n2485, n2486, n2488, n2489, n2490, n2491, n2492,
    n2493, n2494, n2495, n2496, n2497, n2498, n2500, n2501, n2502, n2503,
    n2504, n2505, n2506, n2507, n2509, n2510, n2511, n2512, n2513, n2514,
    n2515, n2516, n2517, n2518, n2519, n2521, n2522, n2523, n2524, n2525,
    n2526, n2527, n2528, n2529, n2530, n2531, n2533, n2534, n2535, n2536,
    n2537, n2538, n2539, n2541, n2542, n2543, n2544, n2546, n2547, n2548,
    n2550, n2551, n2552, n2553, n2554, n2555, n2557, n2558, n2559, n2560,
    n2562, n2563, n2564, n2565, n2566, n2568, n2569, n2570, n2571, n2572,
    n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2584,
    n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2595,
    n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
    n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
    n2617, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
    n2628, n2629, n2630, n2631, n2633, n2634, n2635, n2636, n2637, n2638,
    n2639, n2640, n2641, n2642, n2643, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2670, n2671,
    n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2681, n2682,
    n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2692, n2693,
    n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
    n2704, n2705, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
    n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
    n2726, n2727, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
    n2737, n2738, n2739, n2740, n2742, n2743, n2744, n2745, n2746, n2747,
    n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2756, n2757, n2758,
    n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
    n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2778, n2779, n2780,
    n2781, n2782, n2783, n2785, n2786, n2787, n2788, n2790, n2791, n2792,
    n2793, n2794, n2796, n2798, n2799, n2803, n2804, n2806, n2807, n2808,
    n2809, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2819, n2820,
    n2821, n2822, n2823, n2824, n2825, n2826, n2828, n2829, n2830, n2831,
    n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2840, n2841, n2842,
    n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
    n2864, n2865, n2866, n2867, n2869, n2870, n2871, n2872, n2873, n2874,
    n2875, n2876, n2877, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
    n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2896, n2897,
    n2898, n2899, n2900, n2902, n2903, n2904, n2905, n2907, n2908, n2909,
    n2910, n2912, n2913, n2914, n2915, n2917, n2920, n2921, n2922, n2923,
    n2924, n2926, n2928, n2929, n2930, n2931, n2932, n2933;
  assign z250 = 1'b0;
  assign z000 = ~x0 & ((n268 & n269) | ~n270 | ~n271);
  assign n268 = ~x3 & ~x1 & ~x2;
  assign n269 = x7 & ~x6 & ~x4 & ~x5;
  assign n270 = x1 ? x2 : (~x2 & ~x3 & (x4 | x5 | ~x6));
  assign n271 = x3 | (x1 ? (~x2 | (x4 & x5)) : (x2 | (~x4 & ~x5)));
  assign z001 = n275 | ~n276 | (n273 & ~n274);
  assign n273 = ~x1 & ~x3;
  assign n274 = (x0 | x6 | ((x2 | x4 | x5 | ~x7) & (~x2 | ~x4 | ~x5 | x7))) & (~x0 | ~x2 | ~x4 | x5 | ~x6 | x7);
  assign n275 = ~x0 & ~x3 & ((~x1 & (x2 ? (x4 & ~x5) : (~x4 & x5))) | (x1 & x2 & x4 & x5));
  assign n276 = ~n277 & ((x1 & (~x2 | ~x3)) | (x2 & (x3 ? (x0 | ~x1) : x4)) | (~x3 & ~x4 & ~x0 & ~x2));
  assign n277 = ~x5 & n273 & (x4 ? (~x6 & n279) : (x6 & n278));
  assign n278 = ~x0 & ~x2;
  assign n279 = x0 & x2;
  assign z002 = ~n286 | n281 | n285;
  assign n281 = ~x3 & ((n283 & n284) | (~x1 & ~n282));
  assign n282 = (~x4 | ((~x0 | x5 | ~x6 | (x2 ^ x7)) & (x0 | ~x2 | ~x5 | x6 | ~x7))) & (x5 | x6 | ~x7 | x0 | x2 | x4);
  assign n283 = ~x2 & ~x0 & x1;
  assign n284 = ~x7 & ~x6 & x4 & x5;
  assign n285 = ~x3 & ((x5 & ((~x0 & (x1 ? (x2 & x4) : (~x2 & ~x4))) | (x0 & ~x1 & x2 & x4))) | (x4 & ~x5 & ~x0 & ~x2));
  assign n286 = (~x2 | ~x3 | (x0 & x1)) & (x3 | n287) & (x2 | (~x0 & ~x1) | ~n288);
  assign n287 = (x0 | x1 | ((x2 | (x4 ? (~x5 | x6) : (x5 | ~x6))) & (~x5 | ~x6 | ~x2 | ~x4))) & (~x0 | x2 | ~x4 | x5 | x6);
  assign n288 = ~x3 & ~x4;
  assign z003 = n291 | (x0 ? (~n290 | (~x2 & ~n295)) : (~n296 | (x2 & ~n295)));
  assign n290 = (x1 | ((~x2 | (x3 ? (x4 & (x5 | x6)) : (~x4 | ~x5))) & (~x5 | x6 | x3 | ~x4))) & (~x4 | x5 | ~x6 | ~x1 | x2 | x3);
  assign n291 = x4 & ((~x1 & ~n293) | (n292 & n283 & n294));
  assign n292 = ~x6 & x7;
  assign n293 = x0 ? (x5 | ~x6 | ((x3 | ~x7) & (x2 | ~x3 | x7))) : (~x2 | ~x5 | x6 | (~x3 ^ x7));
  assign n294 = ~x3 & x5;
  assign n295 = x3 ? (x4 & (x5 | x6)) : (~x4 | ~x5 | (~x1 & ~x6));
  assign n296 = (~x4 | ~x6 | ((x2 | x3 | ~x5) & (~x3 | x5))) & (x2 | ~x3 | (x4 & x5 & (x1 | x6)));
  assign z004 = ~n298 | ~n302 | n306 | (~n307 & ~n308);
  assign n298 = ~n299 & n301 & (x5 | ~n279 | n300);
  assign n299 = ~x0 & x2 & (x1 ? (x4 & x5) : (~x4 & ~x5));
  assign n300 = (~x1 | x3 | x4 | x6) & (~x4 | ~x6 | x1 | ~x3);
  assign n301 = x4 ? (~x5 | (x1 & x2) | (~x0 & ~x6)) : (x5 | ((~x1 | (x0 & (x2 | x6))) & (~x0 | x1 | x6)));
  assign n302 = (x2 | n303) & (n304 | ~n305);
  assign n303 = (x0 | ~x3 | x6 | (x1 ? (~x4 | ~x5) : (x4 | x5))) & (x4 | x5 | ~x6 | ~x0 | x1 | x3);
  assign n304 = (x4 | x6 | ~x7 | x0 | x2 | x3) & (~x0 | ~x6 | ((x2 | x3 | ~x4 | ~x7) & (~x2 | ~x3 | x4 | x7)));
  assign n305 = ~x1 & ~x5;
  assign n306 = ~x2 & ((~x0 & ~x1 & ~x4 & (x5 ^ x6)) | (x0 & x1 & x4 & ~x5 & x6));
  assign n307 = ~x4 ^ ~x7;
  assign n308 = (x1 | ((~x0 | x5 | ~x6 | (~x2 ^ x3)) & (~x5 | x6 | x0 | ~x2))) & (x3 | ~x5 | x6 | x0 | ~x1 | x2);
  assign z005 = ~n311 | ~n320 | (n310 & ~n319) | (x5 & ~n318);
  assign n310 = ~x0 & ~x6;
  assign n311 = ~n314 & (n315 | n316) & (~n312 | ~n313 | ~n317);
  assign n312 = ~x5 & ~x6;
  assign n313 = ~x3 & x4;
  assign n314 = ~x1 & ((~x0 & ((~x3 & x5 & x6) | (~x5 & ~x6 & ~x2 & x3))) | (x5 & ~x6 & x0 & ~x3));
  assign n315 = x1 ? (x3 | x4) : (~x3 | ~x4);
  assign n316 = x0 ? ((~x5 | x6) & (~x2 | x5 | ~x6)) : (~x5 | ~x6);
  assign n317 = ~x2 & ~x0 & ~x1;
  assign n318 = x0 ? (x6 | ((x3 | ~x4 | ~x1 | x2) & (x1 | ~x3 | x4))) : (~x6 | (x1 ? (x3 | ~x4) : (~x3 | x4)));
  assign n319 = ((x5 ^ x7) | (x1 ? (x2 | x3) : ~x2)) & (x2 | x4 | x5 | (x1 ? x7 : (x3 | ~x7)));
  assign n320 = ~n322 & (~x6 | ~n321 | n323);
  assign n321 = x0 & ~x1;
  assign n322 = x1 & ((x5 & ((~x0 & (x3 | (x2 & ~x6))) | (~x2 & x3 & ~x6))) | (~x5 & x6 & x0 & ~x2));
  assign n323 = (x7 & (x5 | (~x2 & ~x3 & ~x4))) | (~x5 & ~x7) | (x2 & x3 & x4);
  assign z006 = ~n330 | n325 | ~n326;
  assign n325 = ~x1 & (x0 ? ((x6 & x7 & x2 & x3) | (~x6 & ~x7 & ~x2 & ~x3)) : (x2 ? ((~x6 & x7) | (x3 & x6 & ~x7)) : (x6 & (~x3 | x7))));
  assign n326 = x4 ? n328 : ((x2 | n327) & (~x0 | ~x2 | n329));
  assign n327 = x0 ? (x1 | x3 | ~x7 | (x5 ^ x6)) : (~x1 | ~x3 | x7 | (~x5 ^ x6));
  assign n328 = (~x0 | x1 | ~x6 | (x2 ? (~x3 | x7) : (x3 | ~x7))) & (~x3 | x6 | x7 | x0 | ~x1 | x2);
  assign n329 = (~x1 | x3 | ~x6) & (x1 | ~x3 | x6 | x7);
  assign n330 = (x0 & (x1 ? ~x6 : (x6 & ~x7))) | (x2 & (x1 ? x6 : x3)) | (x1 & ((~x0 & x3 & x6) | (~x2 & ~x6 & ~x7))) | (~x0 & (x6 ? x7 : ~x1)) | (~x1 & ((~x6 & x7) | (~x2 & ~x3)));
  assign z007 = n336 | n337 | ~n338 | (~x4 & (~n332 | ~n333));
  assign n332 = (x2 | ((x1 | x3 | (x0 ? (x5 ^ x7) : (~x5 | x7))) & (x0 | ~x1 | ~x3 | ~x5 | x7))) & (~x3 | x5 | ~x7 | ~x0 | x1 | ~x2);
  assign n333 = (~n292 | ~n283 | ~n335) & (x1 | n334);
  assign n334 = (~x0 | ~x5 | x6 | (x2 ? (~x3 | ~x7) : (x3 | x7))) & (x5 | ~x6 | x7 | x0 | x2 | x3);
  assign n335 = x3 & ~x5;
  assign n336 = ~x3 & ((x0 & ((~x1 & ~x2 & x4 & x7) | (x1 & x2 & ~x4 & ~x7))) | (~x0 & ~x1 & ~x2 & x4 & ~x7));
  assign n337 = (x3 ? (x4 & ~x7) : x7) & (x0 ? (~x1 & x2) : (x1 & ~x2));
  assign n338 = x1 ? (x0 ? (x2 ? (x3 | ~n339) : x7) : (~x2 | x7)) : ((x0 | (x2 ? ~x7 : (~x3 | x7))) & (~x3 | ~x7 | ~x0 | x2));
  assign n339 = ~x7 & ~x6 & x4 & ~x5;
  assign z008 = n341 | n344 | ~n348 | (x3 ? ~n346 : ~n347);
  assign n341 = ~x1 & ((n342 & n339) | (~x4 & ~n343));
  assign n342 = x3 & ~x0 & x2;
  assign n343 = (x5 | x6 | ~x7 | x0 | x2 | x3) & (~x5 | ((x0 | x2 | x3 | ~x6 | x7) & (~x0 | ~x7 | (x2 ? (~x3 | ~x6) : (x3 | x6)))));
  assign n344 = n345 & ((x5 & ((x0 & (x3 ? (x4 & ~x6) : (~x4 & x6))) | (~x0 & ~x3 & ~x4 & ~x6))) | (~x0 & ~x3 & ~x4 & ~x5 & x6));
  assign n345 = ~x1 & ~x2;
  assign n346 = (x1 | (x0 ? (x2 ^ x4) : (~x2 | x4))) & (x0 | ~x1 | x2 | ~x4);
  assign n347 = x2 ? (x0 | (x1 & x4)) : (~x0 | (~x1 & ~x4));
  assign n348 = n350 & (~n349 | ((x2 | ~x3 | x4 | ~x5) & (~x2 | x3 | ~x4 | x5)));
  assign n349 = ~x0 & x1;
  assign n350 = x2 | ~x3 | (x0 ? (x1 | ~n351) : (~x1 | ~n352));
  assign n351 = x4 & ~x5;
  assign n352 = x7 & x6 & ~x4 & ~x5;
  assign z009 = n355 | ~n356 | ~n364 | n375 | (n354 & ~n376);
  assign n354 = ~x1 & x2;
  assign n355 = ~x4 & (x1 ? (x3 & (~x0 ^ ~x2)) : (x2 & ~x3));
  assign n356 = ~n360 & ~n363 & (~n359 | (~n357 & (~x0 | ~n358)));
  assign n357 = ~x2 & ~x3;
  assign n358 = x2 & x3;
  assign n359 = ~x1 & x4;
  assign n360 = ~x2 & x5 & ~n362 & (n288 | n361);
  assign n361 = x3 & x4;
  assign n362 = x0 ? (x1 | ~x6) : (~x1 | x6);
  assign n363 = n354 & n351 & (x0 ? (~x3 & ~x6) : (x3 & x6));
  assign n364 = ~n365 & (x2 | (~n366 & ~n371));
  assign n365 = ~x0 & ~x1 & ((~x4 & ~x5 & ~x2 & x3) | (x2 & x4 & (~x3 ^ x5)));
  assign n366 = x5 & ~n368 & ((n367 & n369) | (n273 & n370));
  assign n367 = x1 & x3;
  assign n368 = x0 ^ ~x6;
  assign n369 = x4 & ~x7;
  assign n370 = ~x4 & x7;
  assign n371 = ~x5 & n373 & ((n372 & n321) | (n349 & n374));
  assign n372 = ~x6 & ~x7;
  assign n373 = x3 & ~x4;
  assign n374 = x6 & x7;
  assign n375 = x1 & ((~x0 & x5 & (x2 ? (~x3 & x4) : (x3 & ~x4))) | (~x2 & ~x5 & (~x3 ^ x4)));
  assign n376 = x0 ? (~x6 | ((~x5 | ~x7 | ~x3 | x4) & (x5 | x7 | x3 | ~x4))) : (~x4 | x6 | (x3 ? (x5 | ~x7) : (~x5 | x7)));
  assign z010 = ~n380 | (x2 ? ~n378 : ~n379);
  assign n378 = (x6 | ((~x1 | ((~x4 | ~x5 | x0 | ~x3) & (x4 | x5 | ~x0 | x3))) & (x0 | x4 | ((x1 | x3 | ~x5) & (~x3 | x5))))) & (x0 | x1 | ~x4 | ~x6 | (~x3 ^ x5));
  assign n379 = x0 ? (x4 ? (x3 ? (~x5 | ~x6) : (x5 | x6)) : ((x1 | ~x6 | (~x3 ^ x5)) & (~x1 | ~x3 | ~x5 | x6))) : ((~x1 | x3 | x4 | ~x5 | ~x6) & (~x4 | x5 | x6 | x1 | ~x3));
  assign n380 = n381 & (x3 ? (n388 & (n382 | n387)) : n383);
  assign n381 = ((~x3 ^ x5) | ((~x0 | (x1 ? (x2 | x4) : (~x2 | ~x4))) & (x0 | ~x1 | ~x2 | ~x4))) & (x0 | (x2 ? ((~x4 | ~x5 | x1 | ~x3) & (x3 | x4 | x5)) : (x3 ? (x4 | ~x5) : (~x4 | x5)))) & (x1 | x4 | (x2 ? (x3 | x5) : (~x3 | ~x5)));
  assign n382 = x2 ^ ~x7;
  assign n383 = (~x5 | ((~n384 | n386) & (x0 | x6 | n385))) & (~x0 | x5 | ~x6 | n385);
  assign n384 = ~x1 & ~x4;
  assign n385 = (x1 | ~x4 | (~x2 ^ ~x7)) & (~x1 | ~x2 | x4 | x7);
  assign n386 = (x0 | ~x6 | (x2 ^ ~x7)) & (~x0 | x2 | x6 | ~x7);
  assign n387 = (~x0 | x1 | x4 | x5 | x6) & (x0 | ~x1 | ~x4 | ~x5 | ~x6);
  assign n388 = x0 ? (~x5 | (x1 ? (x2 | n389) : (~x2 | n390))) : (x5 | (x1 ? (x2 | n390) : (~x2 | n389)));
  assign n389 = x4 ? (x6 | ~x7) : (~x6 | x7);
  assign n390 = x4 ? (x6 | x7) : (~x6 | ~x7);
  assign z011 = n394 | n396 | ~n397 | (~n392 & ~n393) | ~n405;
  assign n392 = ~x3 ^ ~x7;
  assign n393 = (x4 | ((~x6 | (x1 ^ ~x2) | (~x0 ^ ~x5)) & (~x0 | x1 | ~x2 | x5 | x6))) & (~x1 | ~x4 | ((x0 | ((~x5 | ~x6) & (x2 | x5 | x6))) & (~x5 | x6 | ~x0 | x2)));
  assign n394 = ~n395 & x2 & x7;
  assign n395 = (~x0 | ((x1 | ~x4 | (x3 ? (~x5 | x6) : (x5 | ~x6))) & (x4 | x5 | ~x6 | ~x1 | x3))) & (x0 | x1 | x3 | x4 | ~x5 | ~x6);
  assign n396 = n345 & ((~x3 & ((x5 & x6 & x0 & ~x4) | ((~x4 ^ x5) & (x0 ^ x6)))) | (~x0 & x3 & ~x4 & x5 & ~x6));
  assign n397 = ~n398 & n401 & ((~x3 & (x4 | x6)) | (x4 & x6) | ~n400 | (x3 & ~x4 & ~x6));
  assign n398 = ~n399 & ((~x0 & ~x4 & ~x6 & (~x1 ^ ~x2)) | (x0 & x1 & ~x2 & x4 & x6));
  assign n399 = ~x3 ^ ~x5;
  assign n400 = ~x5 & x2 & ~x0 & x1;
  assign n401 = ~n403 & n404 & ((x6 & (x0 | ~x4)) | n402 | (~x0 & ~x6));
  assign n402 = (x1 | ~x2 | x3 | ~x5) & (~x1 | x2 | ~x3 | x5);
  assign n403 = (x4 ^ x6) & ((x0 & ~x1 & x3 & ~x5) | (~x0 & x1 & ~x3 & x5));
  assign n404 = x0 ? (~x5 | ((~x4 | ~x6 | x1 | ~x3) & (x4 | x6 | ~x1 | x3))) : (x1 | ~x4 | x5 | (~x3 ^ ~x6));
  assign n405 = (n406 | n408) & (n407 | (x0 ? (x2 | x4) : (~x2 | ~x4)));
  assign n406 = x3 ^ ~x7;
  assign n407 = (x5 | ((~x1 | x7 | (~x3 ^ ~x6)) & (x1 | ~x3 | x6 | ~x7))) & (x1 | ~x5 | x6 | (x3 ^ ~x7));
  assign n408 = (x1 | x2 | ((~x4 | (x0 ? (x5 | ~x6) : (~x5 | x6))) & (x0 | x4 | (x5 ^ x6)))) & (x4 | ~x5 | x6 | x0 | ~x1 | ~x2);
  assign z012 = ~n415 | (x1 ? ~n410 : (x0 ? ~n414 : ~n413));
  assign n410 = x4 ? n412 : n411;
  assign n411 = (~x6 | ((~x7 | (x0 ? (x2 ? (x3 | x5) : ~x3) : (x2 | x5))) & (x0 | ~x2 | ~x3 | ~x5 | x7))) & (x3 | x6 | (x0 ? (~x5 | x7) : (x2 ? (~x5 | ~x7) : (x5 | x7))));
  assign n412 = (x5 | ~x6 | x7 | x0 | x2 | x3) & (~x5 | (x0 ? (x2 | ((x6 | ~x7) & (x3 | ~x6 | x7))) : (~x2 | ((x6 | x7) & (~x3 | ~x6 | ~x7)))));
  assign n413 = (~x3 | ((x2 | ~x5 | x7 | (x4 ^ x6)) & (x6 | ~x7 | ~x2 | ~x4))) & (~x7 | ((~x2 | x4 | ~x6 | (x3 & x5)) & (~x4 | ~x5 | x6)));
  assign n414 = x4 ? (x2 ? (~x7 | (x3 ? (~x5 | x6) : (x5 | ~x6))) : (x6 | x7 | (x3 ^ ~x5))) : (x5 | ((x3 | ~x6 | x7) & (x2 | ((~x6 | x7) & (~x3 | x6 | ~x7)))));
  assign n415 = n417 & (n416 | n423) & (~x2 | n422);
  assign n416 = ~x5 ^ ~x6;
  assign n417 = (n420 | n421) & (x2 | n418) & (n416 | n419);
  assign n418 = x0 ? ((~x1 | x5 | (x3 ? (x4 | x6) : (~x4 | ~x6))) & (x1 | ~x3 | ~x4 | ~x5 | ~x6)) : ((~x5 | ((~x1 | ((~x4 | x6) & (x3 | x4 | ~x6))) & (x1 | x3 | x4 | x6))) & (x5 | ~x6 | x1 | ~x4));
  assign n419 = (~x0 | x3 | (x1 ? (~x2 | x4) : (x2 | ~x4))) & (x0 | x1 | ~x2 | ~x3 | x4);
  assign n420 = x4 ? (x5 | ~x6) : (~x5 | x6);
  assign n421 = x0 ? (x2 | (x1 ? (~x3 | x7) : ~x7)) : (~x2 | (x1 ? (~x3 | ~x7) : x7));
  assign n422 = (x1 | ((~x0 | ((x4 | ~x5 | x6) & (x5 | ~x6 | ~x3 | ~x4))) & (x0 | x3 | x4 | x5 | x6))) & (x0 | ~x1 | x5 | ((x4 | ~x6) & (~x3 | ~x4 | x6)));
  assign n423 = x1 ? ((x0 | ((x2 | ((~x4 | ~x7) & (~x3 | x4 | x7))) & (x3 | ((~x4 | ~x7) & (~x2 | x4 | x7))))) & (x3 | x4 | ~x7 | ~x0 | x2)) : (x0 ? (~x2 | (~x4 ^ x7)) : (x2 | ((x4 | ~x7) & (x3 | ~x4 | x7))));
  assign z013 = n427 | n430 | ~n436 | (~n425 & ~n426);
  assign n425 = ~x6 ^ ~x7;
  assign n426 = x0 ? ((~x1 | x3 | x4 | (~x2 ^ x5)) & (x2 | ~x3 | x5) & (x1 | (~x2 ^ ~x5))) : ((x1 | (x2 ? x5 : (x4 | ~x5))) & (~x2 | ((~x3 | ~x4 | x5) & (~x1 | x3 | ~x5))) & (x2 | ((~x1 | ((~x4 | ~x5) & (x3 | x4 | x5))) & (~x5 | (~x3 ^ x4)))));
  assign n427 = ~x3 & (x1 ? ~n429 : ~n428);
  assign n428 = x2 ? (x0 ? ((~x5 | ~x6 | x7) & (x6 | ~x7 | ~x4 | x5)) : ((x5 | ~x6 | x7) & (x6 | ~x7 | x4 | ~x5))) : ((~x5 | x6 | ~x7 | x0 | ~x4) & (x5 | ~x6 | x7 | ~x0 | x4));
  assign n429 = x2 ? ((x0 | ((~x5 | x6 | ~x7) & (~x6 | x7 | ~x4 | x5))) & (~x0 | ~x4 | x5 | x6 | x7)) : ((x4 | ((~x0 | (x5 ? (x6 | ~x7) : (~x6 | x7))) & (x6 | ~x7 | x0 | x5))) & (~x5 | ~x6 | x7 | x0 | ~x4));
  assign n430 = x3 & (~n433 | (~n431 & n432));
  assign n431 = (x1 | x6 | ~x7 | (x2 ^ x5)) & (~x1 | x2 | x5 | ~x6 | x7);
  assign n432 = x0 & x4;
  assign n433 = ((x1 ? n434 : n435) | (x0 ? (x2 | x4) : (~x2 | ~x4))) & (x0 | x2 | x4 | (x1 ? n435 : n434));
  assign n434 = x5 ? (x6 | ~x7) : (~x6 | x7);
  assign n435 = x5 ? (~x6 | x7) : (x6 | ~x7);
  assign n436 = ~n439 & n441 & (n437 | n438);
  assign n437 = x6 ^ ~x7;
  assign n438 = x0 ? ((~x5 | (x1 ? (x2 ? (x3 | x4) : (~x3 | ~x4)) : (x2 | x3))) & (~x3 | x5 | x1 | ~x2)) : ((x5 | (x1 ? (x2 ? (x3 | x4) : (~x3 | ~x4)) : (x2 | x3))) & (x1 | ~x2 | ~x5 | (~x3 ^ x4)));
  assign n439 = ~n440 & ((~x0 & x3 & (x1 ? (x2 & ~x4) : (~x2 & x4))) | (x0 & x1 & ~x2 & ~x3 & x4));
  assign n440 = ~x5 ^ ~x7;
  assign n441 = (~n321 | n442) & (x3 | n443 | ~n444);
  assign n442 = (x2 | ~x3 | ~x4 | ~x5 | x7) & (~x2 | x3 | x4 | x5 | ~x7);
  assign n443 = x4 ? (x5 | ~x7) : (~x5 | x7);
  assign n444 = ~x2 & ~x0 & x1;
  assign z014 = ~n446 | ~n457 | (~n437 & ~n468) | (~n425 & ~n469);
  assign n446 = ~n449 & ~n453 & (n447 | n448) & (n455 | n456);
  assign n447 = x3 ? (~x4 | x6) : (x4 | ~x6);
  assign n448 = (~x0 | x1 | x2 | ~x5) & (x0 | ~x1 | ~x2 | x5);
  assign n449 = ~x3 & n278 & ((n451 & n452) | (n450 & n359));
  assign n450 = ~x5 & x6;
  assign n451 = x5 & ~x6;
  assign n452 = x1 & ~x4;
  assign n453 = ~n454 & (x2 ? (~x4 & n321) : (x4 & n349));
  assign n454 = (~x3 | x5 | x6 | x7) & (~x6 | ~x7 | x3 | ~x5);
  assign n455 = (x0 | x1 | ~x2 | x3) & (~x0 | ~x1 | x2 | ~x3);
  assign n456 = (~x4 | ~x5 | x6 | x7) & (x4 | x5 | ~x6 | ~x7);
  assign n457 = n458 & n461 & n465 & ~n466 & (n455 | n467);
  assign n458 = ~x4 | ~x6 | (x3 ? (x5 | ~n459) : ~n460);
  assign n459 = x2 & x0 & ~x1;
  assign n460 = ~x2 & x0 & ~x1;
  assign n461 = (~n463 | ~n464) & (~n351 | ~n462 | ~n374);
  assign n462 = x3 & x2 & ~x0 & x1;
  assign n463 = ~x3 & ~x2 & x0 & ~x1;
  assign n464 = ~x7 & ~x6 & ~x4 & x5;
  assign n465 = ((x1 ^ x6) | ((~x3 | ~x4 | x0 | x2) & (x3 | x4 | ~x0 | ~x2))) & (~x3 | x4 | ~x6 | x1 | ~x2) & (x3 | ~x4 | x6 | ~x1 | x2);
  assign n466 = ~x0 & ~x4 & ((~x1 & ~x2 & ~x3 & x6) | (x1 & x2 & x3 & ~x6));
  assign n467 = x4 ? (~x5 | ~x6) : (x5 | x6);
  assign n468 = x2 ? ((~x4 | ~x5 | x1 | ~x3) & (x0 | (x1 ? (x3 | (~x4 & ~x5)) : (~x3 | ~x4)))) : ((~x0 | (x1 ? (x3 | x4) : (~x3 | x5))) & (x1 | ((~x3 | x4) & (~x4 | ~x5 | x0 | x3))) & (x4 | x5 | ~x1 | x3));
  assign n469 = x1 ? (~x3 | ((x0 | (x2 ? (~x4 | ~x5) : x4)) & (x2 | ((x4 | ~x5) & (~x0 | ~x4 | x5))))) : (x3 | ((~x0 | (x2 ? ~x4 : (x4 | x5))) & (~x2 | ((~x4 | x5) & (x0 | x4 | ~x5)))));
  assign z015 = ~n479 | (x0 ? (~n474 | ~n475) : ~n471);
  assign n471 = x5 ? n473 : n472;
  assign n472 = (x3 | x4 | ((x1 | (x2 ? (x6 ^ x7) : (~x6 | x7))) & (x6 | ~x7 | ~x1 | x2))) & (~x1 | ~x3 | ~x4 | (x2 ? (~x6 | ~x7) : (~x6 ^ x7)));
  assign n473 = x1 ? (x3 | ((x6 | x7 | ~x2 | x4) & (x2 | ~x4 | (x6 ^ x7)))) : ((x4 | x6 | ~x7 | x2 | ~x3) & (~x4 | ~x6 | x7 | ~x2 | x3));
  assign n474 = (x4 | ~x5 | x7 | x1 | ~x2 | ~x3) & (x2 | ((x5 | ~x7 | ~x3 | ~x4) & (x1 | ((x5 | ~x7 | x3 | x4) & (~x5 | x7 | ~x3 | ~x4)))));
  assign n475 = (n437 | n477) & (~x5 | ~n354 | n478) & (x5 | n476);
  assign n476 = (~x1 | ((x4 | ~x6 | ~x7 | x2 | ~x3) & (~x4 | x6 | x7 | ~x2 | x3))) & (x4 | x6 | x7 | x1 | x2 | ~x3);
  assign n477 = (x1 | x4 | (x2 ? (~x3 | x5) : (x3 | ~x5))) & (~x1 | x2 | ~x3 | ~x4 | ~x5);
  assign n478 = (~x3 | ~x4 | x6 | x7) & (x3 | x4 | ~x6 | ~x7);
  assign n479 = n482 & (x0 | n480) & (n440 | n481);
  assign n480 = (x2 | ((x7 | ((x3 | x4 | ~x5) & (~x1 | ~x4 | (x3 ^ x5)))) & (x4 | x5 | ~x7 | x1 | ~x3))) & (x1 | ~x2 | x3 | ~x7 | (~x4 ^ x5));
  assign n481 = (x0 | x3 | (x1 ? (~x2 | x4) : (x2 | ~x4))) & (~x3 | ((~x0 | (x1 ? (x2 | x4) : (~x2 | ~x4))) & (x0 | ~x1 | ~x2 | ~x4)));
  assign n482 = x7 ? (((x0 ^ ~x1) | (x2 ? (x3 | ~x4) : (~x3 | x4))) & (x0 | x1 | ~x2 | ~x3 | ~x4) & (~x0 | ~x1 | x2 | x3 | x4)) : (x0 ? (x3 | (~x2 ^ x4)) : (~x3 | ((x1 | x2 | ~x4) & (~x2 | x4))));
  assign z016 = ~n489 | (x1 ? ~n486 : (x2 ? ~n485 : ~n484));
  assign n484 = (x5 | ((~x0 | ((x6 | ~x7 | ~x3 | x4) & (~x6 | x7 | x3 | ~x4))) & (x0 | x3 | x4 | x6 | ~x7))) & (x0 | x3 | x4 | ~x5 | ~x6 | x7);
  assign n485 = (x0 | ((~x5 | x6 | ~x7 | x3 | ~x4) & (x5 | ~x6 | x7 | ~x3 | x4))) & (~x0 | ~x3 | ~x4 | ~x5 | x6 | ~x7);
  assign n486 = (~x6 | n488) & (x4 | ~x5 | x6 | ~n487 | n406);
  assign n487 = ~x0 & x2;
  assign n488 = (x0 | ~x3 | ~x4 | (x2 ? (x5 | ~x7) : (~x5 | x7))) & (~x0 | x2 | x3 | x4 | x5 | x7);
  assign n489 = ~n490 & ~n491 & n492 & (x3 ? n494 : n493);
  assign n490 = ~x0 & ((x3 & (x1 ? ((~x4 & ~x5) | (x2 & x4 & x5)) : (x4 & ~x5))) | (~x1 & ~x2 & ~x3 & x4 & x5));
  assign n491 = ~n390 & (x0 ? ((~x3 & x5 & ~x1 & x2) | (x1 & ~x2 & x3 & ~x5)) : (~x2 & (x1 ? (~x3 & ~x5) : (x3 & x5))));
  assign n492 = ((x1 ^ ~x2) | ((~x0 | (x3 ? (x4 | ~x5) : (~x4 | x5))) & (x4 | ~x5 | x0 | x3))) & (~x0 | ((x1 | x2 | ~x3 | ~x4 | ~x5) & (~x1 | ~x2 | x3 | x4 | x5)));
  assign n493 = ((x0 ? (x1 | x2) : (~x1 | ~x2)) | (x4 ? (x5 | x6) : (~x5 | ~x6))) & ((x1 ^ ~x2) | ((~x5 | ~x6 | x0 | ~x4) & (x5 | x6 | ~x0 | x4))) & (x0 | x1 | x4 | ((x5 | ~x6) & (x2 | ~x5 | x6))) & (~x4 | ~x5 | x6 | ~x0 | ~x1 | x2);
  assign n494 = ((~x0 ^ ~x6) | ((x1 | ((x4 | x5) & (~x2 | ~x4 | ~x5))) & (~x4 | ~x5 | ~x1 | x2))) & (x2 | ((x0 | ~x1 | ~x4 | x5 | ~x6) & (~x0 | x1 | x4 | ~x5 | x6)));
  assign z017 = ~n502 | (x5 ? ~n498 : (x1 ? ~n496 : ~n497));
  assign n496 = x2 ? ((x0 | ~x3 | ~x4 | ~x6 | ~x7) & (~x0 | x3 | x4 | x6 | x7)) : (x6 ? ((x3 | x4 | ~x7) & (~x0 | ((x4 | ~x7) & (x3 | ~x4 | x7)))) : ((x0 | ((x4 | x7) & (x3 | ~x4 | ~x7))) & (~x3 | ((x4 | x7) & (~x0 | ~x4 | ~x7)))));
  assign n497 = (((~x4 | x7) & (~x3 | x4 | ~x7)) | (x0 ? (x2 | x6) : (~x2 | ~x6))) & (x2 | x3 | ((~x0 | ~x6 | (x4 ^ x7)) & (x6 | ((~x4 | x7) & (x0 | x4 | ~x7)))));
  assign n498 = (x3 | n501) & (~x3 | n499) & (n307 | n500);
  assign n499 = (x1 | x2 | ((~x4 | ~x6 | x7) & (x0 | ~x7 | (~x4 ^ x6)))) & (x4 | x6 | ~x7 | x0 | ~x1 | ~x2);
  assign n500 = (x0 | ((~x3 | ~x6 | ~x1 | x2) & (x3 | x6 | x1 | ~x2))) & (~x0 | x1 | ~x2 | ~x3 | x6);
  assign n501 = ((~x4 ^ x7) | ((~x0 | x1 | ~x2 | ~x6) & (x0 | (x1 ? (~x2 | x6) : (x2 | ~x6))))) & (~x2 | ((~x0 | x1 | ~x4 | x6 | ~x7) & (~x6 | x7 | ~x1 | x4)));
  assign n502 = (~x5 | n506) & (x5 | n503) & (n504 | n505);
  assign n503 = (x6 | ((x1 | ~x2 | ~x4) & (x0 | (x1 ? (~x2 | x4) : (~x3 | ~x4))))) & (~x0 | x1 | ~x2 | x4 | ~x6);
  assign n504 = (x2 | ((~x3 | x5 | ~x6) & (~x0 | ((~x5 | ~x6) & (x3 | x5 | x6))))) & (x0 | ((x3 | x5 | ~x6) & (~x2 | ~x3 | ~x5 | x6)));
  assign n505 = ~x1 ^ ~x4;
  assign n506 = x6 ? ((x0 | (x1 ? (x2 ? (~x3 | x4) : (x3 | ~x4)) : (~x2 | ~x4))) & (~x3 | ~x4 | x1 | ~x2)) : ((~x0 | (x1 ? (x3 | x4) : (x2 | ~x4))) & (x2 | (x1 ? x4 : (x3 | ~x4))));
  assign z018 = n508 | ~n514 | (~n425 & ~n513) | (n452 & ~n512);
  assign n508 = ~x1 & ((x4 & ~n510) | (x0 & n509 & n511));
  assign n509 = ~x2 & x3;
  assign n510 = x3 ? ((~x6 | ((~x0 | x7 | (~x2 ^ ~x5)) & (x0 | x2 | ~x5 | ~x7))) & (x0 | x5 | x6 | (x2 ^ x7))) : (~x6 | ((~x0 | ~x7 | (~x2 ^ ~x5)) & (~x5 | x7 | x0 | ~x2)));
  assign n511 = ~x7 & x6 & ~x4 & x5;
  assign n512 = (x5 | ((~x6 | (x0 ? (x2 ? (x3 | x7) : (~x3 | ~x7)) : (x2 ? (~x3 | x7) : (x3 | ~x7)))) & (x0 | x2 | ~x3 | x6 | ~x7))) & (x0 | ~x2 | x3 | ~x5 | ~x6 | ~x7);
  assign n513 = (x4 & ((~x1 & ((~x2 & ~x5) | (~x0 & x3 & x5))) | (x5 & (x2 | (x0 & x1 & ~x3))))) | ((~x0 | x3) & (x2 ^ ~x5)) | (~x3 & ~x4 & x5 & x0 & ~x2) | (~x5 & ((x0 & (x3 ? x1 : x2)) | (x1 & x2 & ~x3 & ~x4)));
  assign n514 = (n515 | n518) & (~x2 | n516) & (x2 | n517);
  assign n515 = x2 ^ ~x4;
  assign n516 = x0 ? (x1 | (x5 ? (x6 | ~x7) : (~x6 | x7))) : ((~x6 | x7 | ~x3 | ~x5) & (x3 | ((~x5 | x6 | ~x7) & (~x6 | x7 | ~x1 | x5))));
  assign n517 = x5 ? ((x0 | x1 | ~x3 | x6 | ~x7) & (~x6 | x7 | ((~x1 | x3) & (~x0 | (~x1 & x3))))) : ((x0 | (x3 ? (~x6 | x7) : (x6 | ~x7))) & (x6 | ~x7 | (x3 ? ~x0 : x1)));
  assign n518 = (x0 | ((~x1 | ~x3 | ~x5 | x6 | ~x7) & (x1 | x3 | x5 | ~x6 | x7))) & (x5 | x6 | ~x7 | ~x0 | ~x1 | x3);
  assign z019 = n521 | n526 | ~n528 | ~n537 | (~n520 & ~n525);
  assign n520 = ~x3 ^ ~x6;
  assign n521 = ~x3 & ((n339 & n524) | (n522 & ~n523));
  assign n522 = ~x2 & x6;
  assign n523 = (x5 | ((x0 | x1 | x4 | x7) & (~x0 | ~x7 | (x1 ^ x4)))) & (x0 | ~x5 | (x1 ? (x4 | x7) : (~x4 | ~x7)));
  assign n524 = x2 & x0 & x1;
  assign n525 = (~x5 | ((x0 | ~x1 | ~x4 | ~x7) & (~x0 | x2 | x4 | x7))) & ((x0 ^ ~x7) | (x1 ? (x2 | ~x4) : (x4 & (~x2 | x5)))) & (x0 | ~x1 | ~x2 | x4 | x5 | x7);
  assign n526 = ~n527 & ~x6 & n358;
  assign n527 = (x1 | (x0 ? (~x7 | (~x4 ^ x5)) : (~x5 | x7))) & (x0 | ~x4 | ~x5 | x7);
  assign n528 = ~n530 & ~n534 & n536 & (n529 | n535);
  assign n529 = x3 ? (~x5 | x6) : (x5 | ~x6);
  assign n530 = ~n533 & (x3 ? (n487 & n312) : (n531 & n532));
  assign n531 = x5 & x6;
  assign n532 = x0 & ~x2;
  assign n533 = x1 ? (x4 | ~x7) : (~x4 | x7);
  assign n534 = ~x0 & ~x1 & x4 & x5 & (x3 ^ ~x6);
  assign n535 = x0 ? (x1 | ~x4) : (~x1 | x4);
  assign n536 = x4 | ~n312 | ((~x0 | ~x1 | x3) & (x0 | x1 | ~x2 | ~x3));
  assign n537 = ~n538 & ~n541 & ~n546 & ~n550 & (x2 | n540);
  assign n538 = ~n539 & ((x0 & ~x1 & ~x4 & x7) | (~x0 & ~x7 & (~x1 ^ x4)));
  assign n539 = x2 ? (x3 | ~x6) : (~x3 | x6);
  assign n540 = (~x0 | ~x1 | ~x6 | (x3 ? (x4 | x5) : (~x4 | ~x5))) & (x0 | x1 | x3 | ~x4 | x5 | x6);
  assign n541 = x4 & n542 & ((n543 & n544) | (n292 & n545));
  assign n542 = x1 & ~x2;
  assign n543 = x6 & ~x7;
  assign n544 = ~x0 & ~x3;
  assign n545 = x0 & x3;
  assign n546 = ~n549 & (x1 ? n548 : n547);
  assign n547 = x4 & x6;
  assign n548 = ~x4 & ~x6;
  assign n549 = (x0 | x2 | ~x3 | x5) & (~x0 | ~x2 | x3 | ~x5);
  assign n550 = ~n551 & (n552 | (n531 & n288));
  assign n551 = x0 ? (x1 | x2) : (~x1 | ~x2);
  assign n552 = ~x6 & ~x5 & x3 & x4;
  assign z020 = n554 | ~n558 | n563 | (x4 ? ~n557 : ~n562);
  assign n554 = ~x3 & ((~x0 & ~n556) | (~n448 & ~n555));
  assign n555 = x4 ? (x6 ^ ~x7) : (x6 | x7);
  assign n556 = (~x5 | x6 | ~x7 | ~x1 | x2 | x4) & (x1 | ((x6 | ((~x2 | ~x4 | x5 | x7) & (x2 | ~x5 | (~x4 ^ ~x7)))) & (x2 | x4 | ~x6 | (x5 ^ x7))));
  assign n557 = x1 ? ((x0 | ((x2 | ~x5 | x7) & (x5 | ~x7 | ~x2 | ~x3))) & (x2 | x7 | (x5 ? ~x3 : ~x0))) : (~x3 | (x2 ? (x5 | x7) : (~x5 | ~x7)));
  assign n558 = (n559 | n560) & (~x3 | ~n487 | n561);
  assign n559 = ~x2 ^ ~x5;
  assign n560 = x1 ? ((x3 | x4 | ~x7) & (x0 | (~x4 ^ x7))) : (x4 ? ~x7 : (x7 | (~x0 & ~x3)));
  assign n561 = (x1 | x6 | (x4 ? (~x5 | x7) : (x5 | ~x7))) & (~x1 | x4 | x5 | ~x6 | ~x7);
  assign n562 = ((x1 ? (~x3 | x5) : (x3 | ~x5)) | (x0 ? (x2 | ~x7) : (~x2 | x7))) & (~x1 | ~x7 | ((~x2 | x3 | x5) & (~x3 | ~x5 | x0 | x2))) & (x1 | x2 | ~x3 | ~x5 | x7);
  assign n563 = ~n564 & ((x0 & ~x6 & (x3 ? (~x4 & x7) : (x4 & ~x7))) | (~x3 & x6 & (~x4 ^ x7)));
  assign n564 = x1 ? (x2 | ~x5) : (~x2 | x5);
  assign z021 = x1 ? ~n568 : (x5 ? ~n566 : ~n567);
  assign n566 = (x2 | ((x0 | ((x6 | ~x7) & (~x4 | ~x6 | x7))) & (~x3 | (~x6 & ~x7)) & (x6 | (x7 ? ~x4 : (~x0 & x3 & x4))))) & (~x3 | ((~x6 | ~x7 | ~x0 | x4) & (x0 | ~x2 | ~x4 | x6 | x7))) & (~x2 | x3 | ((~x6 | (x4 & ~x7)) & (~x0 | (~x6 & (x4 | ~x7)))));
  assign n567 = x2 ? ((~x3 | x6) & ((~x4 & x7) | (~x3 & x6))) : ((~x6 | ~x7 | ~x0 | x4) & (x3 | (~x6 & (x4 | ~x7))));
  assign n568 = n571 & (x3 | n569) & (~x3 | x4 | ~x6 | n570);
  assign n569 = (x6 | ((x7 | ((x0 | ~x2 | x4 | x5) & (~x0 | (x2 ? (~x4 | x5) : (x4 | ~x5))))) & (x4 | ~x7 | (~x2 ^ ~x5)))) & (x0 | ~x4 | ~x5 | ~x6 | (x2 ^ x7));
  assign n570 = (x0 | ~x2 | x5 | x7) & (x2 | ((x5 | ~x7) & (~x0 | ~x5 | x7)));
  assign n571 = (x3 | ~x6 | (x2 ? (x4 | ~x5) : x5)) & (((~x4 | x6) & (~x3 | (~x4 & x6))) | ((x2 | ~x5) & (x0 | ~x2 | x5))) & (x0 | x2 | ~x5 | (~x3 & x6));
  assign z022 = (x5 & ~n577) | (~x5 & ~n573) | (~n425 & ~n576);
  assign n573 = x0 ? n574 : n575;
  assign n574 = (x4 | ((~x1 | ((x2 | ~x3 | x7) & (~x6 | ~x7 | ~x2 | x3))) & (~x3 | x6 | ~x7 | (x1 & x2)))) & (~x6 | x7 | x1 | ~x3) & (~x4 | ((x3 | x6 | x7) & ((x1 & x2) | (x3 ^ x6))));
  assign n575 = (~x4 | (x3 ^ x6)) & (~x3 | ((x4 | x6 | ~x7) & (~x6 | ((x1 | x2) & x7))));
  assign n576 = (x0 | ((~x4 | ~x5 | x1 | ~x3) & (x4 | x5 | ~x2 | x3))) & (x3 | x4 | ((~x1 | (x5 ? ~x0 : x2)) & (x1 | ~x2 | x5) & (~x0 | (~x2 ^ ~x5))));
  assign n577 = ~n579 & n581 & (n392 | n578) & (n437 | n580);
  assign n578 = (~x0 | x1 | x2 | x4 | x6) & (x0 | ~x1 | ((~x4 | ~x6) & (~x2 | x4 | x6)));
  assign n579 = ~x0 & x1 & ((~x3 & x4 & ~x6) | (~x4 & x6 & x2 & x3));
  assign n580 = (~x0 | ~x3 | x4 | (x1 ^ ~x2)) & (x0 | x1 | x3 | ~x4);
  assign n581 = (x1 & (x2 | (x0 & ~x4))) | (x0 & ~x4 & (x2 | ~x6)) | (x3 & ~x6) | (~x3 & x6) | (~x0 & x4);
  assign z023 = n584 | ~n587 | (~x2 & ~n583);
  assign n583 = x0 ? ((~x1 | ~x3 | ~x4 | x5 | ~x7) & (~x5 | x7 | x1 | x4)) : ((x4 | ~x5 | ~x7) & (x1 | x7 | ((~x4 | ~x5) & (~x3 | x4 | x5))));
  assign n584 = ~x7 & ((~x2 & ~n586) | (x2 & x5 & n349 & ~n585));
  assign n585 = ~x4 ^ ~x6;
  assign n586 = (x3 | x5 | ((x0 | x1 | x4 | ~x6) & (~x0 | ~x1 | ~x4 | x6))) & (x0 | ~x1 | ~x5 | (x4 ^ x6));
  assign n587 = (~n588 | n592) & (n307 | n591) & (n589 | n590);
  assign n588 = x2 & x5;
  assign n589 = x4 ^ ~x6;
  assign n590 = (~x7 | ((x0 | (x1 ? (~x2 | ~x5) : (x2 | x5))) & (~x0 | x1 | x2 | ~x5))) & (~x0 | ~x1 | x5 | x7 | (~x2 ^ x3));
  assign n591 = (x0 & x1 & (x2 | (x3 & ~x5))) | (~x1 & ~x2 & x5) | (~x0 & (x5 | (~x1 & ~x2)));
  assign n592 = (~x0 | ~x1 | x3 | x4 | x7) & (x0 | x1 | (~x4 ^ x7));
  assign z024 = ~n598 | (x3 ? ~n597 : ~n594);
  assign n594 = (x5 | n596) & (~x5 | x6 | x7 | n515 | ~n595);
  assign n595 = x0 & x1;
  assign n596 = (~x4 | (~x2 ^ ~x7) | (x0 ? (x1 | ~x6) : (~x1 | x6))) & (~x0 | ~x1 | x4 | (~x2 ^ (~x6 & ~x7)));
  assign n597 = (x5 | (~x2 ^ ~x7) | (x0 ? (x1 | ~x6) : (~x1 | x6))) & (~x5 | x6 | x7 | ~x0 | ~x1 | x2);
  assign n598 = x0 ? ((x2 | ((~x6 | ~x7 | x1 | ~x5) & (x5 | (x6 ? ~x1 : ~x7)))) & (x1 | x5 | (x6 & (~x2 | x7)))) : ((~x1 | ((~x5 | ~x6) & (x6 | x7 | ~x2 | x5))) & (x1 | ((~x5 | x6) & (~x6 | ~x7 | x2 | x5))) & (~x5 | ((x2 | x6 | ~x7) & (~x6 | (~x2 & x7)))));
  assign z025 = n601 | ~n603 | (~x3 & (~n600 | (~x4 & ~n602)));
  assign n600 = (x6 | ((~x0 | ((~x4 | ~x7 | x1 | ~x2) & (~x1 | x4 | (~x2 ^ ~x7)))) & (x1 | x2 | ~x4 | x7))) & (~x0 | ~x1 | ~x6 | x7 | (~x2 ^ x4));
  assign n601 = (~x1 | (~x2 & (~x6 | ~x7))) & (x1 | (x6 ? x7 : x2)) & (x2 | x6 | x7) & (~x2 | ~x6) & (~x0 | x3);
  assign n602 = (x0 | x1 | x2 | ~x5 | x6 | x7) & (x5 | (~x2 ^ ~x7) | (x0 ? (x1 | ~x6) : (~x1 | x6)));
  assign n603 = x1 ? ((x0 | ~x2 | ~x6) & (x3 | x6 | ~x7 | ~x0 | x2)) : ((x6 | x7 | x2 | ~x3) & (~x0 | x3 | (x2 ? (x6 | x7) : (~x6 | ~x7))));
  assign z026 = n605 | ~n608 | (n288 & (~n606 | ~n607));
  assign n605 = ~x3 & ((x0 & ((x4 & ((~x2 & x7) | (~x1 & x2 & ~x7))) | (x1 & ~x4 & (x2 ^ ~x7)))) | (x2 & x4 & ~x7 & ~x0 & x1));
  assign n606 = (x6 | (~x2 ^ ~x7) | (x0 ? (x1 | ~x5) : (~x1 | x5))) & (~x5 | ~x6 | x7 | ~x0 | x1 | ~x2);
  assign n607 = (~x2 | ((~x0 | x1 | x5 | ~x7) & (x0 | ~x1 | ~x5 | x7))) & (~x0 | x1 | x2 | (x5 ^ x7));
  assign n608 = (x0 & (~x3 | (x1 & ~x7))) | (x2 & x7) | (~x7 & (~x2 | (x1 & ~x3)));
  assign z027 = (~x4 | ~n610) & (n618 | ~n619 | x4 | n614);
  assign n610 = x3 ? n613 : ((~n317 | ~n611) & (~n524 | ~n612));
  assign n611 = x7 & x5 & x6;
  assign n612 = ~x7 & ~x5 & ~x6;
  assign n613 = x0 & x1 & (x2 | (~x5 & ~x6 & ~x7));
  assign n614 = ~n617 & (x3 ? (n321 & n615) : (n349 & n616));
  assign n615 = x5 & x7;
  assign n616 = ~x5 & ~x7;
  assign n617 = ~x2 ^ ~x6;
  assign n618 = (x2 ? (~x3 & ~x6) : (x3 & x6)) & (x0 ? (~x1 & x5) : (x1 & ~x5));
  assign n619 = x3 ? (x0 | (x1 & ~x5)) : (~x0 | (~x1 & x5 & (x2 | ~n372)));
  assign z028 = ~n626 | (x0 ? ~n623 : (n622 | (x6 & ~n621)));
  assign n621 = (x4 | ~x5 | x7 | x1 | x2 | x3) & (~x7 | ((x1 | x2 | ~x3 | ~x4 | ~x5) & (~x1 | ~x2 | x5 | (~x3 ^ x4))));
  assign n622 = n312 & (x3 ? (n542 & n370) : (n354 & n369));
  assign n623 = (~x5 | n624) & (~x1 | x5 | n625);
  assign n624 = (~x1 | ~x2 | x3 | x4) & (x1 | ((x2 | x3 | ~x4 | x6 | ~x7) & (~x2 | ~x3 | x4 | ~x6 | x7)));
  assign n625 = (~x4 | x6 | x7 | (x2 ^ ~x3)) & (~x2 | x3 | x4 | (~x6 & ~x7));
  assign n626 = n630 & n631 & (x1 | n628) & (~n627 | ~n629);
  assign n627 = ~x5 & ~x4 & ~x0 & x1;
  assign n628 = (x5 | x6 | ~x7 | x0 | ~x2 | ~x4) & (~x5 | (x0 ? ((~x2 | ~x4 | ~x6 | ~x7) & (x2 | x4 | x6 | x7)) : (x2 | ~x6 | (~x4 ^ x7))));
  assign n629 = ~x7 & (x2 ^ ~x6);
  assign n630 = ((x2 ? (x4 | x6) : (~x4 | ~x6)) | (x0 ? (x1 | ~x5) : (~x1 | x5))) & (x0 | x1 | ~x4 | (x2 ? (x5 | ~x6) : (~x5 | x6)));
  assign n631 = x0 ? (x4 | (x1 ? x2 : x5)) : (~x4 | ((x1 | x2 | x5) & (~x5 | (~x1 & ~x2))));
  assign z029 = ~n638 | (x0 ? ~n635 : (x2 ? ~n633 : ~n634));
  assign n633 = (x1 | ~x3 | ~x4 | x5 | x6 | x7) & (~x1 | x3 | x4 | ~x5 | ~x6 | ~x7);
  assign n634 = (~x5 | (x1 ? (x4 | (x3 ? (~x6 | x7) : (x6 | ~x7))) : (~x4 | ~x6 | (x3 ^ x7)))) & (x3 | x5 | ((~x6 | x7 | x1 | x4) & (x6 | ~x7 | ~x1 | ~x4)));
  assign n635 = (~x5 | n636) & (x2 | x5 | x6 | n637);
  assign n636 = x1 ? (x4 | ((~x2 | x3 | (~x6 & ~x7)) & (x6 | x7 | x2 | ~x3))) : (~x4 | ((x6 | ~x7 | x2 | ~x3) & (~x6 | x7 | ~x2 | x3)));
  assign n637 = (x1 | x4 | (~x3 ^ ~x7)) & (~x1 | ~x3 | ~x4 | x7);
  assign n638 = ~n639 & ~n640 & ~n642 & n643 & (x2 | n641);
  assign n639 = x3 & n354 & ((x0 & x6 & (x5 ^ x7)) | (~x6 & x7 & ~x0 & x5));
  assign n640 = ~x3 & (x0 ? ((~x5 & x6 & ~x1 & x2) | (x5 & ~x6 & x1 & ~x2)) : (x5 & (x1 ? (~x2 & x6) : (x2 & ~x6))));
  assign n641 = (x0 | x5 | ((~x6 | ~x7 | x1 | ~x3) & (x6 | x7 | ~x1 | x3))) & (~x5 | x6 | x7 | ~x0 | x1 | x3);
  assign n642 = ~n368 & (x1 ? ((x5 & x7 & ~x2 & x3) | (~x5 & ~x7 & x2 & ~x3)) : (~x2 & (x3 ? (x5 & ~x7) : (~x5 & x7))));
  assign n643 = x0 ? ((x1 | (x2 ? (~x5 | x6) : (x5 | ~x6))) & (~x5 | ~x6 | ~x1 | x2)) : (x1 ? (x5 | ((~x3 | x6) & (~x2 | (~x3 & x6)))) : (~x5 | (~x2 ^ ~x6)));
  assign z030 = (~x0 & (~n646 | (~x3 & ~n645))) | ~n651 | (~x3 & ~n650);
  assign n645 = (x6 | ((~x1 | ~x5 | (x2 ? (~x4 | ~x7) : (x4 | x7))) & (x1 | x2 | x4 | x5 | ~x7))) & (x5 | ~x6 | x7 | x1 | x2 | ~x4);
  assign n646 = (~x6 | x7 | n648) & (~x7 | ((~n647 | n649) & (x6 | n648)));
  assign n647 = ~x1 & x3;
  assign n648 = ((x4 & x5) | (x1 ? (~x2 | x3) : (x2 | ~x3))) & (x2 | ~x4 | ~x5 | (~x1 ^ ~x3));
  assign n649 = (~x2 | x4 | x5 | ~x6) & (x2 | ~x4 | ~x5 | x6);
  assign n650 = (x1 | ((x5 | ((~x0 | (x2 ? (~x4 | x6) : (x4 | ~x6))) & (~x4 | x6 | x0 | x2))) & (x4 | ~x5 | x6 | x0 | x2))) & (x0 | ~x1 | ~x2 | ~x4 | ~x5 | ~x6);
  assign n651 = ~n656 & n657 & (n425 | n652) & (~x0 | n653);
  assign n652 = x1 ? ((x0 | x2 | x3 | x4 | x5) & (~x0 | (x2 ? (x3 | x4) : (~x3 | ~x4)))) : ((~x3 | (x0 ? (x2 | x4) : (~x2 | (~x4 & ~x5)))) & (~x0 | x2 | (x4 ? x3 : ~x5)));
  assign n653 = x1 ? n655 : (~x2 | n437 | (~x3 & ~n654));
  assign n654 = x4 & x5;
  assign n655 = (x2 | ~x3 | x4 | ~x5 | ~x6 | ~x7) & (~x2 | x3 | ~x4 | x5 | x6 | x7);
  assign n656 = n509 & ((x0 & x1 & ~x4 & ~x5 & x6) | (~x0 & x4 & (x1 ? (~x5 & ~x6) : (x5 & x6))));
  assign n657 = x2 ? ((x0 | ~x6 | (~x1 ^ ~x3)) & (~x0 | x1 | x3 | x4 | x6)) : (x0 ? ((~x1 | x3 | ~x6) & (~x4 | x6 | x1 | ~x3)) : (~x1 | x6 | (~x3 ^ x4)));
  assign z031 = ~n659 | n663 | ~n669 | (x2 & ~n666);
  assign n659 = (n406 | n661) & (x2 | (n660 & n662));
  assign n660 = ((x4 ^ x7) | (x0 ? (x1 | ~x3) : (~x1 | x3))) & (~x0 | x3 | (x1 ? (x4 | ~x7) : (~x4 | x7))) & (x0 | ~x1 | ~x3 | x4 | ~x7);
  assign n661 = x0 ? (x1 ? (x2 | ~x4) : (~x2 | x4)) : (x1 | (x2 ^ x4));
  assign n662 = ((x1 ^ x3) | ((x5 | ~x7 | ~x0 | x4) & (~x5 | x7 | x0 | ~x4))) & (x1 | x7 | ((x0 | ~x3 | ~x4 | x5) & (x4 | ~x5 | ~x0 | x3)));
  assign n663 = n354 & ((~x0 & x3 & ~x4 & n664) | (x0 & ~x3 & x4 & ~n665));
  assign n664 = x5 & ~x7;
  assign n665 = x5 ^ ~x7;
  assign n666 = (~x1 | x3 | ~x4 | n667) & (x0 | x1 | ~x3 | x4 | ~n668);
  assign n667 = (~x0 | x5 | x6 | x7) & (~x6 | ~x7 | x0 | ~x5);
  assign n668 = ~x5 & (~x6 ^ ~x7);
  assign n669 = ~n670 & (x2 | ((n671 | n672) & (x0 | n673)));
  assign n670 = x2 & (x1 ? ((~x3 & ~x4 & ~x7) | (~x0 & (~x3 ^ x7))) : ((~x4 & x7 & ~x0 & ~x3) | (x4 & ~x7 & x0 & x3)));
  assign n671 = x3 ? (~x5 | ~x6) : (x5 | x6);
  assign n672 = (~x0 | ~x1 | x4 | x7) & (x0 | x1 | ~x4 | ~x7);
  assign n673 = x1 ? (~x7 | ((~x3 | ~x4 | x5 | x6) & (~x5 | ~x6 | x3 | x4))) : (~x4 | x7 | (x3 ? (~x5 | x6) : (x5 | ~x6)));
  assign z032 = n676 | n680 | ~n681 | (x3 ? ~n679 : ~n675);
  assign n675 = (~x0 | ((x2 | ((~x5 | x6 | x1 | ~x4) & (~x1 | x5 | (~x4 ^ x6)))) & (x1 | ~x2 | x4 | x5 | x6))) & (~x4 | x5 | ~x6 | x0 | x1 | x2);
  assign n676 = x1 & ((~x0 & ~n677) | (n532 & ~n399 & ~n678));
  assign n677 = ((x4 ? (~x6 | ~x7) : (x6 | x7)) | (x2 ? (x3 | ~x5) : (~x3 | x5))) & (x2 | x3 | x4 | ~x5 | ~x6 | ~x7);
  assign n678 = x4 ? (~x6 | x7) : (x6 | ~x7);
  assign n679 = x0 ? (~x5 | ((x4 | x6 | x1 | ~x2) & (~x1 | x2 | (~x4 ^ x6)))) : ((x1 | ~x6 | (x2 ? (x4 | x5) : (~x4 | ~x5))) & (~x1 | ~x2 | ~x4 | x5 | x6));
  assign n680 = ~x1 & (((x3 ? (~x4 & ~x5) : (x4 & x5)) & (x0 ^ ~x2)) | ((~x3 ^ x5) & (x0 ? (~x2 & x4) : (x2 & ~x4))));
  assign n681 = n682 & ((x4 & (x2 | (x3 & ~x5))) | ~n349 | (~x4 & (~x2 | (~x3 & x5))));
  assign n682 = (~x0 | ((x2 | n683) & (~x3 | ~n511 | x1 | ~x2))) & (x0 | x1 | ~x2 | n683);
  assign n683 = x3 ? (~x4 | x5) : (x4 | ~x5);
  assign z033 = ~n690 | (x5 ? ~n688 : ~n685);
  assign n685 = (x2 | n687) & (~n543 | ~n686 | ~n288);
  assign n686 = x2 & ~x0 & ~x1;
  assign n687 = x0 ? ((x3 | ((~x1 | ~x7 | (x4 ^ x6)) & (x6 | x7 | x1 | ~x4))) & (x4 | ~x6 | x7 | x1 | ~x3)) : ((~x3 | ((~x1 | ~x7 | (x4 ^ x6)) & (x6 | x7 | x1 | ~x4))) & (x4 | x6 | ~x7 | x1 | x3));
  assign n688 = (~x6 | n689) & (n533 | ((~x0 | x2 | ~x3 | x6) & (x0 | x3 | (x2 ^ ~x6))));
  assign n689 = (~x2 | ((x1 | x4 | (x0 ? (x3 ^ x7) : (~x3 | x7))) & (x0 | ~x1 | ~x4 | (~x3 ^ x7)))) & (~x3 | ~x4 | ~x7 | ~x0 | ~x1 | x2);
  assign n690 = n693 & (x2 ? n692 : n691);
  assign n691 = x0 ? (x1 ? (x3 ? (x4 ? (x5 | x6) : (~x5 | ~x6)) : (x4 | (~x5 ^ x6))) : ((x5 | x6 | ~x3 | x4) & (~x5 | ~x6 | x3 | ~x4))) : (((~x3 ^ ~x6) | (x1 ? (x4 | x5) : (~x4 | ~x5))) & (~x1 | ~x3 | x4 | ~x5 | x6) & (x5 | ~x6 | x1 | x3));
  assign n692 = ((~x5 ^ x6) | ((~x0 | x1 | x3 | x4) & (x0 | ~x3 | (~x1 ^ ~x4)))) & (~x0 | x1 | ~x3 | x4 | x5 | x6) & (x0 | x3 | ((~x1 | (x4 ? (x5 | x6) : (~x5 | ~x6))) & (x5 | x6 | x1 | x4)));
  assign n693 = ((x1 ? (x2 ? (x4 | x5) : (~x4 | ~x5)) : (~x5 | (x2 ^ x4))) | (x0 ^ ~x3)) & (~x4 | x5 | (x0 ? (x1 | ~x3) : (x3 | (x1 ^ ~x2))));
  assign z034 = ~n710 | ~n707 | n706 | n704 | n695 | ~n698;
  assign n695 = ~x2 & ((~x5 & ~n696) | (~x0 & n273 & n697));
  assign n696 = ((~x6 ^ x7) | ((~x0 | x1 | x3 | ~x4) & (x0 | ~x1 | ~x3 | x4))) & (x4 | x6 | ((x0 | x1 | (~x3 ^ x7)) & (~x0 | ~x1 | x3 | ~x7)));
  assign n697 = x7 & x6 & x4 & x5;
  assign n698 = (n699 | n703) & (n683 | n702) & (n700 | n701);
  assign n699 = x4 ^ ~x7;
  assign n700 = x3 ? (x4 | x7) : (~x4 | ~x7);
  assign n701 = (~x0 | ~x1 | x2 | x5 | ~x6) & (x0 | ~x2 | ~x5 | (~x1 ^ ~x6));
  assign n702 = (x0 | x2 | ~x6 | (~x1 ^ ~x7)) & (~x0 | x1 | ~x2 | x6 | x7);
  assign n703 = ((x1 ? (~x5 | x6) : (x5 | ~x6)) | (x0 ? (x2 | ~x3) : (~x2 | x3))) & (x1 | ~x2 | ~x5 | ~x6 | (x0 ^ ~x3));
  assign n704 = ~n705 & (x2 ? ((~x0 & (x3 ? ~x6 : (x5 & x6))) | (~x3 & ~x6 & (x0 | ~x5))) : ((x0 & ((x5 & x6) | (x3 & ~x5 & ~x6))) | (x6 & ((x3 & x5) | (~x0 & ~x3 & ~x5)))));
  assign n705 = x1 ^ ~x4;
  assign n706 = (x2 ? (~x5 & x6) : (x5 & ~x6)) & (x0 ? (~x1 & ~x4) : (x1 & x4));
  assign n707 = n709 & (n708 | ((x0 | x1 | ~x2 | x4) & (~x0 | ~x1 | x2 | ~x4)));
  assign n708 = x3 ? (x5 | ~x6) : (~x5 | x6);
  assign n709 = ~n451 | ((x4 | ~n317) & (~x3 | ~x4 | ~n459));
  assign n710 = (n712 | n713) & (n711 | (x1 ? (x3 | x7) : (~x3 | ~x7)));
  assign n711 = (~x0 | ~x2 | x4 | ~x5 | ~x6) & (x0 | x2 | ~x4 | x5 | x6);
  assign n712 = (x3 | x4 | x5 | x7) & (~x3 | ~x4 | ~x5 | ~x7);
  assign n713 = (~x2 | ~x6 | x0 | ~x1) & (~x0 | x2 | (~x1 ^ ~x6));
  assign z035 = ~n716 | n723 | (~x1 & ~n715) | (~n416 & ~n722);
  assign n715 = x2 ? ((x4 | x5 | ~x7 | x0 | x3) & (~x4 | ~x5 | x7 | ~x0 | ~x3)) : (((x0 ^ ~x3) | ((~x5 | x7) & (~x4 | x5 | ~x7))) & (x4 | ~x7 | (x0 ? (~x3 | x5) : (x3 | ~x5))));
  assign n716 = ~n720 & (x2 | (~n717 & n718 & (~x1 | n721)));
  assign n717 = ~n705 & (((~x6 ^ x7) & (x0 ? (x3 & ~x5) : (~x3 & x5))) | (x0 & x3 & x5 & ~x6 & x7) | (~x0 & ~x3 & ~x5 & x6 & ~x7));
  assign n718 = (x0 | x1 | x3 | ~n719) & (~x0 | ~x1 | ~x3 | ~n351 | ~n374);
  assign n719 = ~x4 & ~x7 & (~x5 ^ ~x6);
  assign n720 = ~n440 & ((x1 & x4 & (x0 ? (~x2 & x3) : (x2 & ~x3))) | (x2 & (~x1 | ~x4) & (~x0 ^ ~x3)));
  assign n721 = (x0 | x3 | ~x4 | ~x5 | x7) & ((x0 ^ ~x3) | ((x5 | ~x7) & (x4 | ~x5 | x7)));
  assign n722 = x1 ? (x2 | ~x4 | (x0 ? (x3 | x7) : (~x3 ^ x7))) : ((x4 | ((x2 | (x0 ? (~x3 ^ x7) : (~x3 | ~x7))) & (x3 | x7 | x0 | ~x2))) & (~x0 | ~x2 | ~x3 | ~x4 | ~x7));
  assign n723 = x2 & ((~n425 & ~n724) | n725 | ~n726);
  assign n724 = (x0 | ((~x1 | (x3 ? (~x4 | ~x5) : (x4 | x5))) & (x1 | x3 | ~x4 | x5))) & (~x0 | x1 | ~x3 | x4 | ~x5);
  assign n725 = ~n406 & ((x0 & ~x1 & ~x4 & n450) | (~x0 & (x1 ? (x4 ? n450 : n451) : (x4 & n451))));
  assign n726 = (~x0 | x3 | ~n451 | ~n727) & (x0 | x1 | ~x3 | ~n352);
  assign n727 = ~x7 & (~x1 ^ ~x4);
  assign z036 = n730 | ~n732 | (x6 ? ~n729 : ~n731);
  assign n729 = x0 ? ((~x4 | x7 | (x1 ? (x2 | ~x3) : (x2 ^ x3))) & (~x1 | x3 | x4 | (x2 & ~x7))) : ((x2 | (x1 ? (~x3 | x4) : (x3 ? (~x4 | x7) : (x4 | ~x7)))) & (~x1 | (x3 ? (x4 | ~x7) : (~x4 | x7))));
  assign n730 = ~n307 & ((~x1 & (x0 ? (x3 ^ x6) : ((x3 & x6) | (x2 & ~x3 & ~x6)))) | (~x0 & x1 & ~x2 & ~x3 & ~x6));
  assign n731 = (x2 | ((~x0 | (x1 ? (x3 ? x4 : (~x4 | x7)) : (x3 ? (~x4 | x7) : (x4 | ~x7)))) & (x0 | x1 | ~x3 | x4 | ~x7))) & (x0 | ((~x4 | x7 | x1 | x3) & (~x1 | ((~x3 | ~x4 | x7) & (~x2 | x3 | x4)))));
  assign n732 = x5 ? (~n734 & ~n735 & (x3 | n733)) : n737;
  assign n733 = x0 ? (~x2 | ((x6 | x7 | ~x1 | x4) & (x1 | (x4 ? (x6 | x7) : (~x6 | ~x7))))) : ((x4 | x6 | ~x7 | ~x1 | x2) & (~x4 | ~x6 | x7 | x1 | ~x2));
  assign n734 = ~n307 & ((x0 & x1 & ~x2 & x3 & x6) | (~x0 & ((x1 & x2 & (x3 ^ x6)) | (~x3 & ~x6 & ~x1 & ~x2))));
  assign n735 = n647 & (x0 ? ~n736 : (x2 & ~n390));
  assign n736 = (~x2 | x4 | x6 | ~x7) & (x2 | ~x4 | ~x6 | x7);
  assign n737 = (~x0 | (n738 & (x3 | n739))) & (n740 | ~n741) & (x0 | ~x3 | n739);
  assign n738 = (~x4 | x6 | ((~x1 | (x2 ? (x3 | x7) : (~x3 | ~x7))) & (x1 | ~x2 | ~x3 | x7))) & (x4 | ~x6 | ~x7 | x1 | x2 | ~x3);
  assign n739 = (~x6 | ((~x1 | (x2 ? (x4 | x7) : (~x4 | ~x7))) & (x1 | ~x2 | ~x4 | x7))) & (x1 | x4 | x6 | (~x2 ^ ~x7));
  assign n740 = x1 ? (~x4 | x6) : (x4 | ~x6);
  assign n741 = ~x0 & ~x3 & (x2 ^ ~x7);
  assign z037 = (~x3 & ~n743) | (~n425 & ~n746) | ~n751 | (x3 & ~n747);
  assign n743 = x1 ? n744 : n745;
  assign n744 = (x7 | ((x0 | ~x6 | (x2 ? (x4 | ~x5) : (~x4 | x5))) & (~x0 | ~x2 | ~x4 | x5 | x6))) & (~x0 | x4 | x6 | ~x7 | (x2 ^ ~x5));
  assign n745 = x0 ? ((x2 | ((x6 | ~x7 | ~x4 | ~x5) & (~x6 | x7 | x4 | x5))) & (~x2 | ~x4 | x5 | x6 | ~x7)) : ((x5 | x6 | ~x7 | x2 | x4) & (~x2 | ~x4 | ~x5 | ~x6 | x7));
  assign n746 = x3 ? ((~x2 ^ x5) | (x0 ? (x1 | x4) : (~x1 | ~x4))) : ((x0 | x1 | ~x2 | x4 | ~x5) & (x2 | ((x0 | x5 | (x1 ^ ~x4)) & (~x0 | ~x1 | ~x4 | ~x5))));
  assign n747 = ~n749 & (~n748 | ~n543 | (x0 ? (~x1 | ~x5) : (x1 | x5)));
  assign n748 = ~x2 & ~x4;
  assign n749 = ~n750 & ((x0 & ~x1 & x4 & x6 & ~x7) | (~x0 & ~x6 & x7 & (~x1 ^ ~x4)));
  assign n750 = x2 ^ ~x5;
  assign n751 = n754 & (x1 | n752) & (n699 | n753);
  assign n752 = (x5 | (x0 ^ ~x2) | (x3 ? (x4 | x7) : (~x4 | ~x7))) & (x2 | ~x5 | ((x0 | ((x4 | x7) & (x3 | ~x4 | ~x7))) & (x3 | x4 | x7)));
  assign n753 = ((~x0 & ~x3) | (x1 ? (x2 | x5) : (~x2 | ~x5))) & (x0 | ~x1 | x3 | (~x2 ^ x5));
  assign n754 = (~x3 | ((x4 | x7 | ~n756) & (x2 | ~x4 | ~x7 | n755))) & (~x4 | ~x7 | ~n756) & (~x2 | x3 | x4 | x7 | n755);
  assign n755 = (x1 | x5) & (~x0 | ~x1 | ~x5);
  assign n756 = x5 & x2 & ~x0 & x1;
  assign z038 = n758 | ~n760 | (n345 & ~n766) | (x0 & ~n765);
  assign n758 = x1 & ((n284 & n342) | (x6 & ~n759));
  assign n759 = x0 ? ((x4 | x5 | ~x7 | ~x2 | x3) & (~x4 | ~x5 | x7 | x2 | ~x3)) : (~x2 | ((~x5 | x7 | x3 | ~x4) & (x5 | ~x7 | ~x3 | x4)));
  assign n760 = n762 & ~n763 & ~n764 & (x0 | n761);
  assign n761 = ((~x4 ^ x6) | ((~x1 | ~x2 | x3 | ~x5) & (x1 | x2 | ~x3 | x5))) & ((x4 ? (x5 | ~x6) : (~x5 | x6)) | (x1 ? (~x2 | ~x3) : (x2 | x3))) & (~x1 | x2 | ~x3 | ~x4 | ~x5 | ~x6) & (x1 | ~x2 | x3 | x4 | x5 | x6);
  assign n762 = ((x1 ? (x2 | x5) : (~x2 | ~x5)) | (x0 ? (x3 | x6) : (~x3 ^ x6))) & (~x0 | x1 | ~x3 | ~x6 | (~x2 ^ x5));
  assign n763 = ~n443 & ((~x0 & x1 & ~x2 & ~x3 & ~x6) | (~x1 & x2 & (x0 ? (x3 ^ x6) : (x3 & x6))));
  assign n764 = ~n440 & ~n705 & ((~x0 & x2 & ~x3 & ~x6) | (~x2 & (x0 ? (x3 ^ x6) : (x3 & x6))));
  assign n765 = (x2 | (((~x4 ^ x6) | (x1 ? (~x3 | ~x5) : (x3 | x5))) & (~x1 | x3 | ~x4 | ~x5 | ~x6) & (x1 | ~x3 | x4 | x5 | x6))) & (x4 | ~x5 | x6 | ~x1 | ~x2 | x3);
  assign n766 = (x5 | x6 | ~x7 | ~x0 | x3 | x4) & (x0 | ((x5 | x6 | ~x7 | ~x3 | x4) & (x3 | ((~x6 | ~x7 | x4 | x5) & (~x4 | ~x5 | x6 | x7)))));
  assign z039 = ~n771 | n776 | (x2 ? ~n768 : (n779 | ~n782));
  assign n768 = ~n770 & (n437 | n724) & (x1 | n389 | n769);
  assign n769 = x0 ? (~x3 | x5) : (x3 | ~x5);
  assign n770 = n349 & (x5 ? (n292 & n288) : (n543 & n361));
  assign n771 = (n774 | ~n775) & (n425 | n772) & (x1 | n773);
  assign n772 = x0 ? ((~x5 | ((~x3 | ~x4 | ~x1 | x2) & (x3 | x4 | x1 | ~x2))) & (x3 | (x2 & x5) | (x1 ^ ~x4))) : ((~x2 | ~x5 | (x1 ? (x3 | ~x4) : (~x3 | x4))) & (~x3 | (x2 & x5) | (x1 ^ ~x4)));
  assign n773 = x0 ? (~x3 | ((x5 | ~x6 | x2 | x4) & (~x5 | x6 | ~x2 | ~x4))) : (x3 | x4 | ~x6 | (x2 ^ ~x5));
  assign n774 = (~x0 | x2 | ~x3 | x5) & (x0 | x3 | (x2 ^ ~x5));
  assign n775 = ~x6 & x1 & x4;
  assign n776 = ~n777 & (x6 ? ~n778 : (n384 & ~n750));
  assign n777 = x0 ^ ~x3;
  assign n778 = (~x4 | ~x5 | x1 | ~x2) & (~x1 | (x2 ? (x4 | ~x5) : (~x4 | x5)));
  assign n779 = ~n777 & (x1 ? (x4 & n781) : (~x4 & n780));
  assign n780 = x7 & ~x5 & ~x6;
  assign n781 = ~x7 & x5 & x6;
  assign n782 = ~n787 & n785 & (~x6 | ~n783 | ~n784 | n699);
  assign n783 = ~x0 & ~x1;
  assign n784 = ~x3 & ~x5;
  assign n785 = (~x0 | ~n367 | ~n786) & (n437 | n705 | n769);
  assign n786 = x7 & ~x6 & ~x4 & x5;
  assign n787 = ~n389 & (x3 ? (x5 & n321) : (~x5 & n349));
  assign z041 = n789 | n795 | ~n799 | (x2 ? ~n793 : ~n794);
  assign n789 = ~x0 & (~n791 | (~x7 & ~n790));
  assign n790 = (~x2 | ((~x4 | ((~x1 | x6 | (x3 ^ x5)) & (~x5 | ~x6 | x1 | ~x3))) & (x1 | x4 | x5 | (~x3 ^ x6)))) & (x1 | x2 | x4 | ~x5 | (~x3 ^ x6));
  assign n791 = (x2 | ~x7 | n792) & (n708 | ((~x4 | ~x7 | x1 | ~x2) & (~x1 | (x2 ? (x4 | ~x7) : (~x4 | x7)))));
  assign n792 = x1 ? ((~x5 | ~x6 | ~x3 | x4) & (x5 | x6 | x3 | ~x4)) : ((~x3 | (x4 ? (~x5 | ~x6) : (x5 | x6))) & (x3 | x4 | x5 | ~x6));
  assign n793 = (x4 | ~x5 | x6 | ~x0 | ~x1 | x3) & (x0 | ((x4 | ~x5 | ~x6 | x1 | ~x3) & (~x1 | (x3 ? (x4 ? (x5 | ~x6) : (~x5 | x6)) : (x6 | (x4 ^ x5))))));
  assign n794 = ((~x3 ^ x6) | ((~x0 | (x1 ? (~x4 | ~x5) : (x4 | x5))) & (x0 | x1 | ~x4 | x5))) & (~x0 | ((~x1 | ~x3 | x4 | ~x5 | ~x6) & (x1 | x3 | ~x4 | x5 | x6))) & (x0 | ~x1 | ((~x5 | x6 | x3 | x4) & (~x3 | ~x6 | (x4 ^ x5))));
  assign n795 = x0 & (n796 | n797 | (x1 & x6 & ~n442));
  assign n796 = n268 & n269;
  assign n797 = ~n798 & ((~x2 & ~n440 & ~n705) | (~x1 & x2 & ~n443));
  assign n798 = x3 ^ ~x6;
  assign n799 = x0 ? ((x1 | ((~x5 | ~x6 | x2 | ~x3) & (~x2 | (x3 ? (x5 | ~x6) : (~x5 | x6))))) & (~x1 | x2 | x3 | x5 | x6)) : (x2 ? ((x3 | ~x5 | ~x6) & (x1 | x6 | (x3 ^ x5))) : ((~x5 | x6 | x1 | x3) & (x5 | (x1 ? (~x3 ^ x6) : (~x3 | ~x6)))));
  assign z042 = ~n807 | (x2 ? (x5 ? ~n801 : ~n802) : ~n803);
  assign n801 = ((~x6 ^ x7) | ((~x0 | x1 | ~x3 | x4) & (x0 | (x1 ? (x3 ^ x4) : (x3 | ~x4))))) & (x0 | ~x1 | ~x3 | x4 | x6 | x7) & (x1 | x3 | ((~x0 | (x4 ? (x6 | x7) : (~x6 | ~x7))) & (x6 | x7 | x0 | x4)));
  assign n802 = (x0 | ((x4 | x6 | ~x7 | x1 | ~x3) & (~x1 | x3 | (x4 ? (x6 | ~x7) : (~x6 | x7))))) & (x1 | ~x3 | ((x4 | ~x6 | x7) & (x6 | ~x7 | ~x0 | ~x4)));
  assign n803 = x6 ? (n806 & (x7 | n804)) : (n805 & (~x7 | n804));
  assign n804 = x0 ? ((~x1 | ~x3 | x4 | x5) & (x1 | (x3 ? ~x4 : (x4 | x5)))) : ((x1 | ~x3 | x4) & (~x1 | x3 | ~x4 | x5));
  assign n805 = (x4 | x5 | ~x7 | x0 | x1 | x3) & ((x1 ? (~x5 | ~x7) : (x5 | x7)) | (x0 ? (~x3 | x4) : (x3 | ~x4)));
  assign n806 = (x3 | (x1 ? (~x5 | x7) : (x5 | ~x7)) | (~x0 ^ ~x4)) & (~x4 | ~x5 | ~x7 | x0 | x1 | ~x3);
  assign n807 = ~n810 & (n425 | n808) & (x2 ? n809 : n812);
  assign n808 = x0 ? ((x3 | (x1 ? (x4 | (x2 & x5)) : (~x4 | (~x2 ^ x5)))) & (~x1 | x2 | ~x3 | ~x4 | ~x5)) : ((x4 | (~x2 ^ x5) | (~x1 ^ ~x3)) & (~x3 | ~x4 | (x1 ? (x2 | x5) : ~x2)));
  assign n809 = (x3 | (x0 ? (x4 | (x1 ? (~x5 | ~x6) : x6)) : (~x4 | (x1 ? (~x5 | x6) : (x5 | ~x6))))) & (x0 | ~x1 | ~x3 | ~x6 | (~x4 ^ x5));
  assign n810 = ~n798 & (x0 ? (x4 & ~n811) : ((~x4 & ~n811) | (~x1 & ~x2 & x4)));
  assign n811 = x1 ? (x2 | x5) : (~x2 | ~x5);
  assign n812 = (~x3 | ~x6 | ((~x0 | x1 | x4) & (~x4 | ~x5 | x0 | ~x1))) & (~x0 | x1 | x3 | x6 | (~x4 ^ x5));
  assign z043 = n816 | ~n819 | ~n821 | (x3 ? ~n815 : ~n814);
  assign n814 = (x7 | (x0 ? (x1 ? (x2 ? (x4 | ~x5) : (~x4 | x5)) : (x4 | (~x2 ^ x5))) : ((~x4 | ~x5 | x1 | x2) & (~x1 | (x2 ? (~x4 | ~x5) : x4))))) & (x4 | ~x7 | (x0 ? (~x1 | x2) : (~x5 | (x1 ^ x2))));
  assign n815 = (x5 | ((x2 | ((~x7 | (x0 ? (x1 ^ ~x4) : (x1 | x4))) & (x0 | x1 | ~x4 | x7))) & (x0 | ~x1 | ~x2 | x4 | ~x7))) & (x0 | x1 | ~x2 | ~x4 | ~x7);
  assign n816 = x1 & ((~x7 & ~n817) | (x7 & ~n818 & ~x2 & x4));
  assign n817 = (x4 | (x0 ^ ~x2) | (x3 ? (~x5 | ~x6) : (x5 | x6))) & (~x4 | ~x5 | x6 | ~x0 | x2 | x3);
  assign n818 = (x0 | x6 | (x3 ^ ~x5)) & (~x0 | x3 | ~x5 | ~x6);
  assign n819 = x5 ? ((~x7 | n820) & (~x3 | x7 | n346)) : ((x7 | n820) & (x3 | ~x7 | n346));
  assign n820 = (~x4 | (x0 ^ ~x2) | (~x1 ^ ~x3)) & (~x3 | x4 | (x0 ? (x1 | ~x2) : (~x1 | x2)));
  assign n821 = (n699 | n822) & (x1 | (x0 ? n823 : n824));
  assign n822 = (~x2 | (x5 ? ((~x3 | x6 | x0 | ~x1) & (~x0 | x1 | x3 | ~x6)) : (x0 ? (x1 ? (x3 | x6) : (~x3 | ~x6)) : (x1 ? (x3 | ~x6) : (~x3 | x6))))) & (x0 | x2 | ((x1 | (x3 ? (~x5 | x6) : (x5 | ~x6))) & (~x5 | ~x6 | ~x1 | x3)));
  assign n823 = (x6 | ((~x2 | ((x3 | x4 | ~x5 | x7) & (~x3 | ~x4 | x5 | ~x7))) & (x2 | ~x3 | ~x4 | ~x5 | ~x7))) & (x2 | x5 | ~x6 | (x3 ? (x4 | x7) : (~x4 | ~x7)));
  assign n824 = (~x5 | ~x6 | x7 | ~x2 | x3 | x4) & (x2 | (x3 ? ((~x6 | ~x7 | ~x4 | ~x5) & (x6 | x7 | x4 | x5)) : (x5 | (x4 ? (x6 | ~x7) : (~x6 | x7)))));
  assign z044 = ~n828 | (x3 & (x0 ? ~n827 : ~n826));
  assign n826 = x4 ? (((~x5 ^ x7) | (x1 ? (x2 | ~x6) : (~x2 | x6))) & (~x1 | ~x2 | ~x5 | x6 | ~x7) & (x1 | x2 | x5 | ~x6 | x7)) : ((x5 | (x1 ^ ~x7) | (~x2 ^ ~x6)) & (x1 | x2 | ~x5 | ~x6 | ~x7));
  assign n827 = (x2 | ((x6 | (x1 ? (x4 ? (x5 | x7) : (~x5 | ~x7)) : (x4 | (~x5 ^ x7)))) & (~x4 | ~x5 | ~x6 | (x1 ^ ~x7)))) & (x1 | ~x2 | ((~x4 | ~x5 | x6 | x7) & (x4 | ~x6 | (~x5 ^ x7))));
  assign n828 = (x1 ? n829 : n830) & (x3 | (n831 & n834));
  assign n829 = ((~x3 ^ x6) | ((x0 | ~x2 | x5) & (x2 | ((~x4 | ~x5) & (~x0 | x4 | x5))))) & (~x5 | ((~x3 | ((x0 | (x2 ^ x6)) & (x2 | x4 | ~x6))) & (~x0 | ~x2 | x3 | x4 | x6))) & (x2 | x3 | x5 | x6 | (x0 & ~x4));
  assign n830 = ((x2 ^ x6) | (x3 ? (~x4 | x5) : (~x5 | (~x0 & x4)))) & ((x3 ^ x5) | ((x0 | x2 | ~x4 | ~x6) & (~x2 | x4 | x6))) & (~x3 | x5 | ~x6 | (x4 ? ~x0 : x2)) & (~x4 | ~x5 | x6 | x0 | ~x2 | x3);
  assign n831 = (~n352 | ~n524) & (n832 | n833);
  assign n832 = x0 ? (x1 | ~x5) : (~x1 | x5);
  assign n833 = (x2 | x4 | ~x6 | x7) & (~x2 | ~x4 | x6 | ~x7);
  assign n834 = (n836 | n838) & (n835 | n678) & (n456 | ~n837);
  assign n835 = (~x0 | ~x1 | x2 | x5) & (x0 | x1 | ~x2 | ~x5);
  assign n836 = x2 ? (x6 | x7) : (~x6 | ~x7);
  assign n837 = ~x2 & ~x0 & ~x1;
  assign n838 = (x0 | ~x1 | x4 | ~x5) & (~x0 | x1 | ~x4 | x5);
  assign z045 = n840 | n844 | ~n845 | ~n854 | (x6 & ~n843);
  assign n840 = ~x0 & (x1 ? ~n842 : ~n841);
  assign n841 = x2 ? ((~x3 | ~x4 | ~x5 | x6 | ~x7) & (x3 | x4 | x5 | ~x6 | x7)) : (x4 | ((x6 | x7 | x3 | ~x5) & (~x7 | (x3 ? (x5 ^ x6) : (x5 | ~x6)))));
  assign n842 = (x7 | (x2 ? (~x3 | (x4 ? (x5 | ~x6) : (~x5 | x6))) : (x3 | ~x4 | (x5 ^ x6)))) & (x3 | x5 | ~x7 | (x2 ? (~x4 | x6) : (x4 | ~x6)));
  assign n843 = (~x3 | x4 | ~x5 | x0 | ~x2) & (x3 | ((~x1 | ((~x4 | ~x5 | ~x0 | x2) & (x4 | x5 | x0 | ~x2))) & (x0 | x1 | x2 | (~x4 ^ x5))));
  assign n844 = ~n585 & ((~x0 & x1 & ~x2 & ~x3 & ~x5) | (~x1 & ((x3 & x5 & ~x0 & ~x2) | (x0 & (x2 ? (x3 & ~x5) : (~x3 & x5))))));
  assign n845 = ~n846 & (x0 ? (~n849 & n851) : (~n542 | ~n848));
  assign n846 = ~n847 & ((x0 & ~x2 & x3 & x4 & ~x6) | (~x3 & ((~x0 & x2 & x4 & ~x6) | (x0 & ~x4 & (x2 ^ ~x6)))));
  assign n847 = ~x1 ^ ~x5;
  assign n848 = ~x6 & x5 & x3 & ~x4;
  assign n849 = ~n798 & n850 & x7 & n345;
  assign n850 = ~x4 & x5;
  assign n851 = (n389 | n402) & (n852 | n853);
  assign n852 = x3 ? (~x6 | ~x7) : (x6 | x7);
  assign n853 = (x1 | ~x2 | x4 | x5) & (~x1 | x2 | ~x4 | ~x5);
  assign n854 = x6 ? (x7 ? n855 : n856) : (x7 ? n856 : n855);
  assign n855 = x0 ? ((x1 | ~x3 | ~x5 | (~x2 ^ x4)) & (x3 | x5 | ((x2 | ~x4) & (~x1 | ~x2 | x4)))) : (x2 ? ((~x3 | x4 | x5) & (~x4 | ~x5 | x1 | x3)) : ((~x3 | ~x4 | x5) & (~x1 | (x3 ? ~x4 : (x4 | ~x5)))));
  assign n856 = ((x1 ? (x2 | x4) : (~x2 | ~x4)) | (x0 ? (x3 ^ x5) : (~x3 | x5))) & (x1 | x2 | ((~x4 | ~x5 | x0 | x3) & (x4 | x5 | ~x0 | ~x3))) & (x0 | ~x2 | ~x5 | ((x3 | x4) & (~x1 | ~x3 | ~x4)));
  assign z046 = ~n860 | ~n872 | (~n858 & ~n859);
  assign n858 = ~x0 ^ ~x3;
  assign n859 = (x7 | ((x1 | ~x2 | x4 | x5 | x6) & (x2 | ((~x5 | ~x6 | x1 | x4) & (~x1 | ~x4 | (~x5 ^ x6)))))) & (x1 | ~x2 | x4 | x5 | ~x6 | ~x7);
  assign n860 = ~n862 & ~n863 & ~n867 & (n368 | n861) & n869;
  assign n861 = ((x1 ? (x3 | x5) : (~x3 | ~x5)) | (x2 ? (~x4 | x7) : (x4 | ~x7))) & (x2 | ((~x1 | x3 | ~x4 | ~x5 | ~x7) & (x1 | ~x3 | x4 | x5 | x7)));
  assign n862 = ~n440 & ((x3 & ((~x0 & x1 & x2 & x4) | (x0 & (x1 ? (~x2 & ~x4) : x4)))) | (~x0 & ~x3 & (~x1 ^ ~x4)));
  assign n863 = ~n443 & (n866 | (~n864 & n865));
  assign n864 = x1 ^ ~x2;
  assign n865 = x0 & ~x3;
  assign n866 = x3 & x2 & ~x0 & ~x1;
  assign n867 = ~n868 & ((n542 & n369) | (n354 & n370));
  assign n868 = (x0 | ~x3 | x5 | x6) & (~x0 | x3 | ~x5 | ~x6);
  assign n869 = (n551 | n871) & (~n870 | ~n283 | ~n361);
  assign n870 = ~x5 & x7;
  assign n871 = (~x3 | x4 | x5 | ~x7) & (x3 | ~x4 | ~x5 | x7);
  assign n872 = ~n873 & ~n874 & ~n875 & ~n876 & (n878 | ~n879);
  assign n873 = n384 & (x0 ? ((~x5 & ~x7 & ~x2 & ~x3) | (x2 & x3 & x5 & x7)) : ((x5 & x7 & x2 & ~x3) | (~x2 & (x3 ? (x5 & ~x7) : (~x5 & x7)))));
  assign n874 = ~n665 & ((x0 & x1 & x2 & ~x3 & ~x4) | (~x0 & ~x2 & x3 & (~x1 ^ ~x4)));
  assign n875 = ~n443 & ((x2 & n349 & (~x3 ^ x6)) | (~x2 & ~x3 & ~x6 & n321));
  assign n876 = ~n877 & (x3 ? (x7 & n542) : (~x7 & n354));
  assign n877 = (x0 | ~x4 | ~x5 | x6) & (~x0 | ~x6 | (x4 ^ x5));
  assign n878 = (~x0 | x2 | x3 | x4 | ~x6) & (x0 | x6 | (x2 ? (~x3 | ~x4) : (x3 | x4)));
  assign n879 = x7 & ~x1 & x5;
  assign z047 = ~n886 | (x2 ? ~n883 : (x0 ? ~n881 : ~n882));
  assign n881 = x4 ? ((x1 | x7 | ((x5 | x6) & (~x3 | ~x5 | ~x6))) & (x5 | x6 | ~x7 | ~x1 | ~x3)) : ((x1 | x3 | x5 | ~x6 | x7) & (~x1 | ((x5 | ~x6 | ~x7) & (x6 | x7 | x3 | ~x5))));
  assign n882 = (x5 | ((~x7 | ((x1 | x3 | x4 | x6) & (~x1 | ((x3 | x4 | ~x6) & (~x4 | x6))))) & (x1 | x3 | ~x4 | x6 | x7))) & (~x4 | ~x5 | ~x6 | (x1 ? (~x3 | ~x7) : x7));
  assign n883 = (x0 | n884) & (~x0 | x1 | ~x5 | n885);
  assign n884 = (~x3 | ((~x4 | ((~x1 | (x5 ? (x6 | x7) : (~x6 | ~x7))) & (~x6 | x7 | x1 | x5))) & (x1 | x4 | x5 | ~x6 | ~x7))) & (x4 | ~x5 | (x1 ? ((x6 | ~x7) & (x3 | ~x6 | x7)) : (x6 | x7)));
  assign n885 = (~x3 | x4 | x6 | x7) & (~x4 | ((x6 | ~x7) & (x3 | ~x6 | x7)));
  assign n886 = ~n887 & n890 & (x4 ? (x2 | n889) : n888);
  assign n887 = ~n416 & ((x0 & ~x2 & ~x3 & (x1 ^ ~x4)) | (x2 & ((~x1 & x3 & x4) | (~x0 & (x1 ? (x3 & ~x4) : x4)))));
  assign n888 = (x0 | x1 | x2 | x5 | ~x6) & (((x2 | ~x3) & (~x0 | ~x2 | x3)) | (x1 ? (~x5 | x6) : (x5 | ~x6)));
  assign n889 = x1 ? (~x6 | (x0 ? ~x3 : x5)) : (x6 | ((~x3 | ~x5) & (x0 | (~x3 & ~x5))));
  assign n890 = (n750 | n892) & (n891 | n893);
  assign n891 = x1 ^ ~x7;
  assign n892 = (x1 | ((x4 | ~x6 | x0 | x3) & (~x0 | (x3 ? (x4 | ~x6) : (~x4 | x6))))) & (x0 | ~x1 | x3 | (x4 ^ x6));
  assign n893 = x5 ? ((x0 | ((x4 | ~x6 | x2 | ~x3) & (~x4 | x6 | ~x2 | x3))) & (~x0 | ~x2 | x3 | x4 | ~x6)) : ((x4 | x6 | x2 | ~x3) & (~x0 | x3 | (x2 ? (x4 | x6) : (~x4 | ~x6))));
  assign z048 = n895 | n900 | (~n425 & ~n899) | (~n437 & ~n898);
  assign n895 = ~x0 & (x1 ? ~n896 : ~n897);
  assign n896 = (~x4 | ((x2 | ~x3 | ~x5 | x6 | ~x7) & (~x2 | x3 | x5 | x7))) & (x5 | ((~x6 | x7 | ~x2 | x4) & (x2 | x3 | x6 | ~x7))) & (x3 | ~x5 | (x2 ? (~x7 | (x4 & x6)) : (x7 | (x4 & ~x6))));
  assign n897 = x3 ? ((~x4 | ((~x6 | x7 | x2 | x5) & (~x2 | (x5 ? (~x6 | x7) : (x6 | ~x7))))) & (x6 | ~x7 | x2 | ~x5)) : (x2 ? (x5 ? (x6 | ~x7) : (x7 | (x4 & ~x6))) : ((x5 | x6 | ~x7) & (~x6 | x7 | x4 | ~x5)));
  assign n898 = (~x3 | (~x2 ^ ~x5) | (x0 ^ (~x1 & x4))) & (~x0 | x3 | x4 | ((~x2 | x5) & (~x1 | x2 | ~x5)));
  assign n899 = x2 ? ((x4 | ~x5 | ~x0 | x3) & (x5 | ((x1 | ~x3 | ~x4) & (x0 | (~x3 & (x1 | ~x4)))))) : ((x3 | x5 | ((~x1 | x4) & (~x0 | (~x1 & x4)))) & (~x5 | (((x1 & ~x4) | (x0 & ~x3)) & (x0 | ~x3))));
  assign n900 = x0 & ((n354 & ~n902) | (~x2 & ~n901));
  assign n901 = ((~x6 ^ x7) & (x1 ^ ~x4)) | (x1 & ~x3 & ~x4) | (~x1 & x3 & x4) | (x5 & x7) | (~x5 & ~x7);
  assign n902 = x4 ? ((x3 | ~x5 | ~x7) & (x5 | ~x6 | x7)) : ((~x5 | x6 | ~x7) & (~x3 | x5 | x7));
  assign z049 = ~n910 | (x3 ? ~n904 : (x5 ? ~n909 : ~n908));
  assign n904 = (x0 | n907) & (n437 | n906) & (n559 | n905);
  assign n905 = (~x4 | ((~x0 | x1 | x6 | ~x7) & (x0 | ((~x6 | ~x7) & (x1 | x6 | x7))))) & (x0 | ~x1 | x4 | x6 | ~x7);
  assign n906 = (~x1 | ((~x0 | x2 | ~x4) & (x4 | x5 | x0 | ~x2))) & (~x0 | x1 | ((~x2 | ~x4 | x5) & (x4 | (x2 & ~x5))));
  assign n907 = (x1 | (x2 ? (~x4 | x5 | (x6 ^ x7)) : (~x5 | ((x6 | x7) & (x4 | ~x6 | ~x7))))) & (x2 | ~x4 | ~x5 | ((x6 | x7) & (~x1 | ~x6 | ~x7)));
  assign n908 = x7 ? ((~x4 | ((~x0 | ~x1 | x2 | ~x6) & (x0 | x6 | (x1 & x2)))) & (~x0 | x1 | x4 | ~x6) & (~x2 | ((x0 | ~x1 | x4 | ~x6) & (~x0 | (x1 ? (x4 | x6) : ~x6))))) : ((x6 | ((~x1 | (~x0 ^ ~x4)) & (~x0 | ((~x2 | ~x4) & (x1 | x2 | x4))))) & (x0 | ~x6 | ((x2 | ~x4) & (x1 | (x2 & ~x4)))));
  assign n909 = x0 ? (x1 ? (x2 | ((~x6 | ~x7) & (~x4 | x6 | x7))) : (x4 | (x6 ^ x7))) : ((~x4 | (~x1 & ~x2) | (~x6 ^ x7)) & (x1 | x4 | ((~x6 | x7) & (x2 | x6 | ~x7))));
  assign n910 = n911 & (x1 ? n913 : n912);
  assign n911 = x1 ? ((~x3 | ~x4 | x6 | x0 | ~x2) & (x2 | x4 | (x0 ? (x3 ^ x6) : (x3 | ~x6)))) : ((~x0 | x2 | x3 | ~x4 | ~x6) & (~x3 | x4 | x6 | x0 | ~x2));
  assign n912 = ((~x0 ^ ~x3) | ((~x5 | x6 | x2 | ~x4) & (x5 | ~x6 | ~x2 | x4))) & ((x0 ? (~x2 | x3) : (x2 | ~x3)) | (x4 ? (~x5 | ~x6) : (x5 | x6)));
  assign n913 = (x4 | ~x5 | x6 | ~x0 | ~x2 | x3) & (x0 | (~x4 ^ x5) | (x2 ? (x3 | ~x6) : (~x3 | x6)));
  assign z050 = (x3 & (n916 | n917)) | ~n918 | (~x4 & ~n915);
  assign n915 = x1 ? ((x3 | x5 | ~x7 | ~x0 | x2) & (x0 | ((~x5 | ~x7 | x2 | ~x3) & (~x2 | ((x5 | x7) & (x3 | ~x5 | ~x7)))))) : (((~x0 ^ ~x2) | ((~x5 | x7) & (~x3 | x5 | ~x7))) & (~x5 | x7 | x2 | ~x3) & (x3 | x5 | ~x7 | x0 | ~x2));
  assign n916 = ~n589 & ((x2 & x5 & x7 & n349) | (~x2 & ~x5 & (x7 ? n349 : n321)));
  assign n917 = n372 & ((x0 & ~x1 & x2 & x4 & x5) | (~x0 & ((x4 & x5 & ~x1 & ~x2) | (x1 & ~x4 & (~x2 ^ x5)))));
  assign n918 = ~n923 & n924 & (x3 | (n919 & n922));
  assign n919 = (~x1 | x7 | n921) & (n920 | (x4 ? (~x6 | ~x7) : (~x6 ^ x7)));
  assign n920 = x0 ? (x1 ? (x2 | ~x5) : (~x2 | x5)) : (x1 | (x2 ^ x5));
  assign n921 = (~x2 | ((~x5 | ~x6 | x0 | ~x4) & (x5 | x6 | ~x0 | x4))) & (x0 | x2 | x5 | (x4 ^ x6));
  assign n922 = (~x0 | x1 | x2 | ~x4 | ~x7) & (x4 | ((x0 | ~x1 | x2 | ~x7) & (~x0 | (x1 ? (~x2 | ~x7) : (x2 | x7)))));
  assign n923 = x4 & ((~x1 & (~x5 ^ x7) & (x0 ^ ~x2)) | (~x0 & x1 & (x2 ? (~x5 & x7) : (x5 & ~x7))));
  assign n924 = (~x0 | x1 | x2 | ~x3 | ~x4 | ~x7) & ((x0 ? (~x1 | x2) : (x1 | ~x2)) | ((~x4 | x7) & (~x3 | x4 | ~x7)));
  assign z051 = n930 | n931 | ~n932 | (x1 & ~n926);
  assign n926 = ~n927 & ~n928 & ((x0 & ~n294) | n736 | (~x0 & ~n335));
  assign n927 = ~n520 & ((~x0 & x5 & (x2 ? (x4 & ~x7) : (~x4 & x7))) | (x0 & ~x2 & ~x4 & ~x5 & x7));
  assign n928 = ~x4 & n929 & (x0 ? n531 : (~x5 & n372));
  assign n929 = x2 & ~x3;
  assign n930 = x5 & ((~x2 & ((x1 & (x0 ? ~x6 : (~x3 & x6))) | (x0 & (x6 ? (~x1 | x3) : ~x3)))) | (~x0 & x2 & ((x3 & ~x6) | (~x1 & (x3 | ~x6)))));
  assign n931 = n312 & (((~x2 ^ x7) & (x0 ? (~x1 & x3) : (x1 & ~x3))) | (x0 & x1 & x2 & ~x3 & ~x7) | (~x0 & ~x1 & ~x2 & x7));
  assign n932 = ~n933 & (x1 | (~n935 & ~n937 & (x4 | n934)));
  assign n933 = ~x5 & (x6 ? (x0 ? (x1 ? (~x2 & ~x3) : (x2 & x3)) : ((~x1 & ~x2 & x3) | (x2 & (x1 | ~x3)))) : ((~x0 & x1 & ~x2 & x3) | (x0 & ~x1 & x2 & ~x3)));
  assign n934 = ((~x0 ^ ~x2) | ((x6 | x7 | ~x3 | x5) & (~x6 | ~x7 | x3 | ~x5))) & (x0 | ~x2 | x5 | ~x7 | (x3 ^ x6));
  assign n935 = ~n529 & ((n278 & n369) | (x0 & ~n936));
  assign n936 = x2 ? (~x4 | x7) : (x4 | ~x7);
  assign n937 = n544 & n369 & (x2 ? n531 : n312);
  assign z052 = n942 | ~n943 | (~x6 & (~n940 | (~x2 & ~n939)));
  assign n939 = (x4 | x5 | ~x7 | x0 | x1 | x3) & (~x3 | ((~x0 | ((x5 | x7 | x1 | ~x4) & (~x5 | ~x7 | ~x1 | x4))) & (x0 | ~x1 | ~x4 | ~x5 | ~x7)));
  assign n940 = (x1 | ~x5 | ~x7 | n941) & (x5 | x7 | ((~n686 | ~n288) & (~x1 | n941)));
  assign n941 = (x0 | ~x2 | ~x3 | x4) & (x3 | (x0 ? (~x2 ^ ~x4) : (x2 | ~x4)));
  assign n942 = n531 & (x1 ? ((x3 & x4 & x0 & ~x2) | (~x3 & ~x4 & ~x0 & x2)) : (x0 ? (x2 ? (x3 & ~x4) : (~x3 & x4)) : (x3 & (~x2 ^ x4))));
  assign n943 = n947 & n949 & (n437 | (n945 & (n944 | n946)));
  assign n944 = x0 ? (~x1 | x2) : (x1 | ~x2);
  assign n945 = (~x0 | x1 | x2 | x3 | x4 | x5) & (x0 | ~x1 | ~x2 | ~x3 | ~x4 | ~x5);
  assign n946 = x3 ? (x4 | x5) : (~x4 | ~x5);
  assign n947 = (x1 | ((~x0 | ((x6 | n948) & (~x2 | ~x6 | n946))) & (x0 | x2 | ~x6 | n946))) & (x0 | ~x1 | ((~x6 | n948) & (x2 | x6 | n946)));
  assign n948 = (~x2 | x3 | x4 | x5) & (~x4 | ~x5 | x2 | ~x3);
  assign n949 = (~x6 | (x7 ? n952 : (n950 | n951))) & (n950 | n953) & (x6 | (x7 ? (n950 | n951) : n952));
  assign n950 = x4 ^ ~x5;
  assign n951 = (~x0 | x1 | ~x2 | x3) & (x0 | x2 | (~x1 ^ ~x3));
  assign n952 = ((x2 ^ x4) | (x0 ? (x1 | ~x3) : (~x1 | x3))) & (~x0 | ~x1 | ~x2 | x3 | x4) & (x0 | x1 | x2 | ~x3 | ~x4);
  assign n953 = (x0 | ~x1 | ~x2 | ~x3 | x6) & (~x0 | x1 | x2 | x3 | ~x6) & ((x3 ^ x6) | (x0 ? (~x1 | x2) : (x1 | ~x2)));
  assign z053 = ~n957 | (~x2 & ~n955) | (~n425 & ~n956);
  assign n955 = x0 ? (x1 ? ((x5 | x7 | ~x3 | x4) & (x3 | (x4 ? (~x5 ^ x7) : (~x5 | ~x7)))) : ((~x5 | ~x7 | ~x3 | ~x4) & (x5 | x7 | x3 | x4))) : ((~x1 | x3 | ~x4 | ~x5 | ~x7) & ((x1 ^ x3) | (x4 ? (x5 | x7) : (~x5 ^ x7))));
  assign n956 = ((x1 ^ ~x5) | ((x3 | x4 | ~x0 | x2) & (x0 | (x2 ? (~x3 | x4) : (x3 | ~x4))))) & (x0 | ((x1 | ~x2 | x3 | x4 | x5) & (~x1 | x2 | ~x3 | ~x4 | ~x5))) & (~x0 | ((x1 | ~x4 | (x2 ? (x3 | ~x5) : (~x3 | x5))) & (~x3 | x4 | ~x5 | ~x1 | x2)));
  assign n957 = ~n959 & ~n961 & (~n958 | ~n339) & (~x2 | n960);
  assign n958 = ~x3 & x2 & x0 & x1;
  assign n959 = x0 & (x1 ? ((~x4 & ~x7 & x2 & ~x3) | (x4 & x7 & ~x2 & x3)) : ((x4 & x7 & ~x2 & ~x3) | (x3 & (x2 ? (x4 ^ x7) : (~x4 & ~x7)))));
  assign n960 = ((~x5 ^ x7) | ((~x0 | x1 | x3 | x4) & (x0 | ~x4 | (x1 ^ x3)))) & (~x4 | x5 | x7 | ~x0 | x1 | x3) & (x0 | x4 | ((~x1 | ~x3 | ~x5 | ~x7) & (x1 | (x3 ? (x5 | x7) : (~x5 | ~x7)))));
  assign n961 = ~x0 & (((x4 ^ x7) & (x1 ? (x2 & ~x3) : (~x2 & x3))) | (~x1 & x2 & x3 & x4 & x7) | (x1 & ~x2 & ~x3 & ~x4 & ~x7));
  assign z054 = ~n967 | ~n970 | (x6 ? ~n956 : ~n963);
  assign n963 = (~x3 | n966) & (x3 | n964) & (n307 | n965);
  assign n964 = x2 ? ((x7 | ((~x4 | ~x5 | x0 | ~x1) & (~x0 | (x1 ? (x4 | ~x5) : (~x4 | x5))))) & (x0 | x4 | ~x7 | (x1 ^ ~x5))) : ((~x0 | ~x1 | x4 | ~x5 | ~x7) & (x0 | x1 | ~x4 | x5 | x7));
  assign n965 = x0 ? (x2 | (x1 ? (~x3 | x5) : (x3 ^ x5))) : ((x3 | ~x5 | ~x1 | x2) & (~x3 | x5 | x1 | ~x2));
  assign n966 = (x1 | (x4 ? (~x5 | x7) : (x5 | ~x7)) | (~x0 ^ ~x2)) & (x0 | ~x1 | ((x5 | x7 | x2 | ~x4) & (~x5 | ~x7 | ~x2 | x4)));
  assign n967 = n969 & (n968 | (x2 ? (x4 | x5) : (~x4 | ~x5)));
  assign n968 = (~x1 | x3 | x7) & (~x0 | (x1 ? x3 : (~x3 | x7)));
  assign n969 = (x1 | ((~x0 | x2 | ~x3 | x4 | x5) & (x0 | ~x2 | x3 | ~x4 | ~x5))) & (x0 | ~x1 | (x3 ^ x5) | (x2 ^ x4));
  assign n970 = (x7 | n971) & (n683 | ((~x0 | (x1 ? (x2 | x7) : ~x2)) & (x1 | (x2 ? x7 : x0))));
  assign n971 = (x0 | ~x3 | x4 | (x1 ? (~x2 | ~x5) : (x2 | x5))) & (x3 | ~x4 | x5 | ~x0 | x1 | x2);
  assign z055 = n973 | ~n976 | ~n983 | (x0 & ~n975);
  assign n973 = ~n974 & (x1 ? ((x3 & x4 & x0 & ~x2) | (~x3 & ~x4 & ~x0 & x2)) : (x0 ? (x2 ? (x3 & ~x4) : (~x3 & x4)) : (x3 & (~x2 ^ x4))));
  assign n974 = x5 ? (x6 | x7) : (~x6 | ~x7);
  assign n975 = ((x2 ^ ~x6) | ((x4 | x5 | ~x1 | x3) & (x1 | (x3 ? (~x4 | x5) : (x4 | ~x5))))) & (x1 | ((x2 | ~x3 | x4 | x5 | x6) & (~x2 | x3 | ~x4 | ~x5 | ~x6)));
  assign n976 = ~n979 & ~n982 & (n977 | n978) & (~n321 | n981);
  assign n977 = (x0 | ~x2 | (~x1 ^ ~x3)) & (~x0 | ~x1 | x2 | x3);
  assign n978 = (~x4 | x5 | x6 | x7) & (~x6 | ~x7 | x4 | ~x5);
  assign n979 = ~n980 & ((~x0 & x2 & (~x1 ^ ~x5)) | (x0 & x1 & ~x2 & x5));
  assign n980 = x3 ? (x4 | ~x6) : (~x4 | x6);
  assign n981 = (~x2 | x3 | x4 | x5 | x6 | x7) & (x2 | ~x3 | ~x4 | ~x5 | ~x6 | ~x7);
  assign n982 = n444 & ((n313 & n611) | (n373 & n612));
  assign n983 = (n437 | n984) & (x0 | n985);
  assign n984 = ((~x0 ^ x4) | (x1 ? (x2 ? (x3 | ~x5) : (~x3 | x5)) : (x2 | (x3 ^ x5)))) & (x1 | ~x2 | ((~x0 | ~x4 | (x3 ^ x5)) & (x4 | x5 | x0 | ~x3))) & (x3 | x4 | ~x5 | x0 | ~x1 | x2);
  assign n985 = x2 ? ((x4 | x5 | ~x6 | x1 | x3) & (~x4 | ~x5 | x6 | ~x1 | ~x3)) : ((~x4 | x5 | x6 | x1 | ~x3) & ((x4 ^ x6) | (x1 ? (x3 ^ x5) : (x3 | ~x5))));
  assign z056 = ~n990 | ~n994 | (~n425 & ~n988) | (~n987 & ~n989);
  assign n987 = x0 ? (x1 | ~x3) : (~x1 | x3);
  assign n988 = ((x3 ? (~x4 | x5) : (x4 | ~x5)) | (x0 ? (~x1 | x2) : (x1 | ~x2))) & ((x3 ^ x5) | ((~x0 | x1 | x2 | ~x4) & (x0 | ~x1 | ~x2 | x4))) & (x0 | x2 | ((x4 | x5 | x1 | ~x3) & (~x4 | ~x5 | ~x1 | x3))) & (~x3 | x4 | x5 | ~x0 | x1 | ~x2);
  assign n989 = (x2 | ~x4 | x5 | ~x6 | x7) & (~x2 | x4 | ~x5 | x6 | ~x7);
  assign n990 = n991 & (n944 | n871) & (~n509 | ~n783 | ~n786);
  assign n991 = (~n460 | ~n993) & (~n664 | ~n361 | ~n992);
  assign n992 = x2 & ~x0 & x1;
  assign n993 = x7 & ~x5 & ~x3 & ~x4;
  assign n994 = n995 & ~n997 & (n951 | (~n269 & ~n996));
  assign n995 = (n443 | n951) & (n440 | n952);
  assign n996 = ~x7 & x6 & x4 & x5;
  assign n997 = ~n389 & ((~x0 & x1 & x2 & x3 & ~x5) | (x0 & ~x1 & ~x2 & ~x3 & x5) | ((~x3 ^ x5) & (x0 ? (x1 & ~x2) : (~x1 & x2))));
  assign z057 = n999 | n1002 | ~n1007 | (~x2 & ~n1006);
  assign n999 = x3 & (x2 ? ~n1001 : ~n1000);
  assign n1000 = x0 ? (x1 ? ((~x6 | ~x7 | x4 | x5) & (x7 | (x4 ? (x5 ^ x6) : (~x5 | x6)))) : ((x6 | ~x7 | ~x4 | ~x5) & (~x6 | x7 | x4 | x5))) : ((~x1 | ~x4 | ~x5 | x6 | x7) & ((x1 ^ x7) | (x4 ? (x5 | ~x6) : (x5 ^ x6))));
  assign n1001 = ((x5 ^ x6) | ((x0 | ~x4 | (x1 ^ x7)) & (~x0 | x1 | x4 | x7))) & (x0 | x4 | ((x1 | (x5 ? (x6 | x7) : (~x6 | ~x7))) & (x6 | ~x7 | ~x1 | ~x5))) & (x5 | ~x6 | x7 | ~x0 | x1 | ~x4);
  assign n1002 = ~x3 & ((~x0 & ~n1003) | (~n585 & ~n1004) | (x0 & ~n1005));
  assign n1003 = x2 ? ((x5 | x6 | ~x7 | x1 | ~x4) & (~x5 | ~x6 | x7 | ~x1 | x4)) : (x1 ? ((x6 | ~x7 | ~x4 | ~x5) & (~x6 | x7 | x4 | x5)) : (~x5 | (x4 ? (x6 | x7) : (~x6 | ~x7))));
  assign n1004 = x1 ? ((~x5 | ~x7 | ~x0 | x2) & (x5 | x7 | x0 | ~x2)) : (x0 ? (x2 ? (x5 | ~x7) : (~x5 | x7)) : (~x7 | (x2 ^ x5)));
  assign n1005 = x1 ? (x5 | ((x6 | ~x7 | x2 | ~x4) & (~x2 | x7 | (~x4 ^ x6)))) : ((~x2 ^ ~x5) | (x4 ? (x6 | x7) : (~x6 | ~x7)));
  assign n1006 = (x4 | ~x6 | x7 | x0 | ~x1 | ~x3) & (~x7 | ((x0 | ~x1 | x3 | x4 | ~x6) & (x1 | ((~x4 | ~x6 | x0 | ~x3) & (~x0 | (x3 ? (x4 | ~x6) : (~x4 | x6)))))));
  assign n1007 = (n1010 | n1011) & (~n487 | n1008) & (n661 | n1009);
  assign n1008 = (~x1 | ((x3 | x4 | x6 | ~x7) & (~x3 | x7 | (x4 ^ x6)))) & (x1 | x3 | x4 | x6 | x7);
  assign n1009 = x3 ? (x6 | ~x7) : (~x6 | x7);
  assign n1010 = x2 ? (~x6 | ~x7) : (x6 | x7);
  assign n1011 = (x0 | ~x1 | x3 | ~x4) & (~x0 | (x1 ? (x3 | x4) : (~x3 | ~x4)));
  assign z058 = ~n1014 | (~n425 & ~n956) | (~n665 & ~n1013);
  assign n1013 = x0 ? (x1 ? ((~x4 | x6 | x2 | ~x3) & (x4 | ~x6 | ~x2 | x3)) : ((~x4 | x6 | x2 | x3) & (~x3 | (x2 ? (x4 ^ x6) : (x4 | ~x6))))) : ((x3 | x4 | ~x6 | ~x1 | x2) & (~x3 | ~x4 | x6 | x1 | ~x2) & ((x4 ^ x6) | (x1 ? (~x2 | x3) : (x2 | ~x3))));
  assign n1014 = ~n1017 & n1019 & n1022 & (n1015 | n1016);
  assign n1015 = ~x4 ^ ~x5;
  assign n1016 = x0 ? (x2 | ((x1 | (x3 ? (x6 | ~x7) : (~x6 | x7))) & (~x6 | x7 | ~x1 | ~x3))) : ((x3 | x6 | ~x7 | ~x1 | x2) & (~x3 | ~x6 | x7 | x1 | ~x2));
  assign n1017 = ~x0 & ((n268 & n1018) | (~n989 & (n273 | n367)));
  assign n1018 = ~x7 & x6 & ~x4 & ~x5;
  assign n1019 = (n1020 | n1021) & (~n288 | ~n317 | ~n615);
  assign n1020 = (~x4 | x5 | x6 | ~x7) & (x4 | ~x5 | ~x6 | x7);
  assign n1021 = (~x0 | x1 | ~x2 | ~x3) & (x0 | (x1 ? (~x2 | x3) : (x2 | ~x3)));
  assign n1022 = (n440 | n1023) & (~n865 | n1024);
  assign n1023 = (x3 | ((x0 | x1 | ~x2 | ~x4) & (~x0 | (x1 ? (x2 | ~x4) : (~x2 | x4))))) & (x0 | ~x1 | ~x3 | (x2 ^ x4));
  assign n1024 = (~x5 | x6 | ~x7 | ~x1 | x2 | x4) & (~x2 | x5 | ((~x6 | x7 | x1 | ~x4) & (~x1 | x6 | (~x4 ^ x7))));
  assign z059 = ~n1036 | n1035 | n1033 | n1031 | n1026 | n1028;
  assign n1026 = ~x1 & (x0 ? ~n981 : ~n1027);
  assign n1027 = x3 ? ((x2 | ((~x6 | ~x7 | ~x4 | ~x5) & (x5 | x6 | x7))) & (x5 | ((~x4 | x6 | x7) & (~x6 | ~x7 | (~x2 & x4))))) : ((~x5 | ((x4 | x6 | x7) & (~x2 | ((x6 | x7) & (x4 | ~x6 | ~x7))))) & (x2 | x5 | ~x7 | (x4 ^ x6)));
  assign n1028 = x1 & ((~x0 & ~n1030) | (~n978 & (n342 | n1029)));
  assign n1029 = ~x3 & x0 & ~x2;
  assign n1030 = (x2 | (x3 ? ((x6 | x7 | x4 | ~x5) & (~x6 | ~x7 | ~x4 | x5)) : (~x5 | ((~x6 | ~x7) & (~x4 | x6 | x7))))) & (x3 | x4 | x5 | x6 | x7);
  assign n1031 = ~n437 & ~n1032;
  assign n1032 = ((x2 ? (x3 | ~x5) : (~x3 | x5)) | (x0 ? (~x1 | x4) : ~x4)) & (x1 | ~x2 | ((~x0 | ~x4 | (x3 ^ x5)) & (x4 | x5 | x0 | ~x3))) & (x2 | ((x4 | (x0 ? (x1 | (x3 ^ x5)) : ((x3 | ~x5) & (~x1 | (x3 & ~x5))))) & (x0 | x1 | ~x4 | (~x3 & x5))));
  assign n1033 = ~x0 & ~n1034;
  assign n1034 = (x2 | (x3 ? (x4 | x6) : (~x4 | ~x6)) | (~x1 ^ x5)) & (x1 | ~x2 | ((x5 | x6 | x3 | ~x4) & (~x3 | ~x5 | (~x4 ^ x6))));
  assign n1035 = ~n974 & ((x1 & ((x3 & x4 & x0 & ~x2) | (~x3 & ~x4 & ~x0 & x2))) | (x0 & ~x1 & (x2 ? (x3 & ~x4) : (~x3 & x4))));
  assign n1036 = ~n1037 & ~n1040 & (n1039 | (x0 ? (x2 | ~x5) : (~x2 | x5)));
  assign n1037 = n321 & ((~x2 & x3 & n1038) | (x2 & ~x3 & x5 & ~n585));
  assign n1038 = ~x6 & ~x4 & ~x5;
  assign n1039 = (~x1 | (x3 ? (x4 | ~x6) : (~x4 | x6))) & (x1 | x3 | x4 | ~x6);
  assign n1040 = ~n1042 & ((x3 & n654 & n349) | (n1041 & ~n315));
  assign n1041 = x0 & ~x5;
  assign n1042 = x2 ^ ~x6;
  assign z060 = ~n1046 | ~n1053 | (~x3 & (x2 | ~n1044) & (~x2 | ~n1045));
  assign n1044 = (x5 | ((x0 | x1 | x4 | ~x6 | x7) & (~x0 | ((x6 | x7 | x1 | ~x4) & (~x1 | (x4 ? (x6 | ~x7) : (~x6 | x7))))))) & (x0 | ~x5 | ((x6 | ~x7 | ~x1 | x4) & (x1 | (x4 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n1045 = (x4 | (~x6 ^ x7) | (x0 ? (x1 | x5) : (~x1 | ~x5))) & (x5 | ~x6 | ~x7 | x0 | ~x1 | ~x4);
  assign n1046 = (x2 ? n1052 : n1051) & (~x3 | (~n1047 & ~n1049));
  assign n1047 = ~x4 & ((n992 & n1048) | (~x5 & n374 & n460));
  assign n1048 = ~x7 & x5 & ~x6;
  assign n1049 = n1050 & ((x5 & ((~x1 & ((x6 & ~x7) | (~x2 & ~x6 & x7))) | (x6 & x7 & x1 & x2))) | (x1 & x2 & ~x5 & (x6 ^ x7)));
  assign n1050 = ~x0 & x4;
  assign n1051 = x0 ? (x1 ? ((~x5 | x7 | x3 | ~x4) & (x5 | ~x7 | ~x3 | x4)) : (x3 | ((x5 | ~x7) & (x4 | ~x5 | x7)))) : ((~x1 | ~x3 | ~x4 | ~x5 | x7) & (x1 | (x3 ? ((x5 | ~x7) & (x4 | ~x5 | x7)) : (~x5 | (~x4 ^ x7)))));
  assign n1052 = (x1 | (x0 ^ ~x3) | (x4 ? (x5 | ~x7) : (~x5 | x7))) & (x0 | ~x1 | ((x5 | ~x7 | x3 | x4) & (~x5 | x7 | ~x3 | ~x4)));
  assign n1053 = (n1054 | n1057) & (n440 | n1056) & (n425 | n1055);
  assign n1054 = ~x0 ^ ~x5;
  assign n1055 = (x3 | ~x4 | ~x5 | x0 | x1 | ~x2) & (~x3 | ((~x0 | x5 | (x1 ? (x2 | ~x4) : (~x2 | x4))) & (x2 | x4 | ~x5 | x0 | ~x1)));
  assign n1056 = (~x4 | (x0 ? (x1 | ~x3) : (~x1 | x3))) & (~x0 | ((~x1 | ~x2 | x3 | x4) & (x1 | x2 | ~x3))) & (x0 | ~x2 | x4 | (~x1 ^ ~x3));
  assign n1057 = (x2 | (((~x3 ^ x7) | (x1 ? (x4 | ~x6) : (~x4 | x6))) & (~x1 | x6 | (x3 ? (~x4 | ~x7) : (x4 | x7))))) & (x1 | ((~x6 | x7 | x3 | ~x4) & (~x2 | ~x3 | x4 | x6 | ~x7)));
  assign z061 = n1069 | ~n1072 | (x1 ? ~n1062 : (~n1059 | ~n1068));
  assign n1059 = x0 ? n1060 : n1061;
  assign n1060 = x2 ? ((~x6 | x7 | x4 | ~x5) & (~x3 | ~x4 | x5 | x6 | ~x7) & (x3 | ((x4 | ~x5 | ~x6) & (x7 | (x4 ? (~x5 ^ x6) : (x5 | x6)))))) : ((x3 | ((x6 | ~x7 | ~x4 | ~x5) & (~x6 | x7 | x4 | x5))) & (x6 | ~x7 | x4 | x5) & (~x3 | ((~x6 | ~x7 | x4 | ~x5) & (~x4 | (x5 ? (x6 | x7) : (~x6 | ~x7))))));
  assign n1061 = x2 ? ((~x3 | x4 | ~x5 | ~x6 | ~x7) & ((x3 ^ ~x7) | (x4 ? (~x5 ^ x6) : (x5 | x6)))) : (x3 ? ((x6 | ~x7 | ~x4 | ~x5) & (~x6 | x7 | x4 | x5)) : ((~x6 | ~x7 | x4 | x5) & (x7 | (x4 ? (x5 ^ x6) : (~x5 | x6)))));
  assign n1062 = ~n1063 & ~n1064 & ~n1065 & (~n850 | ~n544 | ~n1067);
  assign n1063 = ~n585 & ((~x2 & ((~x5 & ~x7 & ~x0 & ~x3) | (x0 & x5 & (x3 ^ x7)))) | (~x0 & x2 & ~x3 & x5 & x7));
  assign n1064 = ~n382 & (x0 ? (~x3 & ~x5 & (x4 ^ x6)) : (x3 & x5 & (~x4 ^ x6)));
  assign n1065 = ~x5 & ~n1066;
  assign n1066 = ((x0 ? (x2 | ~x3) : (~x2 | x3)) | (x4 ? (x6 | x7) : (~x6 | ~x7))) & (x0 | ~x3 | ((x6 | ~x7 | x2 | ~x4) & (~x6 | x7 | ~x2 | x4)));
  assign n1067 = ~x7 & (~x2 ^ ~x6);
  assign n1068 = (~x2 | ((~x0 | ~x3 | (x4 ? ~x6 : (x6 | ~x7))) & (x0 | x3 | ~x4 | x6 | x7))) & (x0 | x2 | ~x7 | (x3 ? (x4 | ~x6) : (~x4 | x6)));
  assign n1069 = ~n406 & ((x2 & n1070 & n783) | (~n1042 & ~n1071));
  assign n1070 = ~x4 & x6;
  assign n1071 = x0 ? (x1 | x4) : (~x1 | ~x4);
  assign n1072 = n1073 & (n1009 | ((x0 | ~x2 | (~x1 ^ ~x4)) & (~x0 | ~x1 | x2 | ~x4)));
  assign n1073 = (~n292 | ~n283 | ~n288) & (n777 | n705 | n1010);
  assign z062 = n1075 | ~n1078 | n1084 | n1087 | (~n437 & ~n1077);
  assign n1075 = x2 & ((~x1 & ~n1076) | (~n406 & ~n387));
  assign n1076 = (x4 | ~x7 | ((x0 | x3 | x5 | ~x6) & (~x0 | ~x5 | (x3 ^ ~x6)))) & (~x5 | x6 | x7 | x0 | x3 | ~x4);
  assign n1077 = (x3 | ~x4 | x5 | x0 | ~x1 | ~x2) & (x2 | ((x4 | ((~x0 | (x1 ? (~x3 | x5) : (x3 | ~x5))) & (x0 | x1 | x3 | x5))) & (x0 | ~x1 | x3 | ~x4 | ~x5)));
  assign n1078 = n1081 & (n1079 | n1083) & (x0 ? n1080 : n1082);
  assign n1079 = x4 ? (x5 | x6) : (~x5 | ~x6);
  assign n1080 = (x4 | x5 | ~x7 | ~x1 | ~x2 | x3) & (x1 | (~x3 ^ x4) | (x2 ? (x5 | ~x7) : (x5 ^ x7)));
  assign n1081 = x0 ? ((x3 | ~x5 | x7 | x1 | ~x2) & (~x1 | x2 | (x3 ? (~x5 | x7) : (x5 ^ x7)))) : (((~x2 ^ ~x7) | (x1 ? (~x3 | x5) : (x3 | ~x5))) & (x3 | x5 | (x1 ? (x2 | ~x7) : (~x2 | x7))));
  assign n1082 = ((~x3 ^ x4) | ((x1 | x2 | x5 | ~x7) & (~x1 | ~x2 | ~x5 | x7))) & (~x5 | ((~x2 | ((x4 | ~x7 | ~x1 | x3) & (~x4 | x7 | x1 | ~x3))) & (~x1 | x2 | (x3 ? (~x4 | ~x7) : (x4 | x7)))));
  assign n1083 = (~x0 | ~x1 | ~x2 | x3 | x7) & (~x3 | (x0 ? (x1 ? (x2 | ~x7) : (~x2 | x7)) : (x1 | (x2 ^ x7))));
  assign n1084 = ~n1085 & ~n1086;
  assign n1085 = x5 ^ ~x6;
  assign n1086 = (x0 | ~x1 | ~x2 | x3 | x4 | x7) & (~x3 | ((x2 | x4 | ~x7 | x0 | ~x1) & (x1 | ((x4 | x7 | x0 | ~x2) & (~x4 | (x0 ? (~x2 ^ ~x7) : (x2 | ~x7)))))));
  assign n1087 = ~x2 & ((~x3 & ~n1089) | (x3 & x5 & n321 & ~n1088));
  assign n1088 = x4 ? (~x6 | ~x7) : (x6 | x7);
  assign n1089 = x0 ? ((~x1 | ~x4 | ~x5 | x6 | x7) & (x1 | x5 | ((~x6 | ~x7) & (x4 | x6 | x7)))) : ((x1 | x4 | ~x5 | ~x6 | ~x7) & (~x1 | ~x4 | x5 | x6 | x7));
  assign z063 = (~x0 & ~n1091) | (x0 & ~n1092) | ~n1094 | (~n437 & ~n1093);
  assign n1091 = x6 ? ((x3 | ((~x1 | ~x4 | (x2 ^ ~x5)) & (x1 | x2 | x4 | x5))) & (x1 | ~x3 | (x2 ? (x4 | ~x5) : (~x4 | x5)))) : (x1 ? ((x2 | (x3 ? ~x4 : (x4 | x5))) & (~x2 | ~x3 | x4 | ~x5)) : (x3 | (x2 ? (~x4 ^ x5) : (~x4 | ~x5))));
  assign n1092 = x2 ? ((~x1 | x3 | x4 | x5 | x6) & (x1 | ((x5 | x6 | x3 | ~x4) & (~x3 | ~x6 | (~x4 ^ x5))))) : ((~x3 | ~x4 | ~x5 | (x1 ^ ~x6)) & (x4 | (x1 ? (x3 ? (x5 | ~x6) : (~x5 | x6)) : (x3 ? (x5 | x6) : ~x6))));
  assign n1093 = x4 ? (x2 ? ((x0 | ~x1 | ~x3) & (x1 | x3 | ~x5)) : ((~x1 | x3 | x5) & (~x0 | (x1 ? x3 : (~x3 | x5))))) : (((x0 & ~x2) | (x1 ? (x3 | ~x5) : (~x3 | x5))) & (x1 | x2 | ~x3 | ~x5) & (x0 | ~x1 | ~x2 | x3));
  assign n1094 = n1099 & (x2 | (~n1095 & ~n1097 & (n535 | n1098)));
  assign n1095 = ~n1096 & ((n595 & n611) | (n783 & n612));
  assign n1096 = x3 ^ ~x4;
  assign n1097 = ~n425 & (x0 ? n351 : n850) & (~x1 ^ x3);
  assign n1098 = (x3 | ~x5 | x6 | x7) & (~x3 | x5 | ~x6 | ~x7);
  assign n1099 = (~n1100 | n1103) & (x3 | n1102) & (~n354 | n1101);
  assign n1100 = ~x0 & x3;
  assign n1101 = x6 ? (~x7 | ((x3 | x4 | x5) & (~x0 | (x3 ? (~x4 | ~x5) : x4)))) : (x7 | ((~x3 | ~x4 | ~x5) & (x0 | (x3 ? ~x4 : (x4 | x5)))));
  assign n1102 = (x0 | ~x1 | ~x2 | ~x5 | ~x6 | ~x7) & (~x0 | x6 | x7 | (x1 ? (x2 | x5) : (~x2 | ~x5)));
  assign n1103 = (~x1 | ~x2 | x5 | x6 | x7) & (x1 | ~x6 | ~x7 | (x2 ^ ~x5));
  assign z064 = n1105 | n1108 | ~n1112 | (x0 & ~n1111);
  assign n1105 = ~x1 & (x4 ? ~n1107 : ~n1106);
  assign n1106 = x7 ? ((~x0 | x2 | x3 | ~x5 | ~x6) & (x0 | ~x3 | x6 | (x2 ^ ~x5))) : ((~x2 | ((x5 | ~x6 | x0 | ~x3) & (~x0 | (x3 ? (~x5 | ~x6) : (x5 | x6))))) & (x0 | x2 | x5 | (~x3 ^ x6)));
  assign n1107 = (~x7 | ((x0 | ~x2 | x3 | x5 | ~x6) & (x6 | ((~x3 | ~x5 | x0 | ~x2) & (x2 | (x0 ? (~x3 ^ x5) : (x3 | x5))))))) & (x2 | x3 | ~x6 | x7 | (~x0 ^ ~x5));
  assign n1108 = x1 & ((n865 & ~n1110) | (~x0 & ~n1109));
  assign n1109 = (~x2 | x4 | x6 | ~x7 | (x3 ^ ~x5)) & (x7 | ((x2 | ~x3 | ~x4 | x5 | ~x6) & (x3 | ~x5 | (x2 ? (~x4 ^ x6) : (x4 | x6)))));
  assign n1110 = (~x2 | x4 | x5 | ~x6 | ~x7) & (x2 | ((x4 | x5 | ~x6 | x7) & (x6 | (x4 ? (x5 ^ x7) : (x5 | ~x7)))));
  assign n1111 = (x7 | (x1 ? ((~x4 | ~x5 | x2 | ~x3) & (x4 | x5 | ~x2 | x3)) : (x2 | x4 | (~x3 ^ x5)))) & (~x2 | ~x5 | ~x7 | ((x3 | x4) & (x1 | ~x3 | ~x4)));
  assign n1112 = ~n1113 & n1116 & (n307 | n1115) & (n425 | n1114);
  assign n1113 = ~n699 & ((~x1 & ((~x0 & ~x2 & x3 & ~x5) | (x0 & (x2 ? ~x5 : (x3 & x5))))) | (~x0 & (x2 ? (~x3 & ~x5) : (x5 & (x1 | ~x3)))));
  assign n1114 = (~x5 | ((~x0 | ((x3 | ~x4 | x1 | ~x2) & (~x1 | x2 | ~x3 | x4))) & (x0 | x1 | x2 | ~x3 | ~x4))) & (x0 | ~x1 | ~x3 | x5 | (x2 ^ x4));
  assign n1115 = (x0 | ~x1 | x2 | x3 | x5) & ((~x1 ^ ~x3) | (x0 ? (x2 | x5) : (~x2 | ~x5)));
  assign n1116 = (n443 | n1117) & (~n313 | ~n615 | ~n992);
  assign n1117 = (~x0 | ~x1 | x2 | x3) & (x0 | x1 | ~x2 | ~x3);
  assign z065 = n1119 | n1122 | ~n1126 | ~n1128 | (~n416 & ~n1125);
  assign n1119 = ~x0 & (x7 ? ~n1121 : ~n1120);
  assign n1120 = x5 ? ((~x2 ^ ~x4) | (x1 ? (x3 | x6) : (~x3 | ~x6))) : ((~x3 | ((x1 | x2 | x4 | x6) & (~x1 | (x2 ? (x4 | ~x6) : (~x4 | x6))))) & (x1 | ~x2 | x3 | ~x4 | ~x6));
  assign n1121 = (~x4 | x5 | ~x6 | x1 | ~x3) & (x2 | x3 | (x5 ^ x6) | (~x1 ^ ~x4));
  assign n1122 = x0 & ((n354 & ~n1124) | (~x2 & ~n1123));
  assign n1123 = ((x4 ? (x5 | x7) : (~x5 | ~x7)) | (x1 ? (x3 | x6) : (~x3 | ~x6))) & (x3 | ~x5 | ~x6 | x7 | (~x1 ^ ~x4));
  assign n1124 = (x3 | ~x4 | x5 | ~x6 | ~x7) & (~x5 | ((x3 | x4 | x6 | ~x7) & (~x3 | (x4 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n1125 = x0 ? ((~x1 | x3 | x4) & (~x3 | ~x4 | x1 | x2)) : ((x1 | x3 | ~x4) & (~x3 | (x1 ? (x2 ^ x4) : (~x2 | x4))));
  assign n1126 = (x0 | n1127) & (n420 | ((x0 | ~x1 | ~x2 | x3) & (~x0 | x2 | (~x1 ^ ~x3))));
  assign n1127 = (x5 | ((~x1 | ((~x2 | ~x3 | x4 | x6) & (x2 | x3 | ~x6))) & (x4 | ~x6 | x1 | x3))) & (~x3 | ~x5 | (x1 ? (x2 | ~x4) : (x6 | (x2 & ~x4))));
  assign n1128 = (~x0 | n1129) & (n1130 | (x1 ? n589 : ~n548));
  assign n1129 = (x2 | x3 | ~x4 | ~x5 | x6) & (x1 | ((~x5 | x6 | x3 | ~x4) & (x5 | ~x6 | ~x3 | x4) & (~x2 | ((~x3 | ~x4 | x5) & (~x5 | ~x6 | x3 | x4)))));
  assign n1130 = (x0 | ~x2 | ~x3 | ~x5 | ~x7) & (x5 | ((~x0 | (x2 ? (x3 | x7) : (~x3 | ~x7))) & (x0 | ~x2 | x3 | ~x7)));
  assign z066 = ~n1143 | (x7 ? (n1138 | ~n1140) : ~n1132);
  assign n1132 = ~n1134 & ~n1136 & (x0 ? n1133 : (~n542 | ~n848));
  assign n1133 = (x1 | ~x2 | x3 | x4 | ~x5 | ~x6) & (x2 | ~x3 | ((x5 | x6 | x1 | x4) & (~x5 | (x1 ? (x4 ^ x6) : (~x4 | x6)))));
  assign n1134 = ~n1135 & (n509 | n929);
  assign n1135 = (x0 | ~x1 | ~x4 | ~x5 | ~x6) & (x5 | ((~x0 | ~x1 | (~x4 ^ x6)) & (x1 | ((~x4 | ~x6) & (x0 | x4 | x6)))));
  assign n1136 = ~n1137 & ((~x2 & ~x3 & x4 & ~x6) | (~x0 & ((~x4 & x6 & x2 & ~x3) | (~x2 & x4 & ~x6))));
  assign n1137 = x1 ^ ~x5;
  assign n1138 = ~n1139 & (x2 ? (x3 & ~n585) : n1070);
  assign n1139 = x0 ? (x1 | x5) : (~x1 | ~x5);
  assign n1140 = (x4 | (n1141 & (x6 | ~n357 | n1137))) & n1142 & (~x4 | ~x6 | ~n357 | n1137);
  assign n1141 = (x0 | x1 | x5 | (x2 ? (~x3 | x6) : ~x6)) & (~x0 | ~x1 | x2 | ~x5 | ~x6);
  assign n1142 = (~n992 | ~n552) & (~n358 | ~n451 | x1 | ~x4);
  assign n1143 = (n585 | n1145) & (~x2 | n1144) & (x1 | x2 | n389);
  assign n1144 = x4 ? (x6 | ((x1 | x3 | ~x7) & (x0 | ~x1 | x7))) : ((~x0 | x3 | x6 | (x1 ^ x7)) & (~x6 | ((x1 | ~x7) & (x0 | ~x1 | ~x3 | x7))));
  assign n1145 = (~x1 | x2 | (x3 ^ x7)) & (~x2 | ((x1 | ~x3 | x7) & (x0 | ~x1 | x3 | ~x7)));
  assign z067 = n1147 | ~n1149 | ~n1150 | ~n1153 | (~n1085 & ~n1148);
  assign n1147 = ~n1088 & ((x0 & ~x1 & x2 & n294) | (~x0 & ((~x2 & n335) | (x1 & x2 & n294))));
  assign n1148 = (x4 | ~x7 | x2 | ~x3) & (~x2 | x3 | ~x4 | x7 | (x0 & x1));
  assign n1149 = ((x5 ^ x7) | (x2 ? (x3 | x4) : (~x3 | ~x4))) & (~x3 | ~x5 | x7 | x0 | ~x2) & (x5 | ~x7 | x2 | x3);
  assign n1150 = (n416 | n1151) & (x4 | x7 | n1152);
  assign n1151 = (~x4 | x7 | x2 | x3) & (~x2 | ~x3 | x4 | ~x7 | (x0 & x1));
  assign n1152 = (~x0 | x6 | ((x1 | x2 | ~x3 | x5) & (~x1 | ~x2 | x3 | ~x5))) & (~x3 | x5 | ~x6 | x0 | ~x1 | ~x2);
  assign n1153 = ~n1155 & ~n1157 & (x0 ? (~x3 | n1154) : n1156);
  assign n1154 = (~x1 | x2 | x4 | x5 | x7) & (x1 | ~x2 | ((~x5 | x7) & (~x4 | x5 | ~x7)));
  assign n1155 = ~n617 & n783 & n654 & ~x3 & x7;
  assign n1156 = (x4 | ~x5 | x7 | x1 | x2 | x3) & (~x1 | ~x2 | ~x3 | ~x4 | x5 | ~x7);
  assign n1157 = ~n389 & ((x2 & x3 & ~x5 & n783) | (~x2 & ~x3 & x5 & ~n1158));
  assign n1158 = ~x0 & ~x1;
  assign z068 = (~x3 | ~n1165) & (x3 | n1160 | n1161 | ~n1162);
  assign n1160 = ~x0 & ((~x4 & ~x5 & x6) | (x1 & x4 & x5 & ~x6));
  assign n1161 = ~x1 & ((x5 & ~x6 & x7 & ~x0 & x4) | (~x5 & x6 & ~x7 & x0 & ~x4));
  assign n1162 = ~n1163 & n1164 & (n390 | (~x0 & ~x5) | (x5 & (x0 | x1)));
  assign n1163 = (~x6 ^ x7) & ((~x0 & x4 & ~x5) | (~x4 & x5 & (x0 | x1)));
  assign n1164 = ~x0 | ~x4 | ~x5 | (x1 & x2) | x6;
  assign n1165 = ~n1166 & n1169 & (x1 ? (x5 | n1171) : n1170);
  assign n1166 = ~n437 & ((~n950 & ~n1168) | (~x5 & ~n864 & n1167));
  assign n1167 = x0 & ~x4;
  assign n1168 = x2 & x0 & x1;
  assign n1169 = (x0 | (x4 ? (~x5 | ~x6) : (x5 | x6))) & (~x5 | ~x6 | x2 | ~x4) & (x1 | ((x5 | x6 | x2 | x4) & (~x4 | ~x5 | ~x6)));
  assign n1170 = (x0 | x4 | ~x5 | x6 | x7) & (~x0 | x5 | ((~x4 | ~x6 | ~x7) & (x6 | x7 | ~x2 | x4)));
  assign n1171 = (x0 | ~x2 | ~x4 | ~x6 | ~x7) & (~x0 | x2 | (x4 ? (~x6 | ~x7) : (x6 | x7)));
  assign z069 = ~n1178 | (x7 ? (n1173 | n1176) : (~n589 & ~n1177));
  assign n1173 = ~x0 & ((x1 & n358 & n1174) | (n268 & n1175));
  assign n1174 = x6 & x4 & ~x5;
  assign n1175 = ~x6 & ~x4 & x5;
  assign n1176 = n1041 & ((x1 & x2) ? (~x3 & n548) : ~n585);
  assign n1177 = x0 ? (x5 | (x1 ^ (~x2 | ~x3))) : (x1 | ~x5);
  assign n1178 = ~n1181 & ~n1180 & (x3 | x7 | ~n279 | n1179);
  assign n1179 = x1 ? (x4 | ~x5) : (~x4 | x5);
  assign n1180 = (x7 | (~x4 & (x0 | x1))) & (~x0 | ~x1 | ~x2) & x5 & (x4 | ~x7);
  assign n1181 = ~x5 & ((~x1 & ~x2 & x4 & ~x7) | (~x0 & (x4 ^ x7)));
  assign z070 = ~n1184 | n1189 | (~x1 & (~n1183 | ~n1188));
  assign n1183 = x0 ? (~x6 | ((x5 | ~x7) & (x2 | ~x5 | x7))) : (~x2 | x6 | (x5 ^ x7));
  assign n1184 = ~n1185 & ~n1186 & n1187 & (~n374 | ~n294 | ~n992);
  assign n1185 = x5 & ((~x6 & (x1 ? (~x0 | ~x2) : x0)) | (~x0 & x6 & (~x1 | ~x2)));
  assign n1186 = ~n950 & n358 & n349 & x6 & x7;
  assign n1187 = ~x1 | ~x6 | ((~x0 | x2 | x5) & (~x5 | x7 | x0 | ~x2));
  assign n1188 = (x7 | ((x0 | x2 | ~x3 | x5 | x6) & (~x0 | ~x2 | ~x6 | (~x3 ^ x5)))) & (x0 | x2 | x6 | ~x7 | (x3 ^ x5));
  assign n1189 = ~x3 & ((n1190 & n1192) | (~x6 & ~n1191));
  assign n1190 = x6 & ~x4 & ~x5;
  assign n1191 = (~x1 | x4 | ((~x0 | ~x2 | ~x5) & (x0 | x2 | x5 | x7))) & (x0 | x1 | x2 | ~x4 | (x5 ^ x7));
  assign n1192 = x2 & x0 & x1;
  assign z071 = ~n1196 | ~n1201 | (~x0 & (n1195 | (~x5 & ~n1194)));
  assign n1194 = (~x7 | (x1 ? ((x4 | x6 | x2 | x3) & (~x2 | ~x3 | ~x4 | ~x6)) : (x6 | (~x2 & ~x3)))) & (x1 | ~x6 | x7 | (~x2 & ~x3 & ~x4));
  assign n1195 = ~x1 & x5 & ~n437 & (x2 | n509 | n313);
  assign n1196 = ~n1198 & ~n1199 & n1200 & (~n358 | ~n321 | ~n1197);
  assign n1197 = ~x7 & ~x6 & ~x4 & ~x5;
  assign n1198 = ~n425 & ((n321 & (~x2 | ~x3)) | (x3 & n654 & n992));
  assign n1199 = ~x6 & n349 & ((n357 & n850) | (n351 & n358));
  assign n1200 = x1 | ~x6 | ((x3 | x4 | x0 | x2) & (~x0 | ~x2 | ~x3));
  assign n1201 = ~x1 | (x0 ? (~x6 | (x2 & (x3 | x4))) : (x6 | (x4 ? (x2 & x3) : (~x2 & ~x3))));
  assign z072 = n1203 | n1207 | ~n1208 | (~x0 & ~n1206);
  assign n1203 = ~x5 & (x4 ? ~n1205 : ~n1204);
  assign n1204 = x0 ? (x1 | ~x2 | ~x3 | (~x6 ^ x7)) : (x2 | x3 | ((~x6 | x7) & (~x1 | x6 | ~x7)));
  assign n1205 = (x0 | ((x1 | x2 | x3 | ~x6 | ~x7) & (~x1 | ~x2 | ~x3 | (x6 ^ x7)))) & (~x0 | ~x1 | ~x2 | x3 | x6 | x7);
  assign n1206 = (x2 | x3 | ((x4 | ~x5 | x7) & (x1 | ~x4 | (x5 ^ x7)))) & (~x1 | ~x2 | ~x3 | ~x4 | ~x5 | ~x7);
  assign n1207 = ~x7 & ((~x0 & x1 & ~x2 & ~x3 & x4) | (x2 & ((~x0 & x1 & x3 & ~x4) | (x0 & (x1 ? (~x3 & ~x4) : (x3 & x4))))));
  assign n1208 = (x2 & ((x1 & x3) | (x0 & (x1 | (x3 & ~n1209))))) | (~x0 & ((~x1 & ~x7) | (~x2 & ~x3))) | (x1 & x7) | (~x1 & ~x7 & (~x2 | ~n1209));
  assign n1209 = ~x7 & x5 & x3 & ~x4;
  assign z073 = n1211 | n1212 | n1214 | (x3 ? n706 : ~n1213);
  assign n1211 = ~x0 & ((~x1 & ((~x2 & x4 & x5) | (~x4 & ~x5 & x2 & ~x3))) | (~x2 & ((x1 & (x4 ^ x5)) | (~x3 & x4 & x5) | (x3 & (~x4 | ~x5)))) | (x1 & x2 & x3 & x4 & x5));
  assign n1212 = x0 & ((~x1 & (~x2 ^ (x3 & (x4 | x5)))) | (~x2 & ~x3 & (~x4 | ~x5)));
  assign n1213 = (~x4 | ~x5 | x6 | ~x0 | ~x1 | x2) & (x0 | x4 | ((x5 | ~x6 | ~x1 | x2) & (~x5 | x6 | x1 | ~x2)));
  assign n1214 = n783 & n1215 & (x2 ? (~x4 & n664) : (x4 & n870));
  assign n1215 = ~x3 & x6;
  assign z074 = ~n1217 | ~n1220 | (n783 & ~n1219) | (x6 & ~n1218);
  assign n1217 = x2 ? ((x0 | x1 | ~x3 | x4 | x5) & ((x3 ^ x5) | (x0 ? (x1 | x4) : (~x1 | ~x4)))) : ((x0 | x3 | ~x5 | (x1 ^ ~x4)) & (~x0 | ~x1 | ~x3 | ~x4 | x5));
  assign n1218 = (~x3 | (~x2 ^ x5) | (x0 ? (x1 | x4) : (~x1 | ~x4))) & (~x1 | x2 | x3 | (x0 ? (~x4 | ~x5) : (x4 | x5)));
  assign n1219 = (~x2 | x3 | x4 | ~x5 | ~x6 | ~x7) & (x2 | ~x4 | x5 | (x3 ? (x6 | x7) : (~x6 | ~x7)));
  assign n1220 = x0 ? ((~x1 | x2 | ~x3 | x4) & (x1 | ((~x3 | ~x4) & (x2 | x3 | x4)))) : ((x1 | x2 | ~x3 | x4) & (x3 | (x1 ? (~x2 ^ x4) : (~x2 | ~x4))));
  assign z075 = ~n1224 | n1234 | (~x4 & ~n1222) | (~x2 & ~n1235);
  assign n1222 = (x3 | n1223) & (~x3 | ~x6 | x7 | ~n349 | n750);
  assign n1223 = (x5 | ((x0 | x1 | x2 | x6 | ~x7) & (~x0 | x7 | (x1 ? (~x2 | ~x6) : (x2 | x6))))) & (x0 | ~x2 | ~x5 | (x1 ? (x6 | x7) : (~x6 | ~x7)));
  assign n1224 = ~n1225 & ~n1227 & n1228 & n1229 & (n798 | n1226);
  assign n1225 = ~x0 & ((x2 & ((~x4 & ~x5 & x1 & ~x3) | (~x1 & (x3 ? (~x4 & x5) : (x4 & ~x5))))) | (x1 & ~x2 & ~x4 & (x3 ^ x5)));
  assign n1226 = (~x4 | x5 | ~x7 | x0 | x1 | x2) & (~x0 | x7 | ((x4 | ~x5 | ~x1 | x2) & (x1 | ~x4 | (~x2 ^ x5))));
  assign n1227 = x4 & ((~x0 & x5 & (~x1 ^ x2)) | (x0 & ~x1 & ~x2 & ~x5));
  assign n1228 = ~x0 | ((x4 | ~x5 | x1 | ~x2) & (~x1 | x2 | ((x4 | x5) & (~x3 | ~x4 | ~x5))));
  assign n1229 = (n1232 | ~n1233) & (x6 | ~n1230 | ~n783 | n1231);
  assign n1230 = x2 & x4;
  assign n1231 = x3 ^ ~x5;
  assign n1232 = (~x1 | x2 | x3 | x6) & (~x3 | ~x6 | x1 | ~x2);
  assign n1233 = ~x7 & ~x5 & ~x0 & x4;
  assign n1234 = ~n750 & ((x1 & ((~x4 & ~x6 & x0 & ~x3) | (~x0 & x3 & (~x4 ^ x6)))) | (x0 & ~x1 & (x3 ? (~x4 & x6) : (x4 & ~x6))));
  assign n1235 = (~x4 | ~x5 | ~x6 | ~x0 | ~x1 | x3) & (x0 | x5 | ((x3 | x4 | ~x6) & (x1 | ~x3 | (x4 ^ x6))));
  assign z076 = ~n1238 | (x0 & ~n1245) | (~x0 & ~n1242) | (x1 & ~n1237);
  assign n1237 = (~x5 | ((x0 | x2 | ~x3 | ~x4 | ~x6) & (x6 | (x0 ? (x2 ? (x3 | x4) : (~x3 | ~x4)) : (x3 | (~x2 ^ ~x4)))))) & (x0 | x5 | ((x4 | ~x6 | x2 | ~x3) & (~x2 | (x3 ? (~x4 | ~x6) : (x4 | x6)))));
  assign n1238 = n1241 & (n665 | n1239) & (n1096 | n1240);
  assign n1239 = (~x0 | x1 | x2 | x3 | x4 | x6) & (x0 | ((x1 | ~x2 | ~x3 | ~x4 | ~x6) & (~x1 | ((x4 | ~x6 | ~x2 | ~x3) & (~x4 | x6 | x2 | x3)))));
  assign n1240 = (x0 | x1 | ~x2 | ~x5 | ~x6) & (~x0 | x2 | (x1 ? (~x5 | ~x6) : (x5 | x6)));
  assign n1241 = x0 ? ((~x1 | x2 | x3 | x5 | x6) & (x1 | (x2 ? (x3 ? (x5 | ~x6) : (~x5 | x6)) : (~x6 | (x3 ^ x5))))) : (x2 ? (x3 ? (~x5 | x6) : (x1 ? (~x5 | ~x6) : (x5 | x6))) : ((~x5 | x6 | x1 | x3) & (x5 | (x1 ? (~x3 ^ x6) : (~x3 | ~x6)))));
  assign n1242 = x1 ? (n1243 | (x2 ? (x3 | x6) : (~x3 | ~x6))) : n1244;
  assign n1243 = x4 ? (x5 | x7) : (~x5 | ~x7);
  assign n1244 = (~x2 | x3 | x4 | ~x5 | ~x6 | ~x7) & ((x3 ^ ~x6) | ((~x2 | x4 | x5 | x7) & (x2 | (x4 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n1245 = ~n1246 & (x1 | ~n509 | ~n339) & (~x1 | ~x6 | n442);
  assign n1246 = ~n798 & ((~x2 & ((x5 & x7 & ~x1 & x4) | (x1 & ~x4 & (~x5 ^ x7)))) | (~x1 & x2 & (x4 ? (~x5 & x7) : (x5 & ~x7))));
  assign z077 = ~n1258 | (x0 ? (n1249 | (~x2 & ~n1248)) : ~n1250);
  assign n1248 = x4 ? ((x1 | ~x3 | (~x6 ^ x7)) & (~x1 | x3 | ~x5 | ~x6 | x7)) : (((~x1 ^ ~x3) | ((x6 | ~x7) & (x5 | ~x6 | x7))) & (x1 | ~x3 | x5 | x6 | x7));
  assign n1249 = n354 & ((x3 & x4 & ~x5 & (x6 ^ x7)) | (x5 & ((~x4 & (x3 ? (x6 ^ x7) : (x6 & x7))) | (~x6 & ~x7 & ~x3 & x4))));
  assign n1250 = n1254 & (n1253 | (~n1251 & ~n1252));
  assign n1251 = x3 & ~x1 & ~x2;
  assign n1252 = ~x3 & x1 & x2;
  assign n1253 = (~x4 | x5 | x6 | ~x7) & (x4 | ((~x6 | x7) & (~x5 | x6 | ~x7)));
  assign n1254 = (~x6 | n1257) & (n437 | n1256) & (x2 | x6 | n1255);
  assign n1255 = (x1 | x3 | x4 | x5 | ~x7) & (~x1 | x7 | (x3 ? (~x4 | ~x5) : (x4 | x5)));
  assign n1256 = (~x1 | x2 | x3 | ~x4) & (x1 | ~x2 | ~x3 | x4 | x5);
  assign n1257 = (~x4 | x5 | ~x7 | x1 | ~x2 | ~x3) & (~x5 | (~x1 ^ ~x3) | (x2 ? (~x4 | x7) : (x4 | ~x7)));
  assign n1258 = ~n1261 & n1262 & (n425 | n1259) & (x1 | n1260);
  assign n1259 = ((~x1 ^ ~x3) | ((~x4 | ~x5 | ~x0 | x2) & (x0 | (x2 ? x4 : (~x4 | x5))))) & (~x3 | ~x4 | ~x5 | x0 | x1 | ~x2) & (~x0 | x3 | ((~x4 | x5 | x1 | ~x2) & (~x1 | x4 | (x2 & x5))));
  assign n1260 = (~x4 | x5 | x6 | ~x0 | x2 | x3) & (x4 | (x0 ? (x5 | (x2 ? (x3 | x6) : (~x3 | ~x6))) : (~x5 | x6 | (x2 ^ x3))));
  assign n1261 = ~n798 & ((~x0 & x1 & ~x2 & ~x4) | (x4 & (x0 ? (x1 ? (~x2 & ~x5) : (x2 & x5)) : (~x1 & (x2 ^ x5)))));
  assign n1262 = (n1071 | n1263) & (~n531 | ~n288 | ~n524);
  assign n1263 = (~x5 | ~x6 | x2 | ~x3) & (~x2 | (x3 ? (x5 | ~x6) : (~x5 | x6)));
  assign z078 = n1265 | ~n1270 | (~n699 & ~n1269) | (~x4 & ~n1268);
  assign n1265 = x1 & (~n1267 | (~x0 & ~n1266));
  assign n1266 = (x5 | ~x6 | x7 | x2 | x3 | x4) & (x6 | ((~x4 | ((x2 | x3 | ~x5 | ~x7) & (~x2 | (x3 ? (~x5 | x7) : (x5 | ~x7))))) & (x2 | ~x3 | x4 | ~x5 | x7)));
  assign n1267 = (~x0 | x2 | ~x3 | ~n511) & ((~n697 & ~n1197) | (x0 ? (x2 | x3) : (~x2 | ~x3)));
  assign n1268 = x0 ? ((x5 | ~x7 | x2 | x3) & (x7 | ((~x1 | ~x2 | x3 | ~x5) & (x1 | ~x3 | (~x2 ^ x5))))) : (x1 | (x2 ? ((x5 | ~x7) & (~x3 | ~x5 | x7)) : (~x3 | (x5 ^ x7))));
  assign n1269 = x1 ? ((x3 | x5 | (x0 ? (~x2 | x6) : (~x2 ^ ~x6))) & (x0 | x2 | ~x3 | ~x5 | ~x6)) : (x0 ? ((x5 | x6 | x2 | ~x3) & (~x5 | ~x6 | ~x2 | x3)) : ((x5 | ~x6 | x2 | ~x3) & (~x5 | x6 | ~x2 | x3)));
  assign n1270 = ~n1271 & ~n1275 & ~n1276 & (~x4 | n1274);
  assign n1271 = ~x1 & (x6 ? ~n1273 : (~n1272 & (x0 ^ ~x2)));
  assign n1272 = (x3 | x4 | ~x5 | x7) & (~x3 | ~x4 | x5 | ~x7);
  assign n1273 = ((~x3 ^ x5) | ((x0 | ~x2 | ~x4 | ~x7) & (~x0 | x2 | x4 | x7))) & (x0 | x2 | x3 | x4 | (x5 ^ x7));
  assign n1274 = (x1 | ((~x5 | x7 | x0 | x2) & (~x2 | ((~x0 | (x3 ? (~x5 | x7) : (x5 | ~x7))) & (x5 | x7 | x0 | ~x3))))) & (x0 | x2 | x5 | ~x7 | (~x1 & x3));
  assign n1275 = ~n1231 & ((x0 & ~x1 & ~x2 & x4 & x7) | (x1 & ((~x4 & ~x7 & ~x0 & ~x2) | ((x4 ^ x7) & (~x0 ^ ~x2)))));
  assign n1276 = ~n1277 & (x0 ? ((~x2 & x4) | (~x1 & x2 & ~x4)) : (x2 & (~x1 ^ ~x4)));
  assign n1277 = x3 ? (~x5 | ~x7) : (x5 | x7);
  assign z079 = ~n1290 | n1289 | n1287 | n1286 | n1279 | n1283;
  assign n1279 = x0 & ((n1280 & ~n1282) | (x6 & ~n1281));
  assign n1280 = ~x2 & ~x6;
  assign n1281 = x1 ? ((x4 | x5 | ~x7 | ~x2 | x3) & (x2 | ~x4 | (x3 ? (~x5 | x7) : (x5 ^ x7)))) : ((x2 | x3 | ~x4 | ~x5 | x7) & (~x2 | ((x5 | x7 | x3 | x4) & (~x3 | (x4 ? (x5 | ~x7) : (~x5 | x7))))));
  assign n1282 = ((~x1 ^ x7) | (x3 ? (~x4 | x5) : (x4 | ~x5))) & (~x1 | x4 | ~x7 | (~x3 ^ ~x5));
  assign n1283 = ~x0 & (x7 ? ~n1284 : ~n1285);
  assign n1284 = x5 ? ((x1 | ~x2 | x3 | x4 | ~x6) & (~x1 | x2 | ~x3 | ~x4 | x6)) : (x4 ? ((~x1 | x2 | x3 | x6) & (x1 | ~x2 | ~x3 | ~x6)) : (x1 ? (~x2 | (~x3 ^ x6)) : (x2 | (~x3 ^ ~x6))));
  assign n1285 = ((x2 ^ x6) | ((~x4 | ~x5 | x1 | ~x3) & (~x1 | (x3 ? (~x4 | x5) : (x4 | ~x5))))) & (x6 | ((~x1 | ~x2 | x3 | ~x4 | ~x5) & (x1 | x5 | (x2 ? (~x3 | x4) : (x3 | ~x4)))));
  assign n1286 = ~n399 & ((~x6 & ((~x1 & x2) | (x0 & (x1 ? (~x2 & x4) : ~x4)))) | (~x4 & x6 & x1 & ~x2) | (~x0 & (x1 ? (x4 & x6) : (x2 & ~x4))));
  assign n1287 = ~n589 & ((~x0 & ~n1288) | (~x2 & n321 & n294));
  assign n1288 = (~x1 | ~x2 | ~x3 | x5) & (x1 | x2 | x3 | ~x5);
  assign n1289 = x5 & n837 & (x3 ? (~x4 & ~x6) : (x4 & x6));
  assign n1290 = (n1291 | n1294) & (n1293 | (~n1292 & (~n313 | ~n615)));
  assign n1291 = x2 ? (x3 | ~x5) : (~x3 | x5);
  assign n1292 = ~x7 & ~x5 & x3 & ~x4;
  assign n1293 = (x0 | ~x1 | x2 | ~x6) & (~x0 | x1 | ~x2 | x6);
  assign n1294 = x1 ? (x4 | x6) : (~x6 | (~x0 & ~x4));
  assign z080 = ~n1296 | ~n1305 | (~n416 & ~n1304) | (~n425 & ~n1303);
  assign n1296 = ~n1297 & ~n1299 & ~n1300 & n1302 & (n307 | n1298);
  assign n1297 = ~n437 & (x2 ? (n349 & ~n946) : (~n858 & ~n1179));
  assign n1298 = x0 ? (x3 | ((x5 | ~x6 | ~x1 | x2) & (~x5 | x6 | x1 | ~x2))) : (x1 | ~x3 | (x2 ? (x5 | ~x6) : (~x5 | x6)));
  assign n1299 = ~x2 & (((x4 ? (x5 & ~x6) : (~x5 & x6)) & (x0 ^ ~x3)) | (x0 & ~x3 & x4 & ~x5 & ~x6) | (~x0 & x3 & ~x4 & x5 & x6));
  assign n1300 = ~x2 & ~n1301 & (x1 ? (~x6 & x7) : (x6 & ~x7));
  assign n1301 = x0 ? (x3 | x4) : (~x3 | ~x4);
  assign n1302 = (~n463 | ~n786) & (~n543 | ~n313 | ~n459);
  assign n1303 = x2 ? ((x0 | ~x1 | ~x3 | ~x4 | x5) & ((x0 ^ ~x5) | ((x3 | x4) & (x1 | ~x3 | ~x4)))) : ((~x4 | ~x5 | ~x0 | x3) & (x4 | x5 | x0 | ~x3));
  assign n1304 = (~x4 | ((x0 | x3 | (x1 ? (x2 | ~x7) : (~x2 | x7))) & (~x0 | ~x1 | x2 | ~x3 | ~x7))) & (~x0 | x1 | ~x3 | x4 | (~x2 ^ ~x7));
  assign n1305 = (~x2 | n1306) & (x0 | (~n1308 & (x4 | n1307)));
  assign n1306 = ((x0 ? (~x5 | ~x6) : (x5 | x6)) | ((x3 | x4) & (x1 | ~x3 | ~x4))) & (x4 | ~x5 | x6 | x1 | ~x3) & (x0 | ((x5 | ~x6 | x3 | ~x4) & (~x3 | ~x5 | ((x4 | x6) & (~x1 | ~x4 | ~x6)))));
  assign n1307 = (x1 | ((x2 | x3 | ~x5 | ~x6 | x7) & (~x2 | ~x3 | x5 | x6 | ~x7))) & (x5 | ~x6 | ~x7 | ~x1 | ~x2 | x3);
  assign n1308 = n367 & n369 & (x2 ? n451 : n450);
  assign z081 = ~n1310 | n1315 | ~n1317 | (x1 & ~n1314);
  assign n1310 = ~n1312 & (x0 | n1311) & (x1 | n1313);
  assign n1311 = (x6 | (x1 ? ((~x5 | x7 | x3 | ~x4) & (x5 | ~x7 | ~x3 | x4)) : (x3 | (x4 ? (x5 | ~x7) : (~x5 | x7))))) & (~x3 | ~x4 | ~x6 | (x1 ? (~x5 | x7) : (x5 | ~x7)));
  assign n1312 = ~n406 & ((~x0 & x1 & ~x4 & x5) | (x0 & ((x4 & x5 & ~x1 & x2) | (x1 & ~x2 & (~x4 ^ x5)))));
  assign n1313 = x0 ? ((x2 | ~x5 | (x3 ? (x4 | x7) : (~x4 | ~x7))) & (x3 | x5 | ((~x4 | x7) & (~x2 | x4 | ~x7)))) : (((x5 ^ x7) | (x2 ? (x3 | x4) : (~x3 | ~x4))) & (~x5 | x7 | x3 | ~x4) & (x4 | x5 | ~x7 | x2 | ~x3));
  assign n1314 = (x0 | ((x5 | ~x7 | ~x3 | ~x4) & (x3 | ((x4 | x5 | x7) & (~x2 | ((x5 | x7) & (~x4 | ~x5 | ~x7))))))) & (x4 | ~x5 | ~x7 | ~x0 | x2 | ~x3);
  assign n1315 = x6 & ((n992 & n993) | (~x2 & ~n1316));
  assign n1316 = (x4 | ~x5 | x7 | x0 | x1 | ~x3) & ((x5 ^ x7) | ((x0 | x1 | x3 | x4) & (~x0 | ~x1 | ~x3 | ~x4)));
  assign n1317 = (~x0 | n1320) & (n665 | n1319) & (n798 | n1318);
  assign n1318 = x0 ? ((x4 | x5 | ~x7 | x1 | x2) & ((x4 ? (x5 | ~x7) : (~x5 | x7)) | (x1 ^ ~x2))) : (~x4 | (x5 ^ x7) | (x1 ^ ~x2));
  assign n1319 = (x0 | x1 | ~x2 | ~x3 | x4) & (~x0 | ((~x1 | ~x2 | x3 | x4) & (~x3 | ~x4 | x1 | x2)));
  assign n1320 = (~x1 | x3 | ~x4 | x5 | x6 | x7) & (x1 | x4 | (x5 ^ x7) | (~x3 ^ ~x6));
  assign z082 = n1322 | n1325 | ~n1329 | (~n437 & ~n1328);
  assign n1322 = x3 & (x2 ? ~n1324 : ~n1323);
  assign n1323 = x1 ? ((x6 ^ x7) | (x0 ? (~x4 | ~x5) : (x4 | x5))) : (x0 ? ((x6 | x7 | ~x4 | x5) & (~x6 | ~x7 | x4 | ~x5)) : (x4 ? (x5 ? (x6 | x7) : (~x6 | ~x7)) : (x5 ? (x6 | ~x7) : (~x6 | x7))));
  assign n1324 = (x5 | ~x6 | ~x7 | ~x0 | x1 | ~x4) & (x0 | ((x1 | ~x4 | ~x5 | ~x6 | ~x7) & (x4 | ((~x6 | x7 | x1 | ~x5) & (~x1 | (x5 ? (x6 | x7) : (~x6 | ~x7)))))));
  assign n1325 = ~x3 & (x1 ? ~n1327 : ~n1326);
  assign n1326 = x4 ? ((~x6 | (x0 ? (x2 ? (x5 | ~x7) : (~x5 | x7)) : (~x7 | (~x2 ^ ~x5)))) & (~x2 | x6 | x7 | (x0 ^ ~x5))) : ((x6 | ((x0 | ~x2 | ~x5 | ~x7) & (~x0 | (x2 ? (x5 | ~x7) : (~x5 | x7))))) & (~x0 | x2 | ~x5 | ~x6 | ~x7));
  assign n1327 = ((~x2 ^ ~x5) | ((~x6 | x7 | ~x0 | x4) & (x6 | ~x7 | x0 | ~x4))) & ((~x4 ^ x7) | ((x0 | ~x2 | x5 | ~x6) & (~x0 | x2 | ~x5 | x6))) & (x0 | x2 | x4 | x7 | (x5 ^ x6));
  assign n1328 = (~x3 | (x0 ? (x4 | (x1 ? (x2 | ~x5) : (~x2 | x5))) : (~x1 | ~x4 | (~x2 ^ ~x5)))) & (x0 | x1 | x2 | x3 | x4 | x5);
  assign n1329 = ~n1331 & ~n1332 & ((x6 & (x2 | n1333)) | (n1330 & ((~x2 & ~x6) | n1333)));
  assign n1330 = (x5 | ((~x0 | ~x1 | ~x2 | x3 | x4) & (x0 | ~x3 | (x1 ? (~x2 | ~x4) : (x2 | x4))))) & (x1 | ~x4 | ((x2 | x3 | ~x5) & (~x0 | (~x5 & (x2 | x3)))));
  assign n1331 = x6 & n384 & ((x0 & (x2 ^ ~x5)) | (~x3 & (~x0 ^ ~x5)));
  assign n1332 = ~n585 & ((~x0 & ~x1 & x2 & ~x5) | (x1 & (x0 ? (~x2 & ~x5) : (x5 & (~x2 | ~x3)))));
  assign n1333 = (~x0 | ~x1 | x3 | x4 | ~x5) & (x0 | ((x4 | ~x5 | x1 | ~x3) & (~x1 | x3 | ~x4 | x5)));
  assign z083 = n1335 | ~n1339 | (~n440 & ~n1338);
  assign n1335 = x3 & ((n1336 & n352) | (~x1 & ~n1337));
  assign n1336 = ~x2 & x0 & x1;
  assign n1337 = (x4 | ((x6 | ((x0 | (x2 ? (~x5 | x7) : (x5 | ~x7))) & (~x0 | ~x2 | x5 | ~x7))) & (x0 | x2 | ~x5 | ~x6 | x7))) & (~x0 | x2 | ~x4 | (x5 ? (~x6 | x7) : (x6 | ~x7)));
  assign n1338 = x0 ? ((~x1 | ((x2 | x6) & (x4 | ~x6 | ~x2 | x3))) & (x2 | (x6 ? (x1 & ~x3) : x3))) : ((~x1 | ((~x2 | ~x4 | x6) & (x4 | ~x6 | x2 | x3))) & (x1 | x2 | ~x3 | x6) & (~x2 | (((x1 & ~x3) | (x4 ^ x6)) & (x3 | ~x4 | x6) & (x1 | ~x3 | ~x6))));
  assign n1339 = ~n1342 & n1344 & (x3 | n1340) & (~x4 | n1343);
  assign n1340 = (n665 | n1341) & (~n284 | ~n460);
  assign n1341 = (x0 | x1 | x2 | x4 | x6) & (~x0 | ~x6 | (x1 ? (x2 | x4) : (~x2 | ~x4)));
  assign n1342 = ~n665 & ((~x1 & ((~x3 & x6 & ~x0 & ~x2) | (x0 & x2 & (~x3 ^ x6)))) | (~x0 & x1 & (~x2 ^ (~x3 & x6))));
  assign n1343 = (x0 | x1 | x2 | x3 | x5 | x6) & ((~x0 ^ x5) | ((~x3 | x6 | x1 | ~x2) & (x3 | ~x6 | ~x1 | x2)));
  assign n1344 = (~x3 | n1346) & (~x2 | x3 | x4 | n1054 | n1345);
  assign n1345 = x1 ^ ~x6;
  assign n1346 = (~x5 | x6 | x7 | ~x0 | x1 | x2) & (x0 | x5 | ~x6 | ~x7 | (x1 ^ x2));
  assign z084 = ~n1357 | n1353 | n1352 | ~n1351 | n1348 | n1350;
  assign n1348 = ~n437 & ~n1349;
  assign n1349 = (x3 | x4 | x1 | ~x2) & (~x1 | ((~x4 | ~x5 | x2 | x3) & (~x3 | ((x0 | ~x2 | (~x4 ^ x5)) & (~x0 | x2 | x4 | x5)))));
  assign n1350 = ~x3 & (x1 ? (~x6 & ((~x0 & x2 & x4) | (~x2 & ~x4))) : (x6 & (~x2 ^ x4)));
  assign n1351 = (~x4 | x5 | x6 | ~x1 | x2 | x3) & (x1 | ~x3 | x4 | (x2 ? (x5 | ~x6) : (~x5 | x6)));
  assign n1352 = ~x2 & x3 & (x1 ? (x6 & (x0 ^ ~x4)) : (x4 & ~x6));
  assign n1353 = x3 & (n1356 | (n278 & ~n1355 & ~x6 & n1354));
  assign n1354 = ~x4 & ~x5;
  assign n1355 = ~x1 ^ ~x7;
  assign n1356 = n654 & ~n1042 & ((~x1 & ~x7) | (~x0 & x1 & x7));
  assign n1357 = ~n1360 & (n425 | n1359) & (x5 | ~n313 | n1358);
  assign n1358 = (~x1 | x2 | ~x6 | x7) & (~x0 | ((~x1 | ~x2 | x6 | x7) & (~x6 | ~x7 | x1 | x2)));
  assign n1359 = (~x1 | ~x2 | x3 | x4) & (x1 | ((~x3 | ((~x2 | (~x4 ^ x5)) & (~x0 | x2 | x4 | x5))) & (x2 | x3 | ~x4 | (x0 & ~x5))));
  assign n1360 = n367 & ((x0 & ~x2 & ~x4 & x5 & x6) | (~x0 & ((~x5 & x6 & ~x2 & x4) | (x2 & (x4 ? (x5 & x6) : (~x5 & ~x6))))));
  assign z085 = n1363 | ~n1364 | (~x7 & ~n1362);
  assign n1362 = (~x2 | ~x3 | x4 | ~x5 | (x0 & x1)) & (x5 | (x3 ? ((x0 | ~x2 | ~x4) & (x2 | x4)) : ((~x0 | x1 | ~x2 | x4) & (x0 | (x1 ? (~x2 | x4) : (x2 | ~x4))))));
  assign n1363 = x2 & ((~x7 & ((~x0 & ~x1 & ~x3 & ~x4) | (x0 & (x1 ? (~x3 & ~x4) : (x3 & x4))))) | (~x3 & x4 & x7 & (~x0 | ~x1)));
  assign n1364 = n1366 & ~n1371 & (n1042 | n1365) & (x0 | n1369);
  assign n1365 = (x0 | ~x3 | ((~x4 | ~x5 | x7) & (x5 | ~x7 | x1 | x4))) & (x3 | ~x4 | x5 | (~x0 & ~x1) | x7);
  assign n1366 = n1368 & (n1367 | (x2 ? (x4 | (x0 ^ ~x1)) : ~x4));
  assign n1367 = x3 ? (x5 | ~x7) : (~x5 | x7);
  assign n1368 = x2 | x4 | ~x7 | (x3 & ~x5);
  assign n1369 = (x5 | n1370) & (~x3 | ~x4 | ~x5 | ~x7 | n617);
  assign n1370 = (~x4 | x6 | x7 | x1 | ~x2 | x3) & (x4 | ~x6 | ~x7 | ~x1 | x2 | ~x3);
  assign n1371 = n654 & n545 & ((~x1 & x6 & (x2 ^ ~x7)) | (~x2 & ~x6 & x7));
  assign z086 = ~n1375 | (~x3 & (n1374 | (~x5 & ~n1373)));
  assign n1373 = (~x1 | ((x0 | ~x2 | x4 | ~x6 | ~x7) & (~x0 | x2 | ~x4 | (~x6 & ~x7)))) & (x0 | x1 | x6 | x7 | (~x2 ^ x4));
  assign n1374 = x5 & n432 & ((~x1 & x2 & x6 & ~x7) | (x1 & ~x2 & (~x6 | ~x7)));
  assign n1375 = ~n1378 & n1379 & (~n509 | n1376) & (x1 | n1377);
  assign n1376 = (x0 | ~x1 | x4 | x5 | ~x6 | ~x7) & (~x0 | ((~x4 | x7 | (x1 ? (x5 | x6) : (~x5 | ~x6))) & (~x1 | ~x5 | (x4 & (~x6 | ~x7)))));
  assign n1377 = (~x0 | ~x3 | ~x4 | ~x5 | ~x6 | ~x7) & (x5 | (x3 ? ((~x4 | x6 | x7) & (~x6 | ~x7 | x0 | x4)) : ((~x4 | x6 | ~x7) & (x0 | ((x6 | ~x7) & (x4 | ~x6 | x7))))));
  assign n1378 = ~x5 & n349 & ((n372 & n361) | (~x3 & ~n389));
  assign n1379 = ((x0 & x1) | (x3 ? (x4 | ~x5) : (~x4 | (~x5 ^ x6)))) & (~x5 | ~x6 | x0 | ~x3) & (x3 | x4 | x5 | (~x0 & (~x1 | x6)));
  assign z087 = n1381 | n1385 | ~n1386 | ~n1389 | (~n307 & ~n1384);
  assign n1381 = ~x3 & ((~x4 & ~n1382) | (n1383 & (~x1 | n542)));
  assign n1382 = x0 ? (~x1 | ~x2 | x7 | (x5 ^ x6)) : (x5 | ~x6 | (x1 & x2) | ~x7);
  assign n1383 = ~x7 & x6 & ~x5 & ~x0 & x4;
  assign n1384 = (~x0 & (x6 | (~x1 & ~x2 & ~x3))) | (x6 & (~x5 | (~x1 & ~x2))) | (x0 & x1 & x2) | (x5 & ~x6);
  assign n1385 = (~x0 ^ ~x2) & (x4 ? (x6 & (~x1 ^ ~x5)) : (x5 & ~x6));
  assign n1386 = n1387 & (~n351 | ~n278 | (x1 ? (~x3 | ~x6) : (x3 | x6)));
  assign n1387 = (x6 | ~n850 | x0 | x2) & (~x0 | ~x2 | (x1 ? ~n1388 : (x6 | ~n850)));
  assign n1388 = ~x6 & x5 & ~x3 & ~x4;
  assign n1389 = ~n1390 & (~n547 | (x0 ? (x1 | x5) : (~x5 | (~x1 & x2))));
  assign n1390 = n450 & n1100 & ((~x1 & ~n699) | (n542 & n370));
  assign z088 = ~n1397 | n1396 | n1395 | n1392 | n1393;
  assign n1392 = ~x1 & ((~x0 & ((~x5 & x7) | (x2 & x5 & ~x7))) | (x6 & ~x7 & ((~x2 & x5) | (x0 & x2 & ~x5))));
  assign n1393 = ~x3 & ((~x6 & ~n1394) | (~n440 & n1192 & ~x4 & x6));
  assign n1394 = (~x0 | ~x1 | ~x2 | x4 | (~x5 ^ x7)) & (x0 | x1 | x2 | ~x4 | x7);
  assign n1395 = x1 & ((~x5 & x6 & ~x7 & x0 & ~x2) | (~x0 & ((x5 & x6 & ~x7) | (~x2 & (x5 ? ~x7 : (~x6 & x7))))));
  assign n1396 = n278 & ((~x1 & x3 & x5 & ~x6 & ~x7) | (x1 & x6 & x7 & (~x3 ^ x5)));
  assign n1397 = ~n1398 & (~n509 | ~n349 | ~n352);
  assign n1398 = (x0 | (x1 & x2)) & (x5 | (~x6 & x7)) & (~x6 | x7) & (~x0 | ~x1 | ~x2) & (~x5 | x6 | ~x7);
  assign z089 = ~n1401 | ~n1402 | ~n1403 | (n278 & ~n1400);
  assign n1400 = (x5 | x6 | x7 | x1 | x3 | ~x4) & (x4 | ((x1 | x3 | ~x5 | x6 | x7) & (~x1 | ~x3 | ~x7 | (~x5 ^ x6))));
  assign n1401 = (~x0 | x6 | (x1 ^ ~x2)) & (~n958 | ~n339) & (x0 | x1 | ~x2 | ~x6);
  assign n1402 = ~x6 | ~n278 | (x3 ? (x1 & (x4 | x7)) : (~x1 & (x4 | ~x7)));
  assign n1403 = ~n1404 & (n437 | (x0 ? (x1 | x2) : (~x1 | (~x2 & ~n361))));
  assign n1404 = ~x3 & ((~x0 & ~x1 & ~x2 & x4 & x6) | (x0 & x1 & x2 & ~x4 & ~x6));
  assign z090 = ~n1408 | (n345 & ~n1406) | (n278 & ~n1407);
  assign n1406 = (x5 | ~x6 | x7 | x0 | x3 | x4) & (~x4 | ((x0 | x3 | x5 | (x6 ^ x7)) & (~x0 | ~x3 | ~x5 | ~x6 | ~x7)));
  assign n1407 = (x1 | x3 | ~x4 | ~x5 | ~x7) & (x4 | ((x1 | x3 | ~x5 | x7) & (~x1 | ~x3 | (~x5 ^ x7))));
  assign n1408 = (x0 | (x1 ? (x7 | (~x2 & (~x3 | ~x4))) : (~x3 | ~x7))) & (~x0 | x1 | x2 | x7) & (~x7 | ((x1 | ~x2) & (~x1 | x2 | x3) & (~x0 | (x2 ? (x3 | x4) : ~x1))));
  assign z091 = n1412 | ~n1413 | n1416 | (x4 & (~n1410 | ~n1417));
  assign n1410 = (x0 | ~x6 | ~x7 | ~n354 | ~n294) & (~x0 | x7 | n1411);
  assign n1411 = (x1 | x2 | ~x3 | ~x5 | ~x6) & (~x1 | ~x2 | x3 | x5 | x6);
  assign n1412 = x0 & ((~x1 & ~x2 & x3 & ~x4) | (x1 & ~x3 & (x2 ^ x4)));
  assign n1413 = (x2 | (x0 ? (~x1 ^ ~x3) : (~x1 | x3))) & n1414 & (x0 | ~x2 | ~x3 | (x1 & ~n654));
  assign n1414 = (~n269 | ~n1415) & (~n450 | ~n288 | ~n317);
  assign n1415 = ~x3 & ~x2 & ~x0 & ~x1;
  assign n1416 = ~x2 & (x0 ? ((x4 & ~x5 & ~x1 & x3) | (~x4 & x5 & x1 & ~x3)) : (~x4 & (x1 ? (x3 & ~x5) : (~x3 & x5))));
  assign n1417 = (~x3 | ~x5 | x6 | ~x0 | x1 | x2) & (x0 | x5 | ((x1 | x2 | x3 | x6) & (~x1 | ~x2 | ~x3 | ~x6)));
  assign z092 = ~n1426 | ~n1424 | n1423 | n1421 | n1419 | n1420;
  assign n1419 = ~x0 & ((~x3 & ~x4 & ~x1 & x2) | (x1 & ((~x3 & x4) | (x2 & x3 & ~x4))));
  assign n1420 = ~x1 & (x2 ? ((~x4 & x5 & x0 & x3) | (x4 & ~x5 & ~x0 & ~x3)) : ((~x4 & x5 & ~x0 & ~x3) | (x4 & (x0 ? (x3 ^ x5) : (x3 & x5)))));
  assign n1421 = ~x1 & ~n1422;
  assign n1422 = x0 ? (~x3 | ((~x5 | x6 | x2 | ~x4) & (x5 | ~x6 | ~x2 | x4))) : (x3 | ((~x5 | x6 | ~x2 | ~x4) & (x2 | x5 | (~x4 ^ x6))));
  assign n1423 = x0 & (x1 ? (x2 ? (~x3 & ~x4) : (x3 & x4)) : (x3 & (~x2 ^ x4)));
  assign n1424 = ~n1425 & (x4 | ~n542 | (x0 ? ~n784 : n1231));
  assign n1425 = ~x5 & n349 & (x4 ? (~x6 & n358) : (x6 & n357));
  assign n1426 = (~x5 | ~x6 | n533 | n1427) & (x3 | x5 | x6 | n1428);
  assign n1427 = x0 ? (x2 | ~x3) : (~x2 | x3);
  assign n1428 = (x0 | x1 | x2 | x4 | ~x7) & (~x0 | ~x1 | ~x2 | ~x4 | x7);
  assign z093 = n1430 | n1433 | ~n1435 | (x3 & x6 & ~n1432);
  assign n1430 = ~x2 & ~n1431;
  assign n1431 = x1 ? ((~x0 | x3 | ~x4 | ~x5 | ~x6) & (x4 | ((x5 | (~x3 & x6)) & (~x0 | (x5 & (~x3 | x6)))))) : ((~x4 | ((x5 | (~x3 & x6)) & (~x0 | (x5 & (~x3 | x6))))) & (x0 | x4 | (~x5 & (x3 | ~x6))));
  assign n1432 = (x4 | x5 | ~x7 | x0 | x1 | x2) & (~x0 | ((x4 | ~x5 | x7 | ~x1 | x2) & (x1 | ~x4 | (x2 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n1433 = ~x3 & ((~x5 & ~n1434) | (n487 & n531 & n727));
  assign n1434 = x0 ? ((x1 | x2 | x4 | ~x6 | ~x7) & (~x1 | ~x2 | ~x4 | x6 | x7)) : (x2 | ~x7 | (x1 ? (~x4 | ~x6) : (x4 | x6)));
  assign n1435 = (~x2 | n1437) & (n1071 | ((~x3 | n1436) & (x2 | x3 | ~x5)));
  assign n1436 = x2 ? (x5 | x6) : (~x5 | ~x6);
  assign n1437 = (~x0 & ~x3 & x5 & x6 & (x1 | x4)) | (~x5 & ((~x1 & ~x4) | (x0 & x3))) | (x1 & x4) | (~x4 & ((x0 & (~x1 | x3)) | (~x1 & (x3 | ~x6))));
  assign z094 = ~n1440 | (x0 & ((n269 & n1251) | (~x7 & ~n1439)));
  assign n1439 = x1 ? ((x4 | ~x5 | ~x6 | x2 | ~x3) & (~x4 | x5 | x6 | ~x2 | x3)) : (~x6 | ((~x2 | ~x3 | ~x4 | x5) & (x2 | (x3 ? (~x4 | ~x5) : (x4 | x5)))));
  assign n1440 = ~n1448 & ~n1447 & n1445 & ~n1443 & ~n1441 & ~n1442;
  assign n1441 = x2 & ((~x1 & ((~x5 & x6 & ~x0 & ~x3) | (x0 & (x3 ? (~x5 & ~x6) : (x5 & x6))))) | (~x0 & x5 & (~x3 ^ x6)));
  assign n1442 = ~x2 & (x5 ? ((x0 & x3 & ~x6) | (~x0 & ~x1 & ~x3 & x6)) : (((~x0 ^ ~x1) & (~x3 ^ x6)) | (~x0 & ~x1 & x3 & ~x6) | (x0 & x1 & ~x3 & x6)));
  assign n1443 = ~n1444 & ~x4 & n783;
  assign n1444 = (~x2 | x3 | x5 | x6 | ~x7) & (x2 | ((x6 | ~x7 | x3 | ~x5) & (~x3 | x5 | ~x6 | x7)));
  assign n1445 = (~x0 | x3 | x6 | ~x7 | n778) & (x0 | ((x7 | n778 | x3 | ~x6) & (~x3 | x6 | (n1446 & (~x7 | n778)))));
  assign n1446 = (~x2 | (x1 ? (~x4 | x5) : (x4 | ~x5))) & (~x1 | x2 | (x4 ^ x5));
  assign n1447 = ~n520 & ((~x0 & ~x1 & ~x2 & x4 & ~x5) | (x0 & ((~x4 & x5 & ~x1 & x2) | (x1 & ~x2 & (~x4 ^ x5)))));
  assign n1448 = n1215 & (x0 ? ((~x1 & ~x2 & x4 & ~x5) | (x1 & x2 & ~x4 & x5)) : (x1 & (x2 ? (~x4 ^ x5) : (~x4 & x5))));
  assign z095 = ~n1456 | (x1 ? ~n1450 : (x5 ? ~n1455 : ~n1454));
  assign n1450 = n1453 & (x0 ? (x2 | n1452) : n1451);
  assign n1451 = (~x4 | (x2 ? ((~x6 | ~x7 | x3 | x5) & (x6 | x7 | ~x3 | ~x5)) : ((~x5 | x6 | ~x7) & (~x6 | x7 | x3 | x5)))) & (x2 | x4 | ((~x3 | x5 | ~x6) & (x6 | x7 | x3 | ~x5)));
  assign n1452 = (~x3 | ~x4 | x5 | ~x6 | ~x7) & (x3 | ((x4 | x5 | ~x6) & (~x4 | ~x5 | x6 | ~x7)));
  assign n1453 = (~x4 | x6 | ~x7 | x0 | ~x2 | ~x3) & ((x0 ^ ~x3) | ((x6 | x7 | x2 | ~x4) & (~x6 | ~x7 | ~x2 | x4)));
  assign n1454 = (~x7 | ((x0 | x2 | x3 | ~x4 | x6) & (x4 | ~x6 | ((x0 | (~x2 & x3)) & (~x2 | x3) & (~x0 | x2 | ~x3))))) & (~x6 | x7 | (x0 ? ((x3 | x4) & (~x2 | ~x3 | ~x4)) : (~x3 | x4)));
  assign n1455 = x4 ? (x6 | (x0 ? ((~x3 | ~x7) & (~x2 | x3 | x7)) : ((~x2 | ~x3 | x7) & (x3 | (x2 & ~x7))))) : (((~x3 ^ x6) | (x0 ? (~x2 | x7) : (x2 | ~x7))) & (~x3 | ~x6 | x7 | x0 | ~x2) & (~x0 | x2 | x3 | x6 | ~x7));
  assign n1456 = (n950 | n1457) & (n467 | n1458);
  assign n1457 = ((~x3 ^ x6) | ((x0 | ~x1 | ~x2 | x7) & (~x0 | ((x2 | ~x7) & (x1 | (x2 & ~x7)))))) & ((x2 ? (x3 | x6) : (~x3 | ~x6)) | (x0 ? (~x1 | x7) : ~x7)) & (x0 | ((x6 | ~x7 | ~x1 | x3) & (x1 | (x3 ? (~x6 | (x2 & ~x7)) : (x6 | x7)))));
  assign n1458 = (~x1 | (x0 ? (x2 | ~x3) : x3)) & (x3 | x7 | x0 | ~x2) & (x1 | ((~x0 | (~x3 ^ x7)) & (~x3 | ~x7 | (x0 & ~x2))));
  assign z096 = n1460 | n1464 | ~n1465 | n1469 | (~x0 & ~n1468);
  assign n1460 = x1 & ((n1461 & n786) | n1463 | (x4 & ~n1462));
  assign n1461 = ~x3 & ~x0 & ~x2;
  assign n1462 = (x5 | ~x6 | ~x7 | ~x0 | x2 | ~x3) & (x0 | x3 | ((x2 | ~x5 | (x6 ^ x7)) & (~x6 | ~x7 | ~x2 | x5)));
  assign n1463 = ~n750 & ~n777 & (x4 ? (~x6 & ~x7) : (~x6 ^ ~x7));
  assign n1464 = ~n705 & ((~x2 & ~x5 & x7) | (x5 & ~x7 & ((x0 & ~x2 & x3) | (x2 & (~x0 | ~x3)))));
  assign n1465 = ~n1467 & ~n1466 & (x3 | x4 | x7 | ~n460);
  assign n1466 = x2 & x3 & ((x0 & ~x1 & (x4 ^ x7)) | (x4 & x7 & ~x0 & x1));
  assign n1467 = ~n440 & (x2 ? (~x3 & ((~x1 & ~x4) | (~x0 & x1 & x4))) : ((x1 & x3 & x4) | (x0 & (x1 ? x4 : (x3 & ~x4)))));
  assign n1468 = (x3 | ((x1 | x2 | x4 | ~x5 | x7) & (~x1 | x5 | (x2 ? (x4 | ~x7) : (~x4 | x7))))) & (x1 | ~x3 | x4 | (x2 ? (~x5 | ~x7) : (x5 | x7)));
  assign n1469 = ~x1 & (x6 ? ~n1470 : (~n750 & ~n700));
  assign n1470 = ((~x4 ^ x7) | (x0 ^ ~x3) | (x2 ^ ~x5)) & (~x0 | ~x2 | ~x3 | ~x4 | ~x5 | ~x7) & (x0 | x2 | x3 | x4 | x5 | x7);
  assign z097 = n1472 | ~n1476 | (n542 & ~n1475) | (~x2 & ~n1474);
  assign n1472 = ~n798 & ~n1473;
  assign n1473 = x0 ? (x4 | ((x2 | x5 | x7) & (x1 | (x2 ? (~x5 ^ x7) : (~x5 | ~x7))))) : ((~x4 | ~x7 | ((x1 | x2 | ~x5) & (~x2 | x5))) & (x7 | ((~x4 | ~x5 | x1 | ~x2) & (~x1 | (x2 ? (x4 | ~x5) : (~x4 | x5))))));
  assign n1474 = (x6 | ((~x0 | ((x4 | x5 | x1 | x3) & (~x1 | ~x3 | ~x4 | ~x5))) & (x5 | ((~x1 | x3 | ~x4) & (x0 | ~x3 | (x1 ^ ~x4)))))) & (x3 | ~x6 | ((~x1 | ~x4 | ~x5) & (x0 | x1 | x4 | x5)));
  assign n1475 = (~x5 | ((x0 | x3 | x4 | ~x6 | ~x7) & (~x4 | ((~x0 | (x3 ? (~x6 | x7) : (x6 | ~x7))) & (x6 | ~x7 | x0 | ~x3))))) & (~x0 | ~x3 | ~x4 | x5 | ~x6 | ~x7);
  assign n1476 = n1480 & ((x0 & (x1 | (x4 & n1477))) | (~x0 & ~x1 & ~x4 & n1477) | (n1263 & (x1 | n1477)));
  assign n1477 = (~x2 | n1478) & (x0 | x2 | x4 | n1479);
  assign n1478 = (~x0 | ~x3 | ~x4 | ~x5 | ~x6 | ~x7) & (x0 | x3 | x4 | x5 | x6 | x7);
  assign n1479 = (~x3 | x5 | ~x6 | x7) & (x3 | x6 | (x5 ^ ~x7));
  assign n1480 = n1482 & ((x2 & n1085) | n1481 | (~x2 & n416));
  assign n1481 = (x0 | x1 | ~x3 | x4) & (~x0 | x3 | (x1 ^ ~x4));
  assign n1482 = (x2 | (x1 ^ ~x4) | (x0 ? (~x3 | ~x5) : (x3 | x5))) & (x1 | ~x2 | ((x4 | ~x5 | x0 | x3) & (~x4 | x5 | ~x0 | ~x3)));
  assign z098 = ~n1490 | (x0 ? ~n1484 : (x4 ? ~n1489 : ~n1488));
  assign n1484 = (x1 | ((~x2 | n1486) & (~x5 | n1485))) & (x5 | n1487) & (~x1 | x2 | n1486);
  assign n1485 = (~x2 | ((x6 | ~x7 | ~x3 | x4) & (~x6 | x7 | x3 | ~x4))) & (x3 | x4 | ((~x6 | ~x7) & (x2 | x6 | x7)));
  assign n1486 = x3 ? (~x4 | ~x5 | (x6 ^ x7)) : (x4 | ((x6 | x7) & (x5 | ~x6 | ~x7)));
  assign n1487 = x1 ? ((x2 | ~x3 | ~x4 | ~x6 | ~x7) & (~x2 | x3 | x4 | x6 | x7)) : (x2 | x3 | (x4 ? (x6 | x7) : (~x6 | ~x7)));
  assign n1488 = ((x3 ? (x5 | ~x6) : (~x5 | x6)) | (x1 ? (~x2 | x7) : (x2 | ~x7))) & (~x1 | ~x5 | ~x6 | ((x3 | ~x7) & (x2 | ~x3 | x7))) & (x1 | x5 | x6 | ((~x3 | x7) & (~x2 | x3 | ~x7)));
  assign n1489 = (x2 | ((x6 | x7 | x3 | ~x5) & (~x3 | ((x6 | ~x7 | ~x1 | ~x5) & (~x6 | x7 | x1 | x5))))) & (x3 | ((~x6 | ~x7 | ~x2 | x5) & ((x6 ^ x7) | (x1 ^ ~x5))));
  assign n1490 = ~n1493 & (n437 | n1491) & (x0 ? n1494 : n1492);
  assign n1491 = (~x3 | (x0 ? (x4 | ((x2 | x5) & (x1 | (x2 & x5)))) : ((~x1 | ((~x4 | x5) & (~x2 | x4 | ~x5))) & (~x4 | (x5 ? x1 : ~x2))))) & (x2 | x3 | ((~x0 | ~x1 | ~x4 | ~x5) & (x0 | x1 | x4 | x5)));
  assign n1492 = x3 ? (x1 ? ((x5 | ~x6 | x2 | x4) & (~x5 | x6 | ~x2 | ~x4)) : (x4 | ~x6 | (~x2 & ~x5))) : ((x6 | ((x1 | x2 | ~x4 | x5) & (~x1 | x4 | (x2 & x5)))) & (~x5 | ~x6 | ~x1 | ~x4));
  assign n1493 = ~n950 & ((x2 & ~x3 & ~x6 & n783) | (~x2 & n595 & (~x3 ^ ~x6)));
  assign n1494 = (~x1 | ~x2 | x3 | x4 | ~x6) & (x1 | ((x2 | x3 | x4 | x5 | x6) & (~x4 | (~x3 ^ x6) | (x2 & x5))));
  assign z099 = n1504 | ~n1505 | (x0 ? ~n1496 : ~n1500);
  assign n1496 = (n585 | n1498) & (x3 | n1497) & (x1 | ~x3 | n1499);
  assign n1497 = (x7 | ((~x1 | x2 | x4 | ~x5 | ~x6) & (~x2 | ((~x1 | x5 | (~x4 ^ x6)) & (x1 | ~x4 | ~x5 | x6))))) & (x5 | ~x7 | ((x1 | x2 | (~x4 ^ x6)) & (~x1 | ~x2 | x4 | x6)));
  assign n1498 = (~x1 | x2 | ~x3 | x5 | ~x7) & (x1 | x3 | (x2 ? (~x5 | ~x7) : (x5 | x7)));
  assign n1499 = (x2 | x4 | x5 | x6 | x7) & (~x2 | ~x5 | (x4 ? (x6 | x7) : (~x6 ^ x7)));
  assign n1500 = ~n1501 & n1502 & ((x7 & (x3 | x6)) | n853 | (~x6 & ~x7));
  assign n1501 = n370 & ((~x1 & ~x2 & x3 & ~x5 & ~x6) | (x1 & x6 & (x2 ? (x3 & ~x5) : (~x3 & x5))));
  assign n1502 = x6 ? ((~x7 | n1503) & (x1 | x2 | n1272)) : ((x7 | n1503) & (~x1 | ~x2 | n1272));
  assign n1503 = (x1 | ~x2 | x3 | ~x4 | x5) & (~x1 | x2 | ~x3 | x4 | ~x5);
  assign n1504 = ~n699 & (x0 ? ((~x2 & (x1 ? (~x3 & ~x5) : x5)) | (~x1 & ~x5 & (x2 | x3))) : ((x1 & x2 & x5) | (~x3 & ~x5 & ~x1 & ~x2)));
  assign n1505 = n1508 & (x2 | n1506) & (n1507 | (x0 ? (~x2 | ~x5) : (x2 ^ ~x5)));
  assign n1506 = (x0 | x1 | x3 | ~x4 | ~x5 | ~x7) & (~x3 | x7 | (~x4 ^ x5) | (~x0 ^ ~x1));
  assign n1507 = (~x1 | x3 | x4 | x7) & (~x4 | ~x7 | x1 | ~x3);
  assign n1508 = n1509 & (~n400 | n700);
  assign n1509 = (~x4 | ~x5 | ~x7 | ~x0 | ~x1 | x2) & (x0 | (x4 ^ x7) | (x1 ? (x2 | x5) : (~x2 | ~x5)));
  assign z100 = n1511 | n1512 | ~n1515 | ~n1517 | (n837 & ~n1514);
  assign n1511 = x5 & (((x3 ^ x6) & (x0 ? (x1 & ~x2) : (~x1 ^ x2))) | (x3 & x6 & (x0 ? (~x1 & x2) : (x1 & ~x2))));
  assign n1512 = n1215 & ((n279 & ~n1513) | (~x2 & n654 & n349));
  assign n1513 = x1 ? (x4 | x5) : (~x4 | ~x5);
  assign n1514 = (~x3 | ~x6 | (~x5 ^ x7)) & (x3 | x4 | ~x5 | x6 | ~x7);
  assign n1515 = ((x0 ? (x1 | ~x2) : (~x1 | x2)) | (n1516 & (x5 | x6))) & (x1 | x5 | ~x6 | (x0 ^ ~x2));
  assign n1516 = (~x3 | ~x4 | ~x5 | x6 | ~x7) & (x3 | ~x6 | ((x5 | x7) & (x4 | ~x5 | ~x7)));
  assign n1517 = (x6 | n1518) & (n1519 | (x0 ^ ~x2));
  assign n1518 = ((x0 ^ ~x2) | ((x1 | (x3 ? (~x4 | x5) : (x4 | ~x5))) & (~x4 | ~x5 | ~x1 | x3))) & (x3 | ~x5 | ((x0 | x1 | x2 | ~x4) & (~x0 | ~x1 | ~x2 | x4)));
  assign n1519 = x1 ? (x3 ? (~x6 | ((x5 | ~x7) & (x4 | ~x5 | x7))) : (x4 | x6 | (x5 ^ x7))) : (x6 | ((~x5 | x7 | x3 | ~x4) & (~x3 | x4 | (~x5 ^ x7))));
  assign z101 = ~n1523 | ~n1528 | (x6 ? (x7 ? ~n1522 : ~n1521) : (x7 ? ~n1521 : ~n1522));
  assign n1521 = x0 ? ((~x1 | x2 | x3 | x4 | x5) & (x1 | ((~x4 | ~x5 | ~x2 | ~x3) & (x2 | (x3 ? (x4 | x5) : (~x4 | ~x5)))))) : (x1 ? ((x4 | x5 | ~x2 | x3) & (~x4 | ~x5 | x2 | ~x3)) : (x2 ? (x3 ? (x4 | x5) : (~x4 | ~x5)) : (x3 | x4)));
  assign n1522 = ((~x4 ^ x5) | (x0 ? (x1 ? (x2 | ~x3) : (~x2 | x3)) : (~x1 | (x2 ^ x3)))) & (x0 | x1 | x2 | ~x3 | (~x4 & ~x5));
  assign n1523 = ~n1525 & n1526 & ~n1527 & (n1524 | (n456 & n467));
  assign n1524 = x0 ? (x1 ? (x2 | ~x3) : (~x2 | x3)) : (~x1 | (x2 ^ x3));
  assign n1525 = (x2 ? (~x4 & x6) : (x4 & ~x6)) & (x0 ? (~x1 ^ ~x3) : (~x1 & ~x3));
  assign n1526 = x4 | ~n345 | ((~x0 | x3 | ~x6) & (x5 | x6 | x0 | ~x3));
  assign n1527 = ~x0 & ((x3 & x4 & ~x6 & ~x1 & x2) | (x1 & ((~x4 & x6 & ~x2 & x3) | (x4 & ~x6 & x2 & ~x3))));
  assign n1528 = x0 ? n1531 : (x1 ? n1529 : n1530);
  assign n1529 = (~x5 | x6 | ~x7 | ~x2 | x3 | x4) & (x5 | ~x6 | x7 | x2 | ~x3 | ~x4);
  assign n1530 = (x2 | ~x3 | x4 | x5 | ~x6 | ~x7) & (~x2 | ((x5 | ~x6 | x7 | x3 | ~x4) & (~x5 | x6 | ~x7 | ~x3 | x4)));
  assign n1531 = x1 ? (~n357 | ~n786) : n1532;
  assign n1532 = (~x2 | ~x3 | ~x4 | x5 | ~x6 | x7) & (x2 | ((x5 | ~x6 | x7 | x3 | ~x4) & (~x5 | x6 | ~x7 | ~x3 | x4)));
  assign z102 = n1535 | ~n1539 | (x7 & ~n1534) | (~n858 & ~n1538);
  assign n1534 = ((~x4 ^ x5) | (x0 ? (x1 ? (x2 | ~x3) : (~x2 | x3)) : (x1 ? (x2 ^ x3) : (x2 | ~x3)))) & (~x0 | ((~x1 | x2 | x3 | x4 | x5) & (x1 | ((~x4 | ~x5 | ~x2 | ~x3) & (x2 | (x3 ? (x4 | x5) : (~x4 | ~x5))))))) & (x0 | (x1 ? ((x4 | x5 | ~x2 | x3) & (~x4 | ~x5 | x2 | ~x3)) : ((x4 | x5 | x2 | x3) & (~x2 | (x3 ? (x4 | x5) : (~x4 | ~x5))))));
  assign n1535 = x5 & ((~n437 & ~n1537) | (x3 & n345 & ~n1536));
  assign n1536 = (x0 | ~x4 | x6 | ~x7) & (~x0 | x4 | ~x6 | x7);
  assign n1537 = (x0 | ~x2 | ~x3 | (~x1 ^ ~x4)) & (x3 | ((~x0 | (x1 ? (x2 | x4) : (~x2 | ~x4))) & (x0 | ~x1 | ~x2 | x4)));
  assign n1538 = (~x7 | ((x1 | ~x2 | ~x4 | x5 | ~x6) & (x2 | ((~x1 | (x4 ? (~x5 | x6) : (x5 | ~x6))) & (x1 | x4 | ~x5 | x6))))) & (~x1 | x2 | x7 | (x4 ? (~x5 | ~x6) : (x5 | x6)));
  assign n1539 = (x7 | n1540) & (x5 | (~n1541 & n1543));
  assign n1540 = x0 ? ((x3 | x4 | x1 | x2) & ((~x2 ^ x4) | (x1 ^ ~x3))) : (((x2 ? (x3 | ~x4) : (~x3 | x4)) | (~x1 & x5)) & (x1 | (x2 ? (x3 ^ x4) : (x3 | ~x4))));
  assign n1541 = ~n1542 & n279 & ~x7 & x4 & ~x6;
  assign n1542 = x1 ^ ~x3;
  assign n1543 = (~n373 | ~n374 | ~n317) & (n515 | n1544 | (~n372 & ~n374));
  assign n1544 = x0 ? (x1 | x3) : (~x1 | ~x3);
  assign z103 = n1547 | ~n1550 | ~n1553 | (n783 & ~n1546);
  assign n1546 = x3 ? ((~x2 | x4 | x5 | x6 | x7) & (x2 | ((~x6 | ~x7 | x4 | x5) & (~x4 | (x5 ? (~x6 | ~x7) : (x6 | x7)))))) : (x2 ? ((x6 | x7 | x4 | ~x5) & (~x6 | ~x7 | ~x4 | x5)) : (~x5 | (x4 ? (x6 | x7) : (~x6 | ~x7))));
  assign n1547 = n1548 & (x0 ? (x1 & n784) : (~x1 & n1549));
  assign n1548 = x2 & ~x4;
  assign n1549 = x6 & x3 & x5;
  assign n1550 = (x0 | (n1551 & (~x1 | ~x6 | n1552))) & (~x6 | n1551) & (~x0 | x1 | n1552);
  assign n1551 = (x1 | ~x2 | ~x3 | ~x4 | x5) & (~x1 | x2 | x3 | x4 | ~x5);
  assign n1552 = (~x2 | x3 | x4 | ~x5) & (x2 | ~x3 | ~x4 | x5);
  assign n1553 = x4 ? ((~x5 | n1555) & (x3 | x5 | n1554)) : ((x5 | n1555) & (~x3 | ~x5 | n1554));
  assign n1554 = (x0 & (x2 | (~x1 & ~x6))) | (~x0 & x1 & ~x2) | (~x1 & x2);
  assign n1555 = x1 ? ((x2 | ~x3 | ~x6) & (x0 | ((~x3 | ~x6) & (x2 | (~x3 & ~x6))))) : ((~x0 | (x2 ^ x3)) & (~x2 | x3 | (x0 & ~x6)));
  assign z104 = ~n1558 | n1563 | (~n416 & ~n1557) | (~x1 & ~n1562);
  assign n1557 = (x0 | ((~x1 | (x3 ? (x2 ? ~x4 : (x4 | x7)) : (~x4 | x7))) & ((~x2 ^ x4) | (x3 & (x1 | ~x7))) & (~x4 | x7 | ~x2 | ~x3) & (x4 | ~x7 | x1 | x3))) & (x3 | (x2 ? ((~x0 | x1 | ~x4) & (~x1 | x4 | x7)) : ((~x1 | ~x4 | x7) & (~x0 | x4 | (~x1 & x7))))) & (~x0 | ~x3 | ((x1 | x4 | (x2 & x7)) & (x2 | ~x4 | (~x1 & x7))));
  assign n1558 = (n420 | n1559) & (~x1 | (n1560 & (x7 | n1561)));
  assign n1559 = (x1 | ((~x2 | (x0 ? ~x3 : (x3 | ~x7))) & (~x0 | x3 | (x2 & x7)))) & (~x1 | x2 | ~x3 | x7) & (x0 | ((x2 | ~x3) & (~x1 | x7 | (x2 & ~x3))));
  assign n1560 = ((x0 ^ ~x2) | ((~x5 | x6 | x3 | ~x4) & (x5 | ~x6 | ~x3 | x4))) & (x3 | x4 | ((x0 | x2 | x5 | ~x6) & (~x0 | ~x2 | ~x5 | x6)));
  assign n1561 = (x4 | x5 | ~x6 | ~x0 | x2 | x3) & (x0 | ((x4 | x5 | ~x6 | ~x2 | x3) & (~x4 | ~x5 | x6 | x2 | ~x3)));
  assign n1562 = x0 ? ((x4 | x5 | ~x6 | ~x2 | x3) & (~x4 | ~x5 | x6 | x2 | ~x3)) : ((x4 | x5 | ~x6 | x2 | x3) & (~x2 | ((~x4 | ~x5 | x6) & (x5 | ~x6 | ~x3 | x4))));
  assign n1563 = ~x1 & ((x3 & ~n1564) | (n1565 & (~x0 ^ ~x7)));
  assign n1564 = (x0 | x2 | x4 | x5 | ~x6 | ~x7) & (x7 | ((x0 | ~x2 | x4 | ~x5 | ~x6) & (~x0 | ((~x2 | ~x4 | ~x5 | x6) & (x2 | x4 | x5 | ~x6)))));
  assign n1565 = ~x6 & x5 & x4 & ~x2 & ~x3;
  assign z105 = n1567 | ~n1568 | (x3 ? ~n1573 : (n1571 | n1572));
  assign n1567 = ~n434 & (x1 ? ((~x2 & x3 & ~x4) | (~x0 & ((x3 & ~x4) | (x2 & ~x3 & x4) | (~x2 & (x3 | ~x4))))) : ((x2 & (~x3 ^ x4)) | (~x3 & (x4 ? ~x2 : x0))));
  assign n1568 = x6 ? ((~x7 | n1569) & (~x3 | ~x5 | x7 | n1570)) : ((x7 | n1569) & (x3 | x5 | ~x7 | n1570));
  assign n1569 = (x0 | ((~x2 | ((~x3 | ~x4 | ~x5) & (~x1 | x4 | x5))) & (~x1 | ((~x4 | (~x3 ^ x5)) & (x2 | ((~x4 | x5) & (~x3 | x4 | ~x5))))))) & (x1 | ((~x2 | (x3 ? (x4 | ~x5) : (~x4 | x5))) & (~x4 | x5 | ~x0 | x3) & (x2 | (x3 ? (x4 ^ x5) : (x4 | ~x5))))) & (~x1 | ((x4 | ~x5 | ~x2 | x3) & (x2 | (x3 ? (~x4 | x5) : (x4 ^ x5)))));
  assign n1570 = x1 ? (x2 ? x0 : ~x4) : (x2 | x4);
  assign n1571 = ~x7 & n531 & (x1 ? ((~x2 & ~x4) | (~x0 & (~x2 | ~x4))) : (x4 & (x0 | x2)));
  assign n1572 = n269 & n524;
  assign n1573 = (~n686 | ~n511) & (~x7 | ~n312 | n1574);
  assign n1574 = (x1 | (~x2 ^ x4)) & (x0 | ((~x2 | ~x4) & (~x1 | x2 | x4)));
  assign z106 = n1576 | n1579 | n1580 | n1581 | (~n425 & ~n1578);
  assign n1576 = ~x5 & ((x0 & ~n1577) | (~x4 & n292 & n278));
  assign n1577 = (x1 | ~x3 | ((x4 | x6 | ~x7) & (~x6 | x7 | ~x2 | ~x4))) & (x3 | x6 | ((~x1 | ~x2 | ~x4 | x7) & (x2 | x4 | ~x7)));
  assign n1578 = ((x4 ^ x5) | (x2 ? (x3 | (x0 & x1)) : (~x3 | (~x0 & ~x1)))) & (x1 | ((~x4 | ~x5 | x0 | ~x2) & (~x0 | ((~x2 | ~x4 | x5) & (~x3 | x4 | ~x5))))) & (~x3 | ~x4 | x5 | x0 | ~x2) & (x2 | ((x3 | x4 | ~x5) & (x0 | ((x4 | ~x5) & (x3 | ~x4 | x5)))));
  assign n1579 = n996 & (x0 ? (~x1 & x2) : (~x2 ^ x3));
  assign n1580 = (~x0 | ((x2 | x4) & (~x1 | ~x3))) & (x0 | x3 | (~x2 & (x1 | ~x4))) & (~x2 | ~x4) & ~n434 & (x2 | ~x3 | x4);
  assign n1581 = ~n1020 & (x2 ? ((~x1 & ~x3) | (~x0 & (~x1 | ~x3))) : (x3 & (x0 | x1)));
  assign z107 = ~n1590 | (x4 ? ~n1588 : (~n1584 | (x1 & ~n1583)));
  assign n1583 = (~x5 | ~x6 | x7 | ~x0 | x2 | x3) & (x6 | ((~x0 | ~x2 | x3 | x5 | ~x7) & (~x3 | ((x0 | ~x2 | ~x5 | ~x7) & (x2 | (x0 ? (x5 ^ x7) : (x5 | ~x7)))))));
  assign n1584 = ~n1587 & (~n459 | ~n1586) & (x5 | ~n543 | ~n1585);
  assign n1585 = ~x3 & ~x0 & x1;
  assign n1586 = ~x7 & ~x6 & ~x3 & x5;
  assign n1587 = ~x1 & (x3 ? (~x6 & x7) : (x6 & ~x7)) & (x0 ^ ~x5);
  assign n1588 = (x0 | n1589) & (~x0 | ~n292 | ~n354 | ~n784);
  assign n1589 = (x6 | ~x7 | ~x3 | ~x5) & (x7 | ((~x1 | ((x3 | ~x5 | ~x6) & (~x2 | ~x3 | x5 | x6))) & (x3 | ~x6 | ((~x2 | ~x5) & (x1 | x2 | x5)))));
  assign n1590 = (n437 | n1594) & (n425 | n1593) & (n1591 | n1592);
  assign n1591 = x3 ? (~x6 | x7) : (x6 | ~x7);
  assign n1592 = x0 ? ((x4 | x5 | x1 | ~x2) & (x2 | (x1 ? (x4 ^ x5) : (~x4 | x5)))) : (x1 ? (~x4 | x5) : (x4 | ~x5));
  assign n1593 = x3 ? ((~x0 | ~x4 | (x1 & x2) | x5) & (x0 | x4 | ~x5) & (x1 | ((x2 | x4 | ~x5) & (x0 | (~x5 & (x2 | x4)))))) : ((~x0 | ((x1 | (x4 ^ x5)) & (~x5 | (x4 ? x2 : ~x1)))) & (x4 | x5 | ~x1 | x2) & (x0 | ((~x4 | x5) & (~x1 | (x5 & (~x2 | ~x4))))));
  assign n1594 = x1 ? ((x3 | ~x4 | x5 | ~x0 | x2) & (x0 | x4 | ((x3 | ~x5) & (~x2 | ~x3 | x5)))) : ((x0 | x2 | x3 | ~x4 | ~x5) & (~x3 | (x0 ? ((~x4 | ~x5) & (x2 | x4 | x5)) : (~x4 | x5))));
  assign z108 = n1596 | ~n1598 | (~n665 & ~n1605) | (x0 & ~n1606);
  assign n1596 = x1 & ((n1029 & n1197) | (x4 & ~n1597));
  assign n1597 = (~x2 | x3 | x5 | x6 | x7) & (x2 | (x6 ^ x7) | (x0 ? (~x3 | x5) : (x3 | ~x5)));
  assign n1598 = ~n1603 & (x0 | n1604) & (x1 | (~n1599 & ~n1601));
  assign n1599 = ~n559 & (x0 ? (x7 & ~n447) : (x3 & n1600));
  assign n1600 = ~x7 & ~x4 & x6;
  assign n1601 = ~x7 & n312 & n1602 & (~x2 ^ ~x3);
  assign n1602 = ~x0 & ~x4;
  assign n1603 = ~n434 & (((~x2 | ~x3) & ((x1 & ~x4) | (x0 & ~x1 & x4))) | (~x1 & ~x2 & ~x3 & x4) | (~x0 & x2 & (x1 ^ ~x4)));
  assign n1604 = x1 ? ((x2 | ~x4 | x5 | x6 | x7) & (~x2 | x4 | ~x5 | ~x6 | ~x7)) : (~x4 | ((~x5 | ~x6 | ~x7) & (x6 | x7 | ~x2 | x5)));
  assign n1605 = (x1 | (x4 ? (x6 | (x0 & ~x2)) : ((~x0 | (x6 ? ~x3 : x2)) & (~x6 | (x3 ? x2 : (x0 & ~x2)))))) & (x0 | ~x2 | ~x3 | ~x4 | ~x6) & (~x1 | (x0 ? (x2 | (~x4 ^ x6)) : (x4 ? ~x6 : (x6 | (~x2 & ~x3)))));
  assign n1606 = (x1 | x4 | x5 | x6 | x7) & (~x5 | ~x6 | ~x7 | (x1 ? (x2 | ~x4) : (x2 ^ x4)));
  assign z109 = ~n1613 | (x2 ? ~n1608 : (x5 ? ~n1611 : ~n1612));
  assign n1608 = (~x6 | n1609) & (x0 | x6 | n1610);
  assign n1609 = (x4 | ((x1 | (x0 ? (x3 ? (x5 | x7) : (~x5 | ~x7)) : (~x5 | x7))) & (x0 | x7 | ((~x3 | ~x5) & (~x1 | x3 | x5))))) & (x0 | ~x4 | ((~x1 | ((~x5 | x7) & (~x3 | x5 | ~x7))) & (x3 | ((~x5 | x7) & (x1 | x5 | ~x7)))));
  assign n1610 = (~x3 | ((x4 | x5 | ~x7) & (~x1 | ((x5 | ~x7) & (~x4 | ~x5 | x7))))) & (x1 | x3 | ((x5 | ~x7) & (x4 | ~x5 | x7)));
  assign n1611 = (~x6 | ((x0 | ~x1 | ~x3 | x4 | ~x7) & (x7 | ((x0 | x1 | ~x3 | ~x4) & (~x0 | (~x1 & (x3 | x4))))))) & (~x1 | x3 | ((~x0 | ~x4 | x7) & (x6 | ~x7 | x0 | x4)));
  assign n1612 = (x6 | ~x7 | ~x0 | x3) & (~x1 | ((x0 | ~x3 | x4 | x6 | x7) & (~x0 | ~x7 | (x6 & (~x3 | x4)))));
  assign n1613 = (~x6 | (x7 ? n1614 : n1615)) & (n434 | n1616) & (x6 | (x7 ? n1615 : n1614));
  assign n1614 = x0 ? ((~x1 | x3 | (x2 ? (x4 | ~x5) : x5)) & (x2 | ~x3 | ~x5) & (x1 | (x2 ? (x5 | (~x3 & ~x4)) : ~x5))) : (x5 ? (x1 ? (x2 | x3) : (~x2 | (~x3 & ~x4))) : (x2 ? ((~x1 | (x3 & x4)) & (x3 | x4)) : ((~x3 | ~x4) & (x1 | (~x3 & ~x4)))));
  assign n1615 = x1 ? (x3 | x4 | (x0 ? (~x2 | x5) : (~x2 ^ ~x5))) : (~x3 | (x0 ? (x2 ? ~x5 : (x4 | x5)) : (x2 ? (~x4 | x5) : (x4 | ~x5))));
  assign n1616 = (x1 | (x0 ? (x2 ? x3 : (~x3 | ~x4)) : (x2 | x3))) & (x0 | x2 | (x3 ? ~x1 : ~x4));
  assign z110 = ~n1618 | ~n1627 | (~x3 & (n1622 | n1624 | ~n1625));
  assign n1618 = n1621 & (x2 ? (x0 | n1620) : n1619);
  assign n1619 = x0 ? ((x1 | x3 | ~x4 | ~x5 | x6) & (~x1 | ~x3 | x4 | x5 | ~x6)) : ((~x4 | x5 | x6 | x1 | ~x3) & (x3 | ((x5 | ~x6 | x1 | x4) & (~x1 | (x4 ? (~x5 | ~x6) : (x5 | x6))))));
  assign n1620 = (x1 | ~x3 | ~x4 | ~x5 | x6) & (x3 | (~x4 ^ x5) | (~x1 ^ x6));
  assign n1621 = x1 ? (x0 ? (x3 | (x2 ? (x4 | x6) : (~x4 | ~x6))) : (~x3 | ~x6 | (x2 ^ x4))) : ((x4 | x6 | x2 | ~x3) & (~x0 | ~x2 | (x3 ? (~x4 | x6) : (x4 | ~x6))));
  assign n1622 = ~n1623 & (~x0 ^ ~x5);
  assign n1623 = (x1 | ~x2 | ~x4 | ~x6 | x7) & (~x1 | ((~x4 | x6 | x7) & (x2 | ((x6 | x7) & (x4 | ~x6 | ~x7)))));
  assign n1624 = ~n425 & ((x0 & x1 & ~x2 & ~x4 & x5) | (~x0 & ~x5 & (x1 ? (~x2 & x4) : (x2 & ~x4))));
  assign n1625 = (~n992 | ~n697) & (x4 | ~n321 | ~n1626);
  assign n1626 = ~x5 & ~x7 & (~x2 ^ ~x6);
  assign n1627 = (n437 | n1628) & (~x3 | (~n1629 & (x1 | ~n1631)));
  assign n1628 = (~x5 | ((~x0 | ((~x1 | x2 | ~x3) & (x3 | ~x4 | x1 | ~x2))) & (x1 | x2 | x3 | (x0 & x4)))) & (~x2 | x4 | ((x1 | ~x3 | x5) & (x0 | (x1 ? (x3 | x5) : ~x3)))) & (x2 | ~x4 | (x1 ? ~x3 : (x3 | x5)));
  assign n1629 = ~n425 & (~n1630 | (~x2 & n654 & n783));
  assign n1630 = (~x0 | x1 | x2 | ~x4) & (x0 | ~x1 | ~x2 | x4);
  assign n1631 = x7 & (~x2 ^ ~x6) & (x0 ? (~x4 & x5) : (x4 & ~x5));
  assign z111 = (x3 & ~n1633) | (~x3 & ~n1636) | ~n1641 | (~x7 & ~n1640);
  assign n1633 = (~x5 | n1635) & (~x4 | x5 | ~n783 | n1634);
  assign n1634 = x2 ? (x6 | x7) : (x6 ^ ~x7);
  assign n1635 = (x4 | ~x6 | ~x7 | x0 | ~x1 | ~x2) & (~x0 | ((x2 | ((~x1 | ~x6 | (x4 ^ x7)) & (x6 | ~x7 | x1 | x4))) & (x1 | ~x2 | x4 | (x6 ^ x7))));
  assign n1636 = (x0 | ~x5 | n1639) & (x5 | ((~n1637 | ~n992) & (~x0 | n1638)));
  assign n1637 = x7 & ~x4 & x6;
  assign n1638 = (x1 | ~x2 | x6 | (x4 ^ x7)) & (x2 | (x1 ? (~x4 | (x6 ^ x7)) : (x4 | (~x6 ^ x7))));
  assign n1639 = x1 ? (~x4 | (x2 ? (~x6 | x7) : (x6 ^ x7))) : ((x2 | x4 | ~x6 | x7) & (~x2 | ~x4 | x6 | ~x7));
  assign n1640 = (x2 | ((x0 | x1 | ~x3 | ~x4 | ~x5) & (x3 | (~x4 ^ x5) | (x0 ^ ~x1)))) & (~x0 | x1 | ~x2 | (x3 ? (x4 | x5) : (~x4 | ~x5)));
  assign n1641 = ~n1646 & ~n1645 & ~n1644 & ~n1642 & ~n1643;
  assign n1642 = x7 & ((~x2 & ((~x4 & ~x5 & ~x0 & ~x3) | (x0 & (x3 ? (~x4 & ~x5) : (x4 & x5))))) | (~x0 & x2 & ~x3 & (x4 ^ x5)));
  assign n1643 = ~x0 & ((x3 & ~x4 & (x2 ^ x7)) | (~x1 & x4 & (x2 ? (x3 & x7) : (~x3 & ~x7))));
  assign n1644 = (x2 ^ ~x7) & ((x3 & x4 & ~x0 & x1) | (x0 & (x1 ? (~x3 & ~x4) : (x3 & x4))));
  assign n1645 = x0 & ((~x3 & ~x4 & x7 & ~x1 & x2) | (x3 & x4 & ~x7 & x1 & ~x2));
  assign n1646 = ~x7 & ~x5 & ~x4 & ~x3 & ~x0 & x2;
  assign z112 = ~n1651 | ~n1658 | n1659 | (x1 ? ~n1648 : ~n1660);
  assign n1648 = x6 ? (~n1602 | n1650) : n1649;
  assign n1649 = (x0 | ~x3 | ~x4 | ~x5 | ~x7) & (x3 | (x0 ? ((~x5 | ~x7 | x2 | x4) & (x5 | x7 | ~x2 | ~x4)) : (~x4 | (x2 ? (~x5 | x7) : (x5 | ~x7)))));
  assign n1650 = (x2 | ~x3 | x5 | ~x7) & (~x2 | x7 | (x3 ^ x5));
  assign n1651 = n1656 & (n585 | n1655) & (x1 | (~n1652 & n1653));
  assign n1652 = x6 & n545 & ((n870 & n1230) | (n748 & n664));
  assign n1653 = (~n1461 | ~n464) & (n1654 | (x3 ? (x5 | x6) : (~x5 | ~x6)));
  assign n1654 = (~x0 | x2 | x4 | ~x7) & (x0 | ~x2 | ~x4 | x7);
  assign n1655 = x0 ? (x7 | ((~x3 | ~x5 | ~x1 | x2) & (x3 | x5 | x1 | ~x2))) : (x1 | x2 | ~x7 | (x3 ^ x5));
  assign n1656 = (x0 | ~x1 | n1657) & (n1079 | ((x0 | x1 | x2 | ~x3) & (~x0 | x3 | (x1 ^ ~x2))));
  assign n1657 = (~x2 | x3 | x4 | x5 | x6) & (~x3 | ~x4 | ~x5 | ~x6);
  assign n1658 = x1 ? ((x4 | (x0 ? (x2 ? (x3 | ~x5) : (~x3 | x5)) : (x2 | (x3 ^ x5)))) & (x3 | ~x4 | x5 | x0 | ~x2)) : (((x2 ? (~x3 | x4) : (x3 | ~x4)) | (x0 ^ ~x5)) & (x0 | ~x2 | x3 | x4 | x5) & (~x4 | ~x5 | ~x0 | ~x3));
  assign n1659 = ~n1085 & ((~x2 & ((~x0 & x1 & ~x3 & x4) | (x0 & x3 & (x1 ^ ~x4)))) | (~x0 & x2 & (x1 ? (x3 & ~x4) : (~x3 & x4))));
  assign n1660 = (x0 | ~x2 | ~x3 | ~x4 | ~x5 | ~x6) & (x4 | ((x0 | x2 | x3 | x5 | ~x6) & (~x0 | x6 | (x2 ? (~x3 | ~x5) : (x3 | x5)))));
  assign z113 = n1662 | ~n1666 | (x3 ? ~n1664 : ~n1665);
  assign n1662 = ~x0 & ((x1 & n509 & n284) | (~x5 & ~n1663));
  assign n1663 = (~x6 | ((~x1 | x3 | ~x4 | (x2 ^ ~x7)) & (x1 | ~x2 | ~x3 | x4 | x7))) & (x4 | x6 | ~x7 | ~x1 | x2 | ~x3);
  assign n1664 = x0 ? (x1 | ((x2 | (x4 ? ~x6 : (x6 | x7))) & (~x4 | ((~x6 | x7) & (~x2 | x6 | ~x7))))) : ((x4 | ~x6 | x7 | ~x1 | x2) & (~x2 | ((x6 | x7 | x1 | ~x4) & (~x7 | (x1 ? (x4 ^ x6) : (x4 | ~x6))))));
  assign n1665 = x0 ? ((~x7 | ((~x4 | ~x6 | x1 | x2) & (~x1 | (x2 ? (x4 | ~x6) : (~x4 | x6))))) & (x1 | ((~x6 | x7 | ~x2 | ~x4) & (x4 | x6 | (x2 & x7))))) : ((~x1 | x2 | x4 | ~x6 | ~x7) & (~x4 | x6 | x7 | x1 | ~x2) & ((~x6 ^ x7) | (x1 ? (~x2 | x4) : (x2 | ~x4))));
  assign n1666 = ~n1667 & ~n1670 & (x4 ? (x5 ? n1669 : n1668) : (x5 ? n1668 : n1669));
  assign n1667 = ~n589 & ((~x0 & ~x1 & x2 & ~x3 & x7) | (~x2 & ((x3 & x7 & x0 & x1) | (~x0 & (x1 ? (~x3 & ~x7) : (x3 & x7))))));
  assign n1668 = x0 ? ((x6 | x7 | ~x1 | x2) & (x1 | ((~x6 | x7 | x2 | x3) & (x6 | (x2 ? (~x3 ^ x7) : (~x3 | ~x7)))))) : ((x1 | x2 | x6 | x7) & (~x1 | ~x6 | (x2 ? (~x3 ^ x7) : (~x3 | ~x7))));
  assign n1669 = (~x6 | ((x2 | (~x0 ^ ~x1) | (~x3 ^ x7)) & (x1 | ~x2 | (x0 ? ~x7 : (x3 | x7))))) & (x0 | x6 | ((~x3 | ~x7 | x1 | ~x2) & (~x1 | (x2 ? x7 : (x3 | ~x7)))));
  assign n1670 = x0 & ((~x4 & ~n1672) | (x4 & ~x7 & n1671 & ~n1436));
  assign n1671 = x1 & ~x3;
  assign n1672 = (x1 | ~x3 | ~x5 | (x2 ? (x6 | ~x7) : (~x6 | x7))) & (x5 | ~x6 | x7 | ~x1 | ~x2 | x3);
  assign z114 = ~n1675 | n1681 | ~n1683 | (~n665 & ~n1674);
  assign n1674 = x0 ? ((~x1 | ~x2 | x3 | x4 | ~x6) & (x2 | ((~x1 | (~x3 & x6)) & (~x6 | (x3 ? x4 : x1))))) : (((x1 ^ x2) | ((~x3 | ~x4) & x6)) & (x1 | ~x2 | (x3 & x4) | ~x6));
  assign n1675 = n1677 & ~n1680 & (n425 | n1676) & (x3 | n1679);
  assign n1676 = (x0 | ~x1 | x2 | x3 | x4 | x5) & (~x3 | ((x1 | ((~x4 | x5 | x0 | ~x2) & (~x0 | (x2 ? ~x5 : (~x4 | x5))))) & (x0 | ~x1 | x2 | ~x5)));
  assign n1677 = (~n283 | ~n1292) & (n1678 | (x2 ? (~x6 | x7) : (x6 | ~x7)));
  assign n1678 = (~x0 | x1 | x3 | x5) & (x0 | ~x1 | ~x5 | (~x3 ^ x4));
  assign n1679 = (x0 | ~x1 | x2 | (x4 ? (x5 | x7) : (~x5 | ~x7))) & (~x0 | x1 | ~x2 | ~x5 | ~x7);
  assign n1680 = n1671 & ((x2 & ~n667) | (x0 & ~x2 & n531));
  assign n1681 = x3 & ((~x1 & ~n1682) | (n351 & n543 & n283));
  assign n1682 = (x7 | ((x0 | x2 | x4 | ~x5 | ~x6) & (x5 | (x0 ^ ~x2) | (x4 ^ x6)))) & (~x5 | x6 | ~x7 | ~x0 | ~x2 | x4);
  assign n1683 = x1 ? (x3 | n1685) : (n1684 & (x3 | ~x4 | n1686));
  assign n1684 = x0 ? ((x6 | x7 | x3 | x5) & (~x3 | ((x6 | ~x7 | x2 | ~x5) & (~x6 | x7 | ~x2 | x5)))) : ((x2 | x3 | x5 | ~x6 | x7) & (~x7 | ((~x5 | ~x6 | x2 | x3) & (~x2 | x6 | (x3 ^ x5)))));
  assign n1685 = (x5 | x6 | ~x7 | ~x0 | ~x2 | x4) & (~x6 | ((x2 | x4 | x5 | x7) & (x0 | ((~x5 | ~x7 | x2 | ~x4) & (x4 | x5 | x7)))));
  assign n1686 = (~x0 | x2 | ~x5 | x6 | ~x7) & (x0 | x7 | (x2 ? (x5 | x6) : (~x5 | ~x6)));
  assign z115 = ~n1694 | (x5 ? ~n1690 : (x0 ? ~n1688 : ~n1689));
  assign n1688 = (x6 | x7 | ((x1 | ~x2 | x3 | x4) & (x2 | (x1 ? (~x3 ^ x4) : (~x3 | ~x4))))) & (~x4 | ~x6 | ~x7 | (x1 ? (x2 | x3) : ~x3));
  assign n1689 = (~x6 | ~x7 | ((~x1 | ~x2 | ~x3 | x4) & ((x1 ^ ~x3) | (~x2 ^ ~x4)))) & (x4 | x6 | x7 | ((x2 | ~x3) & (~x1 | (x2 & ~x3))));
  assign n1690 = (~n686 | ~n1693) & (n1542 | n1692) & (x2 | n1691);
  assign n1691 = x0 ? (~x1 | ((~x6 | ~x7 | x3 | x4) & (~x3 | ~x4 | x6 | x7))) : (x1 | x3 | ~x4 | (x6 ^ x7));
  assign n1692 = (x0 | x2 | x4 | x6 | x7) & (~x4 | (x0 ^ ~x2) | (x6 ^ x7));
  assign n1693 = x7 & x6 & ~x3 & x4;
  assign n1694 = ~n1696 & n1697 & ~n1700 & (n437 | n1695) & ~n1701;
  assign n1695 = (~x4 | ((x0 | x1 | ~x2 | x3) & (~x0 | ~x1 | x2 | ~x3 | ~x5))) & ((x4 & x5) | ((x0 | ~x1 | x2 | ~x3) & (~x0 | x1 | (x2 ^ x3)))) & (~x2 | x3 | (x0 ? (~x1 | x4) : (x1 | ~x5)));
  assign n1696 = ~n520 & ((~x0 & ~n853) | (x2 & n654 & n321));
  assign n1697 = ~n1699 & (~x3 | ~n1070 | ~n460) & (n740 | ~n1698);
  assign n1698 = x5 & x3 & ~x0 & x2;
  assign n1699 = ~x0 & ((~x1 & ~x2 & x3 & x4 & ~x6) | (x1 & x2 & ~x3 & ~x4 & x6));
  assign n1700 = ~n950 & ((~x0 & ~x1 & ~x2 & ~x3 & x6) | (~x6 & ((x2 & x3 & ~x0 & x1) | (x0 & (x1 ? (~x2 & x3) : (x2 & ~x3))))));
  assign n1701 = n357 & ((~x0 & x1 & x4 & ~x5 & ~x6) | (x6 & ((~x0 & ~x1 & ~x4 & ~x5) | (x0 & (x1 ? (~x4 & ~x5) : (x4 & x5))))));
  assign z116 = n1704 | ~n1706 | ~n1713 | (~x1 & ~n1703);
  assign n1703 = (x3 | ((x2 | ((~x5 | x7 | x0 | x4) & (~x4 | (x0 ? (~x5 ^ x7) : (x5 ^ x7))))) & (x0 | ~x2 | x5 | (x4 ^ x7)))) & (x4 | x5 | ~x7 | x0 | x2 | ~x3);
  assign n1704 = ~x5 & ((~x0 & ~n1705) | (n292 & n361 & n459));
  assign n1705 = (x4 | ~x6 | x7 | x1 | x2 | x3) & (~x1 | ((x4 | ~x6 | ~x7 | x2 | ~x3) & (~x4 | x6 | x7 | ~x2 | x3)));
  assign n1706 = n1708 & n1709 & (n1707 | n1712) & (n425 | n1711);
  assign n1707 = x4 ? (~x5 | x6) : (x5 | ~x6);
  assign n1708 = (x3 | ~x4 | x7 | ~x0 | x1 | ~x2) & ((~x2 ^ x4) | (x1 ^ ~x3) | (~x0 ^ ~x7));
  assign n1709 = ~n1710 & (n811 | (~n288 & ~n361) | (~x0 & ~x7) | (x0 & x7));
  assign n1710 = (x3 ^ x7) & ((~x0 & x1 & x2 & x4) | (x0 & ~x1 & ~x2 & ~x4));
  assign n1711 = (x3 | x4 | ~x5 | ~x0 | ~x1 | x2) & (~x3 | ~x4 | x5 | x0 | x1 | ~x2);
  assign n1712 = (~x0 | ~x1 | x2 | ~x3 | x7) & (x0 | x1 | ~x2 | x3 | ~x7);
  assign n1713 = ~n1715 & ~n1716 & (~x5 | ~n1602 | n1714);
  assign n1714 = (~x3 | ((x1 | x2 | x6 | ~x7) & (~x1 | ~x2 | ~x6 | x7))) & (~x1 | x2 | x3 | (~x6 ^ x7));
  assign n1715 = ~x4 & n367 & ((x0 & ~x2 & x5 & ~x7) | (~x0 & x7 & (~x2 ^ ~x5)));
  assign n1716 = ~n467 & ((~x0 & x1 & ~x2 & x3 & ~x7) | (x0 & x7 & (x1 ? (~x2 & x3) : (x2 & ~x3))));
  assign z117 = ~n1722 | (x6 ? ~n1720 : (n1718 | n1719));
  assign n1718 = ~n891 & ((x2 & ~x3 & x4 & ~x5) | (~x0 & x3 & x5 & (~x2 ^ ~x4)));
  assign n1719 = x7 & n1167 & (x3 ? (x5 & n354) : (~x5 & n542));
  assign n1720 = (~n317 | ~n1209) & (~x2 | n1721);
  assign n1721 = (~x4 | ((x0 | ~x1 | ~x7 | (~x3 ^ x5)) & (x1 | x7 | ((x3 | ~x5) & (~x0 | ~x3 | x5))))) & (x3 | x4 | x5 | ((x1 | x7) & (x0 | ~x1 | ~x7)));
  assign n1722 = ~n1724 & ~n1725 & ~n1726 & ~n1727 & (~x0 | n1723);
  assign n1723 = (x2 | ((x1 | ~x3 | ~x4 | ~x5 | ~x6) & (~x1 | ((x5 | ~x6 | x3 | x4) & (~x5 | x6 | ~x3 | ~x4))))) & (x1 | ~x2 | ((~x5 | ~x6 | ~x3 | x4) & (x3 | x5 | (x4 ^ x6))));
  assign n1724 = x1 & x2 & ((~x3 & ~x4 & x5) | (~x0 & x3 & (~x4 ^ x5)));
  assign n1725 = ~x2 & (x1 ? (x3 ? (x4 & ~x5) : ((x4 & x5) | (~x0 & ~x4 & ~x5))) : ((~x3 & x4 & ~x5) | (~x4 & x5 & x0 & x3)));
  assign n1726 = (x3 ^ x5) & ((x1 & ~x2 & ~x4 & ~x6) | (~x1 & (x2 ? (x4 & ~x6) : (~x4 & x6))));
  assign n1727 = n783 & ((~x2 & x3 & x5 & ~n585) | (x2 & (x3 ? n1728 : (~x5 & ~n585))));
  assign n1728 = x6 & ~x4 & x5;
  assign z118 = n1730 | ~n1734 | (~n699 & ~n1733);
  assign n1730 = ~x3 & ((x0 & ~n1731) | (x6 & ~n1732 & ~x0 & x5));
  assign n1731 = (x5 | x6 | ~x7 | ~x1 | x2 | ~x4) & (x4 | ((~x1 | ((x6 | x7 | x2 | x5) & (~x6 | ~x7 | ~x2 | ~x5))) & (x5 | ~x6 | x7 | x1 | ~x2)));
  assign n1732 = (x1 | ~x2 | x4 | x7) & (x2 | ~x4 | ~x7);
  assign n1733 = x6 ? ((x3 | (x0 & x1) | (x2 ^ x5)) & (~x2 | ((x0 | (x1 ? (~x3 | x5) : ~x5)) & (~x0 | x1 | ~x3 | x5)))) : (x2 ? (x3 | x5) : (~x3 | ~x5));
  assign n1734 = n1737 & n1738 & (x5 ? n1736 : n1735);
  assign n1735 = (~x6 | (x0 ? (~x1 | x3 | (~x2 ^ x4)) : (~x3 | ((x2 | ~x4) & (x1 | ~x2 | x4))))) & (~x3 | x6 | (x2 ? (~x4 | (x0 & x1)) : x4));
  assign n1736 = (x4 & (~x2 | (x0 & x1))) | (x6 & (~x3 | (~x0 & ~x1))) | (x3 & ~x6) | (x2 & ~x4);
  assign n1737 = (~n464 | ~n866) & (~n870 | ~n313 | ~n460);
  assign n1738 = (x0 | n1740) & (n1739 | (x3 ? n1085 : ~n531));
  assign n1739 = (x0 | ~x1 | ~x2 | x4 | x7) & (~x0 | ((x2 | ~x4 | ~x7) & (x4 | x7 | x1 | ~x2)));
  assign n1740 = (x1 | ~x3 | ~x5 | (x2 ? (~x4 | ~x7) : (x4 | x7))) & (x3 | x5 | (x2 ? (x4 | x7) : (~x4 | ~x7)));
  assign z119 = ~n1745 | (~x4 & (~n1743 | (~n425 & ~n1742)));
  assign n1742 = (x0 | x1 | x3 | ~x5) & (x5 | (x0 ? (x1 ? (~x2 | x3) : (x2 | ~x3)) : (~x1 | ~x3)));
  assign n1743 = (x6 | n1744) & (~x3 | ~x5 | ~x6 | x7 | ~n317);
  assign n1744 = (x0 & ((x1 & x2) | ~x7)) | (~x3 & (~x5 | ~x7)) | (x3 & x5 & x7) | (~x7 & (x1 ? ~x5 : ~x2));
  assign n1745 = n1748 & (n399 | n1746) & (n1054 | n1747);
  assign n1746 = (x0 & x1 & (x2 | (x6 & ~x7))) | (~x1 & ((~x4 & x7) | (~x2 & ((~x4 & ~x6) | (~x0 & x6 & ~x7))))) | (~x6 & x7) | (x4 & x6 & ~x7) | (~x0 & ~x4 & (~x6 | x7));
  assign n1747 = (~x4 | x6 | ~x7 | x2 | ~x3) & (x7 | ((~x4 | ~x6 | x2 | x3) & (x1 | ((x3 | ~x4 | ~x6) & (x4 | x6 | x2 | ~x3)))));
  assign n1748 = (n437 | n1749) & (n1750 | (x2 ? n589 : ~n1070));
  assign n1749 = (~x1 | ~x2 | ((x4 | ~x5 | ~x0 | x3) & (~x4 | x5 | x0 | ~x3))) & (x0 | x1 | x2 | x3 | x4 | x5) & (~x4 | (x0 ? (~x3 | (x1 & x2) | x5) : (x3 | ~x5)));
  assign n1750 = x0 ? ((~x5 | ~x7 | x1 | ~x3) & (x5 | x7 | ~x1 | x3)) : (~x3 | ~x7 | (~x1 ^ ~x5));
  assign z120 = ~n1757 | (x1 ? ~n1752 : (x4 ? ~n1755 : ~n1756));
  assign n1752 = n1754 & (x3 | n1753);
  assign n1753 = (x5 | ~x6 | x7 | x0 | ~x2 | ~x4) & (~x0 | x4 | ((~x6 | ~x7 | x2 | x5) & (~x2 | (x5 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n1754 = (x0 | ((~x5 | ~x7 | ~x2 | x4) & (x6 | x7 | ~x4 | x5))) & (x2 | x4 | ((~x5 | ~x6 | ~x7) & (x6 | x7 | ~x0 | x5)));
  assign n1755 = (~x6 | ~x7 | x0 | ~x5) & (x7 | ((~x0 | ~x2 | ~x3 | ~x5 | ~x6) & (x6 | ((x2 | x3 | x5) & (x0 | (x5 & (x2 | ~x3)))))));
  assign n1756 = (~x7 | (x0 ? (~x6 | (~x5 & (~x2 | ~x3))) : (x5 | x6 | (x2 ^ ~x3)))) & (~x0 | ~x2 | x5 | x6 | x7);
  assign n1757 = (n434 | n1758) & (n665 | n1759);
  assign n1758 = (x0 | ~x1 | ~x2 | ~x3 | ~x4) & ((x1 & x2) | (~x0 ^ ~x4));
  assign n1759 = (~x4 & ((~x2 & ((~x0 & ~x1) | (~x3 & x6))) | (~x1 & x6) | (~x0 & (x6 | (~x1 & ~x3))))) | (x4 & ~x6 & (x1 | x2 | x3)) | (x0 & ((x1 & (x4 | (x2 & x3))) | (x4 & ~x6) | (x2 & x3 & x6)));
  assign z121 = ~n1767 | (x4 ? ~n1763 : (x0 ? ~n1761 : ~n1762));
  assign n1761 = (x1 | ((x5 | ~x6 | x7) & (~x5 | x6 | ~x7) & (~x2 | x3 | (x5 ^ x7)))) & (x2 | x3 | (x5 ? (x6 | ~x7) : (~x6 | x7)));
  assign n1762 = (~x2 & ((~x6 & ~x7) | (x3 & x6 & x7) | (~x1 & ~x3 & (~x6 | ~x7)))) | (x2 & (x1 | (~x3 & x6 & x7))) | (x5 & x7) | (~x7 & (~x5 | (~x3 & ~x6)));
  assign n1763 = (n1042 | n1765) & (~x0 | x1 | n1766) & (x0 | n1764);
  assign n1764 = ((x5 ? (~x6 | x7) : (x6 | ~x7)) | (x1 ^ ~x2)) & (x5 | x6 | ~x7 | x2 | ~x3) & (~x2 | ((x1 | (x3 ? (x5 | ~x7) : (~x5 | x7))) & (~x5 | x6 | ~x7 | ~x1 | ~x3)));
  assign n1765 = (x0 | x1 | ~x3 | ~x5 | x7) & (~x0 | ((x3 | x5 | x7) & (~x5 | ~x7 | x1 | ~x3)));
  assign n1766 = x2 ? ((x5 | ~x6 | x7) & (x3 | ~x5 | ~x7)) : ((~x5 | x6 | ~x7) & (~x3 | x5 | x7));
  assign n1767 = x6 ? (x7 ? n1769 : n1768) : (x7 ? n1768 : n1769);
  assign n1768 = x0 ? (~x1 | ~x5 | (~x2 ^ (x3 | x4))) : ((x1 | x2 | x3 | ~x5) & (~x1 | ~x2 | x5));
  assign n1769 = x1 ? (x0 ? (x5 | (x2 & (x3 | x4))) : ~x5) : ((x5 | ((~x2 | (~x0 ^ ~x3)) & (x0 | (x3 ? x2 : ~x4)))) & (~x0 | x2 | (x3 & x4) | ~x5));
  assign z122 = ~n1779 | n1778 | n1776 | n1773 | n1771 | n1772;
  assign n1771 = ~x4 & ((x0 & ((x3 & x6 & x1 & ~x2) | (~x3 & ~x6 & ~x1 & x2))) | (x1 & x2 & ~x3 & x6) | (~x0 & (x1 ? (x2 ? x6 : (~x3 & ~x6)) : (x2 ? (x3 & ~x6) : (~x3 & x6)))));
  assign n1772 = x4 & ((x2 & ((~x0 & (x1 ? (~x3 & x6) : (x3 & ~x6))) | (x0 & ~x1 & ~x3 & ~x6))) | (x0 & ~x2 & x3 & (~x1 ^ x6)));
  assign n1773 = ~x4 & (n1774 | n1775 | (n374 & n459 & n335));
  assign n1774 = ~n425 & ((~x0 & x1 & ~x2 & x3) | (x0 & ((x1 & ~x2 & ~x3) | (x3 & x5 & ~x1 & x2))));
  assign n1775 = ~x3 & n349 & (x2 ? (~x5 & n372) : (x5 & n374));
  assign n1776 = x0 & (x1 ? (n357 & n1777) : (n358 & n1038));
  assign n1777 = x6 & x4 & x5;
  assign n1778 = n1050 & ((x1 & x2 & x3 & n450) | (~x1 & ~x3 & (x2 ? n451 : n450)));
  assign n1779 = (n437 | n1780) & (~x4 | (~n1781 & (x3 | n1782)));
  assign n1780 = (x0 | ((~x1 | ~x2 | ~x3 | ~x4 | ~x5) & (x1 | (x2 ? (x3 | x4) : ~x3)))) & (x1 | x2 | (x3 ? x4 : ~x0));
  assign n1781 = ~n425 & ((x0 & ~x1 & x2 & x3) | (x1 & ~x2 & (~x0 | n784)));
  assign n1782 = (~x5 | x6 | x7 | ~x0 | ~x1 | x2) & (x0 | x1 | ((~x6 | x7 | x2 | ~x5) & (x6 | ~x7 | ~x2 | x5)));
  assign z123 = ~n1787 | (~x5 & ~n1784) | (x5 & n357 & ~n1786);
  assign n1784 = (~x2 | n1785) & (~n543 | ~n288 | ~n317);
  assign n1785 = x0 ? ((x4 | ~x6 | ~x7 | x1 | ~x3) & (~x4 | x6 | x7 | ~x1 | x3)) : (x3 | ((~x6 | x7 | ~x1 | x4) & (x1 | ~x4 | (~x6 ^ x7))));
  assign n1786 = (x0 | x1 | ~x4 | ~x6 | ~x7) & (~x1 | (x0 ? (~x4 | (~x6 ^ x7)) : (x4 | (x6 ^ x7))));
  assign n1787 = ~n1788 & ~n1789 & ~n1790 & (x4 | n1712) & n1791;
  assign n1788 = x4 & ((~x2 & (x0 ? (x3 & ~x7) : (x1 ? (x3 & x7) : (~x3 & ~x7)))) | (x0 & ~x1 & x2 & (~x3 ^ x7)));
  assign n1789 = (x3 ^ x4) & ((~x0 & x1 & (x2 ^ x7)) | (x0 & ~x1 & ~x2 & x7));
  assign n1790 = n357 & ((x0 & x1 & x4 & ~x5 & x7) | (~x0 & ~x4 & ~x7 & (~x1 ^ ~x5)));
  assign n1791 = ~n1792 & (~x2 | n1793);
  assign n1792 = (x2 ^ x7) & (x0 ? (~x3 & ~x4) : (~x1 & x3));
  assign n1793 = (~x3 | (x5 ^ x7) | (x0 ? (x1 | x4) : (~x1 | ~x4))) & (x0 | x3 | ~x5 | x7 | (x1 ^ ~x4));
  assign z124 = n1796 | n1797 | ~n1799 | (~x3 & ~n1795) | ~n1801;
  assign n1795 = (~x4 | (x0 ? (x2 | (x1 ? (~x5 | ~x6) : (x5 | x6))) : (~x2 | (x1 ? (~x5 | x6) : (x5 | ~x6))))) & (x0 | ~x1 | x4 | ~x6 | (~x2 ^ x5));
  assign n1796 = ~x2 & (x0 ? (x1 ? (x3 & ~x4) : (~x3 ^ x4)) : (x1 ? (~x3 & x4) : (x3 & ~x4)));
  assign n1797 = ~n1798 & x5 & n1050;
  assign n1798 = (~x1 | ~x2 | x3 | ~x6 | x7) & (x1 | x2 | (x3 ? (x6 | x7) : (~x6 | ~x7)));
  assign n1799 = n1800 & (~n1548 | ((x0 | ~x1 | x3 | ~x5) & (~x0 | x1 | (x3 ^ x5))));
  assign n1800 = ~x3 | ((~x0 | x1 | ~x2 | ~x4) & (x0 | x4 | (x1 ? (x2 | ~n312) : ~x2)));
  assign n1801 = x4 ? n1802 : ((~n459 | ~n1586) & (x5 | n1803));
  assign n1802 = (~x0 | ~x1 | x2 | ~x3 | x5) & (x0 | ((x1 | x2 | ~x3 | x5) & (~x2 | (x1 ? (x3 ^ x5) : (x3 | ~x5)))));
  assign n1803 = x0 ? ((x1 | ~x2 | ~x3 | ~x6 | ~x7) & (~x1 | x2 | x3 | x6 | x7)) : (~x1 | ((~x6 | x7 | x2 | ~x3) & (x6 | ~x7 | ~x2 | x3)));
  assign z125 = n1807 | ~n1808 | ~n1812 | (x0 ? ~n1806 : ~n1805);
  assign n1805 = (~x4 | x5 | x6 | ~x1 | x2 | ~x3) & (x1 | ((x4 | ~x5 | x6 | x2 | ~x3) & (~x2 | ~x4 | (x3 ? (~x5 | x6) : (x5 | ~x6)))));
  assign n1806 = (x3 | ~x6 | ((x1 | ~x2 | x4 | ~x5) & (x2 | (x1 ? (x4 ^ x5) : (~x4 | x5))))) & (~x4 | x5 | x6 | x1 | ~x2 | ~x3);
  assign n1807 = ~n368 & ((~x1 & ~x2 & x3 & x4 & x5) | (~x3 & ~x4 & (x1 ? (~x2 ^ ~x5) : (~x2 & ~x5))));
  assign n1808 = ~n1809 & n1811 & (n1010 | n1810);
  assign n1809 = ~x1 & ((x3 & x4 & ~x5 & ~x0 & x2) | (~x2 & (x3 ^ x5) & (x0 ^ ~x4)));
  assign n1810 = (~x0 | x1 | ~x3 | x4 | x5) & (x0 | ~x1 | x3 | ~x4 | ~x5);
  assign n1811 = ((x4 ^ x5) | ((x0 | ~x2 | (~x1 ^ ~x3)) & (~x0 | ~x1 | x2 | ~x3))) & (x3 | x4 | ~x5 | x0 | ~x1 | ~x2) & ((x0 ? (x1 | ~x2) : (~x1 | x2)) | (x3 ? (x4 | ~x5) : (~x4 | x5)));
  assign n1812 = x2 ? n1814 : (~n1813 & (~x5 | n672 | n798));
  assign n1813 = n1354 & ((~x0 & x1 & x3 & x6 & x7) | (~x3 & ((~x0 & ~x1 & ~x6 & x7) | (x0 & (x1 ? (~x6 & x7) : (x6 & ~x7))))));
  assign n1814 = (x4 | n1815) & (x0 | ~n647 | ~n996);
  assign n1815 = (x3 | ((~x0 | ((x6 | ~x7 | x1 | ~x5) & (~x6 | x7 | ~x1 | x5))) & (x5 | x6 | ~x7 | x0 | ~x1))) & (x0 | ~x3 | x6 | x7 | (~x1 ^ ~x5));
  assign z126 = n1818 | ~n1820 | ~n1824 | (x1 ? ~n1819 : ~n1817);
  assign n1817 = (x5 | ((x0 | (x2 ? (~x3 | (~x4 ^ x6)) : (x3 | (~x4 & ~x6)))) & (~x0 | x2 | ~x3 | x4 | ~x6))) & (~x4 | ~x5 | ((~x2 | x3 | x6) & (x0 | x2 | ~x3 | ~x6)));
  assign n1818 = ~n416 & ((~x4 & (x0 ? (x1 ? (~x2 & x3) : (x2 & ~x3)) : (x1 ? (~x2 ^ x3) : (~x2 & x3)))) | (x0 & ~x2 & x4 & (~x1 ^ ~x3)));
  assign n1819 = x3 ? (~x4 | ~x5 | (x2 ? x0 : x6)) : ((x4 | ((~x0 | (x2 ? (~x5 | x6) : (x5 | ~x6))) & (x5 | ~x6 | x0 | ~x2))) & (x0 | ~x4 | (x2 ? (x5 | x6) : (~x5 | ~x6))));
  assign n1820 = n1821 & (n420 | ((x1 | (x0 ? (x2 ^ x3) : (~x2 | x3))) & (x0 | ~x1 | x2 | ~x3)));
  assign n1821 = x4 ? (x7 | ((~x6 | n1822) & (x1 | x6 | n1823))) : (~x7 | ((x6 | n1822) & (~x1 | ~x6 | n1823)));
  assign n1822 = (~x0 | ~x5 | (x1 ? (x2 | ~x3) : (~x2 | x3))) & (x5 | (x0 ^ ~x2) | (x1 ^ ~x3));
  assign n1823 = (x0 | x2 | ~x3 | x5) & (~x0 | x3 | (x2 ^ ~x5));
  assign n1824 = (x1 | n1825) & (x0 | ~x1 | n1829);
  assign n1825 = (n1826 | n1828) & (~n269 | ~n1461) & (~x5 | n1827);
  assign n1826 = ~x2 ^ ~x3;
  assign n1827 = (x7 | ((x0 | ~x2 | x3 | x4 | ~x6) & (~x0 | ((~x2 | ~x3 | ~x4 | x6) & (x2 | x3 | x4 | ~x6))))) & (~x4 | x6 | ~x7 | x0 | x2 | ~x3);
  assign n1828 = (x0 | ~x5 | (x4 ? (~x6 | ~x7) : (x6 | x7))) & (~x0 | x4 | x5 | ~x6 | ~x7);
  assign n1829 = (~x5 | ((~x7 | ((~x2 | (x3 ? (x4 | x6) : (~x4 | ~x6))) & (x2 | x3 | ~x4 | x6))) & (x2 | ~x3 | x4 | ~x6 | x7))) & (~x4 | x5 | x6 | x7 | (~x2 ^ ~x3));
  assign z127 = ~n1831 | n1843 | (~n437 & ~n1842);
  assign n1831 = n1839 & n1837 & ~n1836 & ~n1832 & ~n1835;
  assign n1832 = ~x2 & ((~x4 & ~n1833) | (x5 & n361 & ~n1834));
  assign n1833 = ((~x0 ^ ~x7) | ((~x5 | ~x6 | ~x1 | x3) & (x5 | x6 | x1 | ~x3))) & (x0 | ~x1 | x5 | (x3 ? (~x6 | ~x7) : (x6 | x7)));
  assign n1834 = (x0 | x1 | x6 | ~x7) & (~x0 | (x1 ? (~x6 | ~x7) : (x6 | x7)));
  assign n1835 = ~n515 & ((~x5 & ((~x0 & (x1 ? (x3 & x6) : (~x3 & ~x6))) | (x0 & ~x1 & ~x3 & x6))) | (x0 & x5 & x6 & (~x1 ^ ~x3)));
  assign n1836 = ~n1591 & ((~x0 & x1 & ~x2 & x4 & x5) | (x0 & ~x5 & (x1 ? (~x2 & ~x4) : (x2 & x4))));
  assign n1837 = (~x2 | x3 | ~x4 | n1838) & (~x3 | ((~x4 | ~n686 | ~n312) & (x2 | x4 | n1838)));
  assign n1838 = (~x0 | x1 | ~x5 | x6) & (x0 | (x1 ? (x5 | x6) : ~x6));
  assign n1839 = (~x1 | n1840) & (n425 | n1841);
  assign n1840 = (x4 | x5 | ~x6 | x0 | x2 | x3) & (x6 | (x0 ? (x2 | (x3 ? ~x4 : (x4 | ~x5))) : (~x2 | ~x5 | (x3 ^ x4))));
  assign n1841 = ((~x2 ^ x4) | ((x0 | x1 | x3 | ~x5) & (~x0 | x5 | (x1 ^ ~x3)))) & (~x0 | x1 | x2 | x3 | x4) & (x0 | ~x5 | ((~x3 | ~x4 | x1 | ~x2) & (~x1 | (x2 ? (x3 | ~x4) : (~x3 | x4)))));
  assign n1842 = ((x2 ? (x3 ^ x4) : (x3 | ~x4)) | (x0 ? (x1 | ~x5) : (~x1 | x5))) & (x0 | x1 | x2 | x3 | x4) & (~x3 | ((x0 | x1 | x2 | ~x4 | x5) & (x4 | ((~x0 | ~x1 | x2 | ~x5) & (x0 | ~x2 | (x1 ^ x5))))));
  assign n1843 = x2 & ((~x1 & ~n1844) | (n351 & n374 & n1585));
  assign n1844 = (x0 | ~x4 | x5 | (x3 ? (~x6 | ~x7) : (x6 | x7))) & (~x5 | ((x4 | x6 | ~x7 | x0 | ~x3) & (~x0 | ((~x6 | ~x7 | x3 | ~x4) & (x6 | x7 | ~x3 | x4)))));
  assign z128 = ~n1848 | (x5 & ~n1854) | (~x5 & ~n1853) | (x7 & ~n1846);
  assign n1846 = (~x4 | n1847) & (x2 | x4 | n1231 | (~x1 ^ ~x6));
  assign n1847 = x2 ? ((x1 | ((x3 | x5 | x6) & (~x0 | ~x6 | (~x3 ^ x5)))) & (x0 | ~x1 | x3 | (~x5 ^ x6))) : (~x3 | ~x5 | (x1 ^ x6));
  assign n1848 = n1850 & (x7 | (~n1849 & (~n531 | ~n373 | ~n459)));
  assign n1849 = n357 & (x1 ? (x6 & ((~x4 & ~x5) | (~x0 & x4 & x5))) : (~x6 & ((x4 & x5) | (x0 & ~x4 & ~x5))));
  assign n1850 = (n1345 | n1852) & (n1851 | (~n342 & ~n1029));
  assign n1851 = (x1 | x4 | x5 | ~x7) & (~x4 | (x1 ? (~x5 | x7) : (x5 ^ x7)));
  assign n1852 = (~x4 | x5 | x7 | ~x2 | x3) & (~x3 | ((x2 | x7 | (x4 ^ x5)) & (x0 | ~x2 | (x4 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n1853 = x1 ? (x2 ? (x4 | ((x3 | ~x7) & (x0 | ~x3 | x7))) : (~x4 | (~x3 ^ x7))) : ((x4 | x7 | ~x2 | x3) & (~x4 | ~x7 | x2 | ~x3) & ((~x4 ^ x7) | (x0 ? (~x2 | ~x3) : (x2 | x3))));
  assign n1854 = x7 ? ((x0 | ((~x1 | ~x3 | x4) & (x1 | x2 | x3 | ~x4))) & (~x1 | x2 | ~x3 | x4) & (x1 | ~x2 | ((x3 | x4) & (~x0 | ~x3 | ~x4)))) : (x1 ? (x3 | x4) : (x2 ? (x3 | ~x4) : (~x3 | x4)));
  assign z129 = n1858 | n1860 | ~n1861 | (~x3 & (n1856 | n1857));
  assign n1856 = (~x2 ^ ~x7) & ((~x0 & x4 & x5 & ~x6) | (~x4 & (~x5 ^ x6)));
  assign n1857 = n654 & ((x0 & ~x1 & ~x2 & ~x6 & x7) | (x6 & ((x0 & ((~x2 & ~x7) | (~x1 & x2 & x7))) | (x1 & ((~x0 & x2 & x7) | (~x2 & ~x7))))));
  assign n1858 = ~n1859 & (~x0 | n321);
  assign n1859 = x2 ? (x3 ? (x4 ? (~x5 | x6) : (x5 ^ x6)) : (x4 ? (x5 | ~x6) : (~x5 | x6))) : (x4 ? ((x5 | x6) & (~x3 | ~x5 | ~x6)) : (x5 | ~x6));
  assign n1860 = n595 & ((~x6 & ((x2 & ~x3 & ~x4 & x5) | (~x2 & x4 & (~x3 | ~x5)))) | (~x2 & x6 & ((~x4 & ~x5) | (x3 & x4 & x5))));
  assign n1861 = (x3 | ~x4 | ~x5 | ~x6 | ~n317) & (~x3 | n1862 | (x4 ? (x5 | ~x6) : (~x5 | x6)));
  assign n1862 = x7 ? (~x2 | (x0 & x1)) : x2;
  assign z130 = ~n1866 | ~n1867 | (~n864 & ~n1864) | (~n425 & ~n1865);
  assign n1864 = (x4 & ((x6 & ~x7) | (~x0 & ((x5 & x6) | (~x3 & ~x7))))) | (~x3 & (~x5 | (x6 & ~x7))) | (x3 & x5 & x7) | (~x6 & ((~x4 & x7) | (x3 & x5 & (x0 | ~x4))));
  assign n1865 = x3 ? ((x1 | x2 | x5) & (x0 | (x1 ? (~x2 | x5) : (x2 | ~x4)))) : (x4 | ~x5 | (x1 ^ x2));
  assign n1866 = (~n462 | ~n284) & (n399 | n678 | n1168);
  assign n1867 = (n1868 | n1869) & (x3 | ~x7 | n1870);
  assign n1868 = (x1 | x2) & (x0 | ~x1 | ~x2);
  assign n1869 = (x3 | ~x4 | ~x5 | x6 | ~x7) & (~x3 | ((x6 | ~x7 | ~x4 | x5) & (x4 | ~x6 | x7)));
  assign n1870 = (~x0 | ((x1 | x2 | ~x4 | ~x5 | ~x6) & (~x1 | ~x2 | x4 | x5 | x6))) & (x0 | ~x1 | ~x4 | ~x5 | ~x6);
  assign z131 = n1872 | ~n1875 | (~n950 & ~n1874);
  assign n1872 = ~x7 & ((~x3 & ~n1873) | (x3 & x6 & ~n1015 & ~n1168));
  assign n1873 = (x5 | ((x4 | ~x6) & (~x0 | ~x1 | ~x2 | ~x4 | x6))) & (~x4 | ~x5 | ~x6 | (x0 & x1 & x2));
  assign n1874 = (x0 | x6 | x7) & (x1 | ((x6 | x7 | x2 | x3) & (x0 | ~x6 | ~x7 | (x2 & x3))));
  assign n1875 = ~n1876 & ~n1877 & n1879 & (~x0 | x6 | n1878);
  assign n1876 = (~x1 ^ ~x2) & ((~x4 & ~x6 & x7) | (x0 & x4 & (~x6 ^ x7)));
  assign n1877 = x7 & ((~x0 & x1 & ((x4 & x6) | (x2 & ~x4 & ~x6))) | (~x1 & ~x2 & ((~x4 & ~x6) | (x0 & x4 & x6))));
  assign n1878 = (x1 | x2 | ~x3 | ~x4 | x7) & (~x1 | ~x2 | x3 | x4 | ~x7);
  assign n1879 = ~n374 | ((~n686 | ~n361) & (~n850 | ~n866));
  assign z132 = ~n1882 | (~x1 & (n1881 | (x0 & n509 & n464)));
  assign n1881 = ~x0 & x7 & ((n358 & n1174) | (n357 & n1175));
  assign n1882 = ~n1885 & n1887 & (x6 | ~n1883 | (n864 & n1884));
  assign n1883 = x0 & x5;
  assign n1884 = (~x1 | ~x2 | x3 | x4) & (x1 | x2 | ~x3 | ~x4);
  assign n1885 = ~n440 & ~n1886;
  assign n1886 = x0 ? ((x3 & ((x1 & x2) | (x4 & ~x6))) | (x2 & ~x6) | (x1 & (~x6 | (x2 & x4)))) : (~x1 & (((~x3 | ~x4) & x6) | (~x2 & (x6 | (~x3 & ~x4)))));
  assign n1887 = (~n686 | ~n1888) & (~n450 | ((~n686 | ~n373) & (x2 | ~n783)));
  assign n1888 = x6 & ~x3 & ~x5;
  assign z133 = ~n1891 | n1892 | n1894 | (x0 ? ~n1890 : ~n1893);
  assign n1890 = (~x4 | x6 | x7 | x1 | x2 | ~x3) & (~x1 | ~x2 | x3 | x4 | (x6 ^ x7));
  assign n1891 = (x7 | (x1 ^ ~x2) | (~x0 ^ x6)) & (~x0 | ~x6 | ((x2 | ~x7) & (x1 | (~x7 & (x2 | x3)))));
  assign n1892 = n719 & n509 & n321;
  assign n1893 = (x1 | x6 | ~x7) & (~x6 | (x1 ^ (x2 | x7)));
  assign n1894 = n1230 & (x0 ? (n1671 & n612) : (n647 & n611));
  assign z134 = n1897 | ~n1899 | (~x1 & (~n1896 | (~x0 & ~n1898)));
  assign n1896 = (~x4 | x5 | x7 | x0 | ~x2 | ~x3) & (x2 | x4 | ((~x5 | x7 | x0 | x3) & (~x0 | ~x3 | (~x5 ^ x7))));
  assign n1897 = ~x7 & (x0 ? ((x1 & x2 & ~x3 & ~x4) | (x3 & x4 & ~x1 & ~x2)) : (~x1 & (x2 ? (x3 & ~x4) : (~x3 & x4))));
  assign n1898 = (x5 | ~x6 | x7 | x2 | x3 | x4) & (~x2 | ~x3 | ~x4 | ~x5 | (x6 ^ x7));
  assign n1899 = (x0 | ((~x1 | ~x7) & (x1 | x2 | ~x3 | x7))) & (~x1 | ((~x0 | x2 | x7) & (~x7 | ~n339 | ~x2 | x3))) & (x3 | x7 | x1 | ~x2) & (~x0 | ((x7 | ~n339 | ~x2 | x3) & (x1 | (x2 ? x7 : (x3 | ~x7)))));
  assign z135 = ~n1903 | n1904 | n1905 | (~x1 & (~n1901 | ~n1902));
  assign n1901 = (x0 | x2 | x3 | x4 | ~x5) & (~x3 | ((x0 | x2 | x4 | x5) & (~x0 | (x2 ? (~x4 | x5) : (x4 | ~x5)))));
  assign n1902 = (x0 | ~x6 | ((x4 | x5 | x2 | x3) & (~x2 | ~x3 | ~x4 | ~x5))) & (~x0 | ~x2 | ~x3 | ~x4 | ~x5 | x6);
  assign n1903 = (~x2 | ((x3 | x4 | x0 | ~x1) & (~x0 | x1 | (x3 & x4)))) & (x0 | ~x1 | x2 | ~x4) & (~x3 | (x0 ? (x1 | ~x4 | (x2 & ~n996)) : (~x1 | x2)));
  assign n1904 = ~x0 & ~x2 & ~x3 & (~x1 ^ ~x4);
  assign n1905 = n544 & n312 & ((n1906 & n369) | (n345 & n370));
  assign n1906 = x1 & x2;
  assign z136 = n1910 | (n487 & ~n1908) | (~x1 & ~n1909);
  assign n1908 = (~x4 & (~x1 | ~x3)) | (~x3 & (~x1 | (~x5 & ~x6 & ~x7))) | (x3 & x4 & x5 & x6 & x7) | (~x1 & (~x5 | ~x6));
  assign n1909 = (~x2 | x3 | (x4 & (x5 | x6 | x7))) & (~x3 | ((~x6 | ~x7 | ~x4 | ~x5) & (x2 | (~x4 & ~x5))));
  assign n1910 = x1 & ~x2 & (~x3 | (~x4 & ~x5));
  assign z137 = n1912 | ~n1913;
  assign n1912 = ~x2 & ((x0 & x1 & x3 & x4 & ~x5) | (~x4 & ((x1 & ~x3 & ~x5) | (x0 & (x5 ? x1 : ~x3)))));
  assign n1913 = n1414 & ~n1918 & (~x4 | (~n1914 & n1916 & n1919));
  assign n1914 = ~n1915 & (x0 ? (~x2 & ~x7) : (x2 & x7));
  assign n1915 = (x3 | x5 | x6) & (~x1 | ~x3 | ~x5 | ~x6);
  assign n1916 = (~x2 | ~x7 | ~n321 | n671) & (x2 | x7 | n1917);
  assign n1917 = (x5 | x6 | x0 | x3) & (~x0 | x1 | ~x3 | ~x5 | ~x6);
  assign n1918 = (~x2 | (~x4 ^ x5)) & (x2 | (x4 ^ x5)) & (~x0 | ~x1) & (x3 | x5) & (~x3 | ~x4 | ~x5);
  assign n1919 = (~x5 | x6 | x2 | ~x3) & (~x2 | ~x6 | ((x1 | x3 | x5) & (x0 | ((x3 | x5) & (x1 | ~x3 | ~x5)))));
  assign z138 = (~x7 & (n1922 | n1923)) | ~n1925 | (x4 & ~n1921);
  assign n1921 = (x1 | ((x5 | x6 | (~x3 ^ x7)) & (~x0 | ~x5 | ~x6 | (~x3 ^ ~x7)))) & (x0 | ((x6 | ~x7 | x3 | x5) & (~x3 | ((x5 | x6 | x7) & (~x6 | ~x7 | ~x1 | ~x5)))));
  assign n1922 = ~x0 & (x1 ? (n509 & n1777) : (n929 & n1038));
  assign n1923 = n1924 & ((x5 & ~n1096) | (x4 & ~x5 & ~n798));
  assign n1924 = ~x2 & x0 & x1;
  assign n1925 = ~n1926 & ~n1927 & ~n1928 & (x0 | ~n269 | ~n273);
  assign n1926 = ~x4 & (x3 ? (x5 & (~x0 | ~x1)) : (~x5 & (x0 | x1 | x6)));
  assign n1927 = x4 & ((~x3 & (~x0 | ~x1) & (x5 ^ x6)) | (~x0 & ~x1 & x3 & x5 & x6));
  assign n1928 = n595 & n1929 & ((x3 & ~x4 & x5) | (x4 & (x5 ? ~n520 : ~x3)));
  assign n1929 = ~x2 & x7;
  assign z139 = ~n1932 | (~x3 & ~n1931);
  assign n1931 = (~x4 | x5 | x6 | ~x7 | ~n317) & (x4 | x7 | ~n1192 | (x5 ^ x6));
  assign n1932 = (~x5 | n1934) & (n307 | n1933) & (n420 | n1168);
  assign n1933 = (x1 & x2 & (x0 | (~x3 & x6))) | (~x5 & x6) | (x5 & ~x6) | (~x0 & ((~x2 & x6) | (~x1 & (x6 | (~x2 & ~x3)))));
  assign n1934 = (x3 | ((~x0 | ~x1 | ~x2 | x4 | x6) & (x0 | ~x4 | ~x6))) & (x0 | ~x4 | (x1 & x2) | ~x6);
  assign z140 = n1937 | ~n1938 | (n542 & ~n1936);
  assign n1936 = (x0 | ~x3 | ~x5 | ~x6 | x7) & (~x0 | ((x5 | ~x6 | x7) & ((~x3 & ~x4) | (x5 ? (x6 ^ x7) : (x6 | ~x7)))));
  assign n1937 = ~n1301 & (x5 ? (~x6 ^ x7) : (x6 ? (~x7 & n1906) : x7));
  assign n1938 = ~n1940 & (n1939 | (~n780 & (~x5 | n425)));
  assign n1939 = x0 ? (x1 | (~x3 & ~x4)) : (x3 & x4);
  assign n1940 = x6 & ~x7 & (x0 ? (~x1 & ~x5) : (x5 & (~x1 | ~x3)));
  assign z141 = ~n1944 | n1946 | (n1602 & ~n1942) | (~x6 & ~n1943);
  assign n1942 = (~x1 | ~x2 | ~x3 | x5 | ~x6 | x7) & (~x5 | x6 | ~x7 | x1 | x2 | x3);
  assign n1943 = (~x0 | ~x1 | ~x2 | x3 | x4) & (x0 | ~x4 | ((x1 | x2 | x3 | ~x7) & (~x1 | ~x2 | ~x3 | x7)));
  assign n1944 = ~n1945 & ((x0 & (x6 | (x1 & x2))) | (~x0 & ((~x6 & ~x7) | (~x1 & ~x2 & x7))) | (x6 & x7) | (x1 & x2 & ~x7));
  assign n1945 = n958 & n339;
  assign n1946 = ~x0 & ((~x1 & ~x2 & x3 & ~x6 & x7) | (x1 & x2 & ~x3 & x6 & ~x7));
  assign z142 = n1948 | n1950 | (n1602 & (~n1949 | (~x7 & ~n1288)));
  assign n1948 = ~x0 & ((x1 & ((x4 & x7 & x2 & x3) | (~x3 & ~x7))) | (~x7 & (x3 ? (~x1 | ~x2) : (x2 | x4))));
  assign n1949 = x1 ? (~x2 | ~x3 | ~x5 | (x6 ^ x7)) : (x2 | x3 | x5 | (~x6 ^ x7));
  assign n1950 = x0 & x7 & (~x1 | ~x2 | (~x3 & ~x4));
  assign z143 = ~n1952 | ~n1953;
  assign n1952 = (~x0 | x1 | ~x2 | ~x3) & (~x1 | (x2 & (x3 | x4) & (x0 | (x3 & (x4 | ~n451)))));
  assign n1953 = (x3 | x5 | x6 | n1428) & (~x3 | ~n487 | n1513);
  assign z144 = n1956 | ~n1958 | (n1929 & ~n1955) | (x1 & ~n1957);
  assign n1955 = x0 ? ((x4 | x5 | ~x6 | x1 | ~x3) & (~x4 | ~x5 | x6 | ~x1 | x3)) : ((~x1 | ~x3 | ~x4 | x5 | x6) & (x1 | ((~x5 | ~x6 | ~x3 | ~x4) & (x5 | x6 | x3 | x4))));
  assign n1956 = x3 & ((x0 & ~x1 & ~x2 & ~x4 & x5) | (~x0 & ((x4 & ~x5 & ~x1 & x2) | (x1 & (x2 ? (~x4 & ~x5) : (x4 & x5))))));
  assign n1957 = (~x0 | x2 | x3 | ~x4 | ~x5 | ~x6) & (x0 | ~x3 | ((x5 | ~x6 | x2 | ~x4) & (~x5 | x6 | ~x2 | x4)));
  assign n1958 = n1319 & ((~n929 & (~x0 | ~x1)) | (~n509 & (~n929 | (x0 & x1 & ~n339))));
  assign z145 = n1960 | n1963 | n1965 | ~n1966 | (~x1 & ~n1964);
  assign n1960 = ~x5 & ((n522 & ~n1962) | (~x6 & ~n1961));
  assign n1961 = x0 ? (~x2 | x3 | (x1 ? (~x4 | x7) : (x4 | ~x7))) : (x2 | ((x1 | x4 | ~x7) & (~x4 | x7 | ~x1 | ~x3)));
  assign n1962 = (x0 | ~x1 | x3 | ~x4 | ~x7) & (~x0 | ~x3 | (x1 ? (~x4 | ~x7) : (x4 | x7)));
  assign n1963 = x1 & ((~x3 & x4 & ~x5 & ~x0 & x2) | (~x2 & ((x0 & x4 & (~x3 ^ x5)) | (~x4 & x5 & ~x0 & x3))));
  assign n1964 = ((x2 ? (x3 | ~x6) : (~x3 | x6)) | (x0 ? (x4 | x5) : (~x4 | ~x5))) & (~x3 | ~x6 | ((~x4 | ~x5 | ~x0 | ~x2) & (x0 | x2 | x4 | x5)));
  assign n1965 = ~x3 & x5 & (x0 ? (~x1 ^ ~x4) : (x1 & x4));
  assign n1966 = n1969 & ~n1967 & (x2 | ~x4 | ~n664 | n1968);
  assign n1967 = (~x0 ^ ~x3) & (x1 ? (~x4 & ~x5) : (x4 ^ x5));
  assign n1968 = (~x0 | ~x1 | x3 | x6) & (x0 | x1 | ~x3 | ~x6);
  assign n1969 = (~n992 | ~n848) & (~x3 | ~n1354 | ~n686);
  assign z146 = n1972 | ~n1975 | (~n1971 & ~n1981) | (~n705 & ~n1980);
  assign n1971 = x2 ? (~x5 | ~x7) : (x5 | x7);
  assign n1972 = ~x2 & (n1974 | (~x0 & ~n1973));
  assign n1973 = (x1 | ((x5 | x6 | ~x7 | x3 | x4) & (~x3 | ~x4 | ~x5 | ~x6 | x7))) & (~x1 | x3 | x4 | x5 | ~x6 | ~x7);
  assign n1974 = n595 & ((~x3 & x5 & ~x6 & (~x4 ^ ~x7)) | (x3 & x4 & ~x5 & x6 & ~x7));
  assign n1975 = ~n1977 & ~n1978 & (x0 | n1979) & (~n929 | n1976);
  assign n1976 = (x0 | x1 | x4 | ~x5 | ~x6 | ~x7) & (~x0 | x5 | x6 | (x1 ? (~x4 | x7) : (~x4 ^ ~x7)));
  assign n1977 = x4 & n321 & ((~x2 & ~x3 & x5 & ~x6) | (x3 & (x6 ? ~x5 : x2)));
  assign n1978 = ~n505 & ((~x0 & x2 & x3 & x5 & x6) | (x0 & ~x2 & ~x5 & (~x3 | ~x6)));
  assign n1979 = ((~x3 ^ x6) | ((x1 | x2 | ~x4 | x5) & (~x1 | ~x2 | x4 | ~x5))) & (~x1 | x2 | ((x5 | x6 | x3 | ~x4) & (~x5 | ~x6 | ~x3 | x4)));
  assign n1980 = (x5 & ((x2 & x3) | (~x0 & x6 & (x2 | x3)))) | (~x2 & ((~x5 & ~x6) | (~x3 & (~x5 | (x0 & ~x6))))) | (x0 & ~x5 & (x3 | ~x6));
  assign n1981 = (~x0 | x1 | ~x3 | x4 | ~x6) & (x0 | ((x4 | x6 | x1 | ~x3) & (~x1 | ~x4 | (~x3 ^ x6))));
  assign z147 = (~x0 & ~n1983) | (x3 & ~n1986) | (~x3 & ~n1987) | (x0 & ~n1988);
  assign n1983 = x2 ? n1985 : n1984;
  assign n1984 = x1 ? (x3 ? (~x4 | x6 | (x5 ^ x7)) : (~x6 | ((x5 | x7) & (x4 | ~x5 | ~x7)))) : ((~x3 | ~x4 | ~x5 | ~x6 | x7) & (x6 | ((~x5 | ~x7 | x3 | ~x4) & (x4 | (x3 ? (x5 ^ x7) : (x5 | ~x7))))));
  assign n1985 = (x5 | x6 | ~x7 | x1 | ~x3) & ((~x1 ^ ~x4) | ((x6 | x7 | ~x3 | ~x5) & (x3 | ~x6 | (~x5 ^ x7))));
  assign n1986 = (x0 | ((~x2 | x5 | ~x6) & (~x5 | ((x1 | x2 | ~x4 | x6) & (~x1 | (x2 ? (x4 | x6) : ~x6)))))) & (x2 | ((x4 | (x1 ? (x5 | (~x0 & x6)) : (~x5 | ~x6))) & (~x0 | ((x5 | x6) & (x1 | ~x5 | ~x6))))) & (~x0 | x1 | ~x2 | ~x5 | x6);
  assign n1987 = x2 ? ((~x0 | ((x5 | x6 | ~x1 | x4) & (x1 | ~x5 | ~x6))) & (x0 | ((~x5 | x6) & (x5 | ~x6 | x1 | ~x4))) & (~x5 | (x1 ? (x4 | ~x6) : (~x4 | x6)))) : ((x1 | ((~x4 | x5 | x6) & (x0 | ~x5 | ~x6))) & (~x0 | x5 | ~x6) & (x0 | ((~x4 | ~x5 | ~x6) & (~x1 | x5 | x6))));
  assign n1988 = (~n313 | n1990) & (n1591 | n1989) & (n564 | n852);
  assign n1989 = (~x1 | x2 | ~x4 | x5) & (x1 | x4 | (~x2 ^ ~x5));
  assign n1990 = (x1 | x2 | ~x5 | ~x6 | ~x7) & (~x1 | ~x2 | x5 | x6 | x7);
  assign z148 = ~n1992 | n2007 | (~n425 & ~n2010) | (~x0 & ~n2009);
  assign n1992 = n2003 & n1999 & ~n1998 & ~n1993 & ~n1996;
  assign n1993 = ~x3 & ((~x6 & ~n1994) | (n543 & n349 & ~n1995));
  assign n1994 = (x4 | x5 | ~x7 | x0 | x1 | x2) & (~x4 | ((~x0 | x7 | ((~x2 | x5) & (~x1 | x2 | ~x5))) & (x0 | ~x1 | ~x2 | ~x5 | ~x7)));
  assign n1995 = x2 ? (~x4 | ~x5) : (x4 | x5);
  assign n1996 = ~n1997 & (x2 ? n351 : n850);
  assign n1997 = (x0 | ~x1 | x3 | (~x6 ^ x7)) & (~x3 | ((~x0 | x1 | x6 | ~x7) & (x0 | (x1 ? (~x6 | ~x7) : (x6 | x7)))));
  assign n1998 = ~n437 & (x2 ? (n783 & n288) : (n595 & n361));
  assign n1999 = ~n2002 & (n2000 | n2001) & (~n543 | ~n373 | ~n459);
  assign n2000 = x1 ? (x4 | ~x6) : (~x4 | x6);
  assign n2001 = (x0 | ~x2 | x3 | ~x5) & (~x0 | x2 | ~x3 | x5);
  assign n2002 = ~x1 & x4 & ~x5 & x6 & (~x0 ^ ~x3);
  assign n2003 = ~n2005 & (n832 | n2004) & (~x5 | ~n865 | n2006);
  assign n2004 = (~x2 | ~x3 | x4 | x6 | ~x7) & (x2 | x3 | ~x4 | (~x6 ^ x7));
  assign n2005 = ~x6 & (x0 ? ((x4 & x5 & ~x1 & x3) | (~x4 & ~x5 & x1 & ~x3)) : ((~x1 & ~x3 & x4 & ~x5) | (x1 & x3 & ~x4 & x5)));
  assign n2006 = x1 ? (x2 ? (x4 | x6) : (~x4 | ~x6)) : (~x6 | (x2 ^ x4));
  assign n2007 = x3 & ((n1336 & n511) | (~x1 & ~n2008));
  assign n2008 = (x5 | x6 | ~x7 | ~x0 | x2 | x4) & (~x6 | x7 | ((x0 | x2 | ~x4 | ~x5) & (~x0 | x5 | (x2 ^ x4))));
  assign n2009 = x2 ? ((x1 | ~x3 | ~x4 | ~x5 | ~x6) & (~x1 | x5 | (x3 ? (~x4 | x6) : (x4 | ~x6)))) : ((x1 | ~x3 | x4 | ~x5 | ~x6) & (x6 | ((x4 | ~x5 | x1 | x3) & (~x1 | (x3 ? (x4 | x5) : (~x4 | ~x5))))));
  assign n2010 = x1 ? ((~x4 | ~x5 | x0 | ~x3) & (x2 | (x0 ? (x3 | (~x4 ^ x5)) : (~x3 | ~x4)))) : ((x0 | x2 | x3 | ~x4 | ~x5) & (x4 | (~x2 & x5) | (x0 ^ ~x3)));
  assign z149 = ~n2018 | (x1 ? (n2016 | n2017) : ~n2012);
  assign n2012 = (n1436 | n2014) & (~x0 | ~x3 | n2015) & (x0 | n2013);
  assign n2013 = (x4 | ((x2 | ~x3 | ~x5 | x6 | x7) & (~x6 | ((x2 | x3 | x5 | ~x7) & (~x2 | (x3 ? (x5 | x7) : (~x5 | ~x7))))))) & (~x3 | ~x4 | ~x7 | (x2 ? (x5 | ~x6) : (~x5 | x6)));
  assign n2014 = (x0 | ~x3 | ~x4 | x7) & (~x0 | (x3 ? (x4 | ~x7) : (~x4 | x7)));
  assign n2015 = (x2 | x4 | ~x5 | x6 | x7) & (~x2 | x5 | ~x6 | (~x4 ^ ~x7));
  assign n2016 = ~n307 & ((~x3 & n531 & n532) | (~x0 & x3 & ~n1436));
  assign n2017 = n1280 & ((x5 & x7 & x3 & ~x4) | (~x3 & ((~x5 & x7 & ~x0 & ~x4) | (x5 & ~x7 & x0 & x4))));
  assign n2018 = ~n2019 & n2020 & ~n2024 & (x7 | n2023);
  assign n2019 = ~x2 & ((~x1 & ~x3 & ~x4 & x5 & x7) | (~x5 & (x1 ? (x3 ? (~x4 & x7) : (x4 & ~x7)) : (x3 ? (~x4 & ~x7) : (x4 & x7)))));
  assign n2020 = ~n2022 & ~n2021 & (~x3 | ~x5 | ~n354 | n307);
  assign n2021 = x4 & (x1 ? (~x7 & ((~x2 & x3) | (~x0 & x2 & ~x3))) : (x7 & ((x2 & ~x3) | (x0 & ~x2 & x3))));
  assign n2022 = x2 & ~x4 & (x1 ? (x7 & (~x0 | ~x3)) : (~x3 & ~x7));
  assign n2023 = (x0 | x1 | x2 | x3 | ~x4 | ~x5) & ((x2 ? (~x3 | ~x4) : (x3 | x4)) | (x0 ? (x1 | x5) : (~x1 | ~x5)));
  assign n2024 = n1929 & ((~x0 & ~x1 & x3 & (x4 ^ x5)) | (x1 & ~x3 & (x0 ? (~x4 & ~x5) : (x4 & x5))));
  assign z150 = ~n2031 | (x2 ? ~n2028 : (x5 ? ~n2027 : ~n2026));
  assign n2026 = (x1 | ((x0 | ~x3 | x4 | x6 | x7) & (~x4 | ((x6 | ~x7 | x0 | ~x3) & (~x0 | (x3 ? (~x6 | ~x7) : (x6 | x7))))))) & (x0 | ~x1 | x3 | x4 | x7);
  assign n2027 = (x0 | x1 | x3 | x4 | ~x6 | ~x7) & (~x1 | ((~x3 | ((~x6 | x7 | ~x0 | x4) & (x0 | (x4 ? (~x6 | x7) : (x6 | ~x7))))) & (~x0 | x3 | x6 | (x4 ^ x7))));
  assign n2028 = (~x6 | n2029) & (x1 | x6 | n2030);
  assign n2029 = x0 ? (x1 | (x3 ? (x4 ? (x5 | x7) : (~x5 | ~x7)) : (~x4 | ~x5))) : ((~x4 | ~x5 | x7 | x1 | ~x3) & (~x1 | ((~x5 | ~x7 | x3 | x4) & (~x3 | ~x4 | x5 | x7))));
  assign n2030 = (~x0 | ~x3 | x5) & (~x5 | ((x0 | ~x3 | x4 | ~x7) & (x3 | (x0 ? (x4 ^ x7) : (~x4 | x7)))));
  assign n2031 = ~n2032 & ~n2034 & ~n2035 & ~n2036 & (~n269 | ~n1461);
  assign n2032 = x2 & ~n2033;
  assign n2033 = (x0 | ~x3 | ~x4 | ~x5 | ~x6 | ~x7) & (x6 | ((x0 | ~x3 | x4 | x5 | x7) & (x3 | ((~x0 | (x4 ? (x5 | x7) : (~x5 | ~x7))) & (~x5 | ~x7 | x0 | ~x4)))));
  assign n2034 = x0 & ((x2 & ~x3 & ~x4 & x5 & x6) | (~x2 & ((x3 & x5 & (x4 | ~x6)) | (~x5 & ((~x4 & x6) | (~x3 & (~x4 | x6)))))));
  assign n2035 = ~x0 & (x2 ? (x3 ? (x4 ? (~x5 & ~x6) : (x5 & x6)) : (x5 & (~x4 ^ x6))) : (x3 ? ((~x5 & x6) | (x4 & x5 & ~x6)) : (x4 & ~x5)));
  assign n2036 = ~n665 & ((x0 & ~x2 & ~x3 & x4 & ~x6) | (~x0 & ~x4 & (x2 ? (~x3 & x6) : (x3 & ~x6))));
  assign z151 = n2038 | n2042 | ~n2043 | ~n2047 | (~x2 & ~n2041);
  assign n2038 = ~x1 & ((x5 & ~n2039 & x0 & x3) | (~x3 & (~n2040 | (~x0 & ~x5 & ~n2039))));
  assign n2039 = (x2 | ~x4 | x6 | ~x7) & (~x2 | x4 | ~x6 | x7);
  assign n2040 = (x5 | x6 | ~x7 | x2 | x4) & (~x0 | ~x6 | ((x5 | ~x7 | x2 | ~x4) & (~x5 | x7 | ~x2 | x4)));
  assign n2041 = (~x4 | ((x0 | x1 | x3 | x5 | ~x6) & (~x1 | ~x5 | (x0 ? (~x3 ^ ~x6) : (~x3 | x6))))) & (~x0 | x3 | x4 | ~x6 | (x1 ^ ~x5));
  assign n2042 = (x3 ^ x6) & ((~x0 & (x1 ? (x4 ^ x5) : (x4 & x5))) | (~x4 & ~x5 & x0 & ~x1));
  assign n2043 = ~n2045 & ~n2046 & (n437 | n2044) & (~n686 | ~n552);
  assign n2044 = (~x3 | ((x0 | ~x1 | ~x2 | ~x4 | ~x5) & (~x0 | ((x1 | ~x4 | x5) & (x4 | ~x5 | ~x1 | x2))))) & (x0 | x3 | x4 | (x1 ^ ~x5));
  assign n2045 = ~n585 & ((~x0 & ~x1 & x2 & ~x3 & ~x5) | (x0 & x3 & (x1 ? (~x2 & ~x5) : x5)));
  assign n2046 = ~n390 & ((~x0 & ~x1 & ~x2 & x3 & ~x5) | (x0 & x2 & ~x3 & (~x1 ^ ~x5)));
  assign n2047 = ~n2049 & (n425 | n2048);
  assign n2048 = x0 ? (x3 | (x1 ? ((x4 | ~x5) & (x2 | ~x4 | x5)) : (~x4 | (~x2 ^ x5)))) : (x1 ? ((x4 | x5 | x2 | ~x3) & (~x4 | ~x5 | ~x2 | x3)) : (~x3 | x4 | (~x2 & ~x5)));
  assign n2049 = x1 & ((~x0 & ~n2050) | (n509 & n351 & x0 & n292));
  assign n2050 = ((x4 ^ x6) | ((x2 | x3 | ~x5 | ~x7) & (~x2 | ~x3 | x5 | x7))) & (~x5 | ~x6 | x7 | x2 | ~x3 | ~x4);
  assign z152 = n2052 | ~n2053 | n2057 | ~n2061 | (n345 & ~n2060);
  assign n2052 = ~n1054 & ((~x2 & (x1 ? (~x4 ^ x7) : (~x3 & (x4 ^ x7)))) | (~x4 & ~x7 & x1 & ~x3) | (~x1 & x2 & x3 & x4 & x7));
  assign n2053 = (n699 | n2056) & (n585 | n2055) & (~n1336 | ~n2054);
  assign n2054 = ~x7 & ~x5 & x3 & x4;
  assign n2055 = (x3 | ~x5 | ~x7 | ~x0 | x1 | ~x2) & (x2 | ((x5 | ((x0 | x1 | ~x3 | ~x7) & (~x0 | (x1 ? (~x3 | ~x7) : (x3 | x7))))) & (~x5 | x7 | x0 | ~x1)));
  assign n2056 = (~x1 | ((x0 | ~x2 | ~x5) & (x3 | x5 | ~x0 | x2))) & (~x0 | x1 | (x2 ? x5 : ~x3));
  assign n2057 = x2 & ((~x6 & ~n2059) | (~x0 & n367 & n2058));
  assign n2058 = ~x7 & x6 & x4 & ~x5;
  assign n2059 = (~x4 | ~x5 | x7 | ~x0 | x1 | x3) & (~x7 | (x1 ? (x3 | x5) : (~x3 | ~x5)) | (x0 ^ ~x4));
  assign n2060 = (x5 | ~x6 | ~x7 | x0 | x3 | ~x4) & (~x0 | ((x3 | x4 | x5 | ~x6 | ~x7) & (~x3 | ((~x6 | ~x7 | ~x4 | ~x5) & (x6 | x7 | x4 | x5)))));
  assign n2061 = (x0 | n2062) & (n589 | n2063);
  assign n2062 = (~x2 | ((x5 | x7 | ~x3 | x4) & (x1 | x3 | ~x4 | ~x7))) & (~x5 | ((~x1 | x2 | ~x3 | x4 | ~x7) & (x1 | ((x4 | x7) & (x2 | ~x4 | ~x7)))));
  assign n2063 = (x0 | x2 | ((x5 | x7 | x1 | ~x3) & (~x5 | ~x7 | ~x1 | x3))) & (~x2 | ((x0 | ~x1 | ~x3 | x5 | ~x7) & (x7 | ((x0 | x1 | x3 | x5) & (~x0 | (x1 ? (x3 | x5) : (~x3 | ~x5)))))));
  assign z153 = ~n2073 | ~n2071 | n2070 | n2065 | n2068;
  assign n2065 = ~x0 & ((n374 & ~n2067) | (~x7 & ~n2066));
  assign n2066 = (~x2 | ((~x4 | x5 | ~x6 | x1 | ~x3) & (~x5 | ((~x1 | ~x6 | (~x3 ^ x4)) & (x1 | x3 | x4 | x6))))) & (~x1 | x2 | x5 | (x3 ? (~x4 | x6) : (x4 | ~x6)));
  assign n2067 = (x1 | x2 | x3 | ~x4 | x5) & (~x2 | ((~x4 | ~x5 | x1 | ~x3) & (~x1 | x5 | (~x3 ^ x4))));
  assign n2068 = x0 & ((~x2 & ~n2069) | (n354 & ~n440 & ~n447));
  assign n2069 = (x5 | x6 | ~x7 | x1 | ~x3 | x4) & ((x3 ? (~x5 | ~x6) : (x5 | x6)) | (x1 ? (x4 | x7) : (~x4 | ~x7)));
  assign n2070 = ~x6 & n358 & ((n1354 & n321) | (~x0 & ~n1179));
  assign n2071 = ~n2072 & (n1085 | ((x0 | ~n1251) & (~n1906 | n1301)));
  assign n2072 = ~x2 & (x0 ? ((~x5 & x6 & ~x1 & ~x3) | (x5 & ~x6 & x1 & x3)) : (~x3 & x5 & (~x1 ^ x6)));
  assign n2073 = n2075 & ~n2077 & n2078 & (x2 | n2074);
  assign n2074 = x0 ? ((~x1 | ~x3 | x5 | ~x6 | ~x7) & (x1 | x3 | ~x5 | x6 | x7)) : (~x5 | ((~x1 | ~x3 | x6 | ~x7) & (x1 | x3 | ~x6 | x7)));
  assign n2075 = (~n1336 | ~n2076) & (~n686 | (~n1888 & (~n292 | ~n784)));
  assign n2076 = x5 & ~x3 & ~x4;
  assign n2077 = ~n362 & ((n1354 & n509) | (n654 & n929));
  assign n2078 = ~n2080 & (n2079 | n671);
  assign n2079 = x0 ? (x1 | ~x2) : (~x1 | x2);
  assign n2080 = (x1 ? (~x3 & x5) : (x3 & ~x5)) & (x0 ? (~x2 & x4) : (x2 & ~x4));
  assign z154 = n2082 | ~n2087 | (x6 ? (x7 ? ~n2085 : ~n2086) : (x7 ? ~n2086 : ~n2085));
  assign n2082 = ~x1 & ((n278 & ~n2084) | (x0 & ~n2083));
  assign n2083 = x2 ? (x7 | ((~x5 | ~x6 | ~x3 | x4) & (x5 | x6 | x3 | ~x4))) : (~x3 | ~x7 | (x4 ? (~x5 | ~x6) : (x5 | x6)));
  assign n2084 = x3 ? (x7 | (x4 ? (~x5 | ~x6) : (x5 | x6))) : (x4 | ~x7 | (x5 ^ x6));
  assign n2085 = x1 ? ((x2 | ((x4 | x5 | x0 | x3) & (~x0 | ~x3 | (x4 & x5)))) & (x0 | ~x2 | (x3 ? x4 : (~x4 | ~x5)))) : ((x3 | x4 | ~x0 | ~x2) & (x0 | ~x4 | (x2 ^ x3)));
  assign n2086 = (x2 | ((~x1 | ((x4 | x5 | ~x0 | x3) & (x0 | ~x3 | (~x4 ^ x5)))) & (~x0 | x1 | x3 | (~x4 & ~x5)))) & (x1 | ~x2 | (x0 ? (~x3 | ~x4) : (x3 | (x4 & x5))));
  assign n2087 = ~n2088 & n2090 & (x3 ? n2092 : n2091);
  assign n2088 = x1 & (x0 ? (n509 & n284) : ~n2089);
  assign n2089 = (x5 | ~x6 | ~x7 | ~x2 | x3 | ~x4) & (x2 | ((x3 | x4 | ~x5 | x6 | x7) & (~x3 | ((x6 | ~x7 | ~x4 | ~x5) & (~x6 | x7 | x4 | x5)))));
  assign n2090 = x1 ? ((x0 | ~x2 | ~x3 | ~x4 | ~x6) & (x3 | (x0 ? (x2 ? (x4 | ~x6) : (~x4 | x6)) : (x2 ? (x4 | x6) : (~x4 | ~x6))))) : (x0 ? (~x4 | (x2 ? (x3 | ~x6) : (~x3 | x6))) : (~x3 | x4 | (~x2 ^ x6)));
  assign n2091 = (x2 | x4 | (x0 ? (x1 ? (~x5 | x6) : (x5 | ~x6)) : (~x5 | (x1 ^ x6)))) & (x0 | ~x2 | ~x4 | x6 | (x1 ^ ~x5));
  assign n2092 = (x4 | x5 | ~x6 | ~x0 | x1 | ~x2) & (x2 | ((x0 | x1 | ~x4 | x5 | ~x6) & (~x0 | ~x5 | (x1 ? (~x4 | ~x6) : (x4 | x6)))));
  assign z155 = (~x4 & ~n2094) | (~x3 & ~n2100) | ~n2097 | (x4 & ~n2101);
  assign n2094 = (x1 | n2095) & (~n444 | n2096);
  assign n2095 = (~x0 | ~x2 | ~x3 | ~x5 | ~x6 | ~x7) & (x2 | ((x5 | ((~x3 | ~x6 | x7) & (x0 | ((~x6 | x7) & (~x3 | x6 | ~x7))))) & (x0 | x3 | ~x5 | (x6 ^ x7))));
  assign n2096 = (x3 | ~x5 | ~x6 | x7) & (~x3 | x5 | (x6 ^ x7));
  assign n2097 = (~n509 | n2099) & (~x3 | n2098) & (x3 | n515 | n891);
  assign n2098 = x2 ? ((x1 | (x4 ^ x7)) & (x0 | ~x1 | (~x4 ^ x7))) : ((x0 | x1 | ~x4 | x7) & (~x0 | ~x1 | x4 | ~x7));
  assign n2099 = x1 ? (~x7 | ((~x4 | x5) & (x0 | x4 | ~x5))) : (x7 | ((x4 | ~x5) & (~x0 | ~x4 | x5)));
  assign n2100 = (((~x0 | x1 | x2 | x4) & (~x2 | ~x4 | x0 | ~x1)) | (x5 ^ x7)) & (~x1 | x2 | x4 | ((x5 | ~x7) & (~x0 | ~x5 | x7))) & (x1 | ~x2 | ~x4 | ((~x5 | x7) & (x0 | x5 | ~x7)));
  assign n2101 = (~x6 | ((x7 | n2103) & (x0 | ~x7 | n2102))) & ~n2104 & (x6 | ((~x7 | n2103) & (~x0 | x7 | n2102)));
  assign n2102 = (~x1 | ~x2 | x3 | x5) & (x1 | x2 | ~x3 | ~x5);
  assign n2103 = (~x0 | x1 | ~x2 | x3 | x5) & (x0 | ~x1 | x2 | ~x3 | ~x5);
  assign n2104 = ~n891 & n532 & x3 & n531;
  assign z156 = n2110 | ~n2111 | (~x1 & ~n2106) | (x6 & ~n2107);
  assign n2106 = (x3 | ((~x0 | ((~x2 | x5 | ~x6) & (~x5 | x6 | x2 | x4))) & (x5 | ((~x2 | x4 | ~x6) & (x0 | x2 | ~x4))))) & (x0 | ((x4 | ~x5 | x2 | ~x3) & (~x2 | x6 | ((x4 | x5) & (~x3 | ~x4 | ~x5)))));
  assign n2107 = ~n2109 & (x7 | n2108) & (~x5 | ~x7 | ~n373 | ~n459);
  assign n2108 = (~x3 | ~x4 | ~x5 | x0 | x1 | ~x2) & (x2 | ((x3 | ~x4 | x5 | x0 | ~x1) & (~x0 | ((~x4 | x5 | x1 | x3) & (x4 | ~x5 | ~x1 | ~x3)))));
  assign n2109 = ~n2102 & (x0 ? (~x4 & ~x7) : (x4 & x7));
  assign n2110 = ~n1158 & ((x2 & ~x3 & ~x4 & ~x5 & ~x6) | (~x2 & (x3 ? (x4 ? (x5 & x6) : (x5 ^ x6)) : (x4 ? (~x5 & ~x6) : (x5 & x6)))));
  assign n2111 = ~n2114 & ~n2115 & (x6 | (~n2113 & (x4 | n2112)));
  assign n2112 = (~x3 | x5 | ((x0 | ~x1 | ~x2 | x7) & (~x0 | x1 | (~x2 ^ x7)))) & (x0 | x3 | ~x5 | ((~x2 | x7) & (~x1 | x2 | ~x7)));
  assign n2113 = n361 & ((~x0 & ~x1 & ~x2 & ~x5 & ~x7) | (x0 & x5 & (x1 ? (~x2 & x7) : (x2 & ~x7))));
  assign n2114 = ~n1231 & ((~x0 & (n1230 | (~x1 & x6 & n748))) | (~x1 & n1230) | (x0 & x1 & ~x6 & n748));
  assign n2115 = n349 & ((~x2 & x3 & ~x4 & x5 & x6) | (x2 & ((x3 & x4 & x5 & ~x6) | (~x3 & ~x4 & ~x5 & x6))));
  assign z157 = (~x1 & ~n2117) | (x1 & ~n2119) | ~n2123 | (~n392 & ~n2122);
  assign n2117 = (~n342 | ~n464) & (x3 | n2118);
  assign n2118 = (x5 | ~x6 | ~x7 | ~x0 | x2 | ~x4) & (x0 | ((x2 | x4 | x5 | ~x6 | x7) & (x6 | ((x2 | x4 | x5 | ~x7) & (~x2 | (x4 ? (x5 | x7) : (~x5 | ~x7)))))));
  assign n2119 = (x0 | n2121) & (n2120 | ((~x0 | x4 | x5 | ~x6) & (x0 | (x4 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n2120 = x2 ? (x3 | ~x7) : (~x3 | x7);
  assign n2121 = (~x2 | ~x3 | ~x4 | x5 | ~x6 | x7) & (x2 | x3 | ((x6 | ~x7 | x4 | ~x5) & (~x4 | ~x6 | (~x5 ^ x7))));
  assign n2122 = (x6 | ((~x0 | ~x4 | ~x5 | (x1 ^ ~x2)) & (x5 | (x0 ? (x1 | x4) : (x1 ? (~x2 | x4) : (x2 | ~x4)))))) & (~x5 | ~x6 | (x0 ? (x4 | (x1 & x2)) : (x1 | ~x4)));
  assign n2123 = n2125 & (n864 | n2124) & (~n451 | ~n313 | ~n460);
  assign n2124 = x3 ? ((x5 | ~x6 | x0 | x4) & (~x4 | ((x5 | x6) & (~x0 | ~x5 | ~x6)))) : (x0 ? (x4 ? (x5 | ~x6) : (~x5 | x6)) : (x4 ? (~x5 | x6) : (x5 ^ x6)));
  assign n2125 = (~x3 | n2127) & (n2126 | (~x1 ^ ~x2));
  assign n2126 = (~x0 | x3 | x4 | ~x5 | x6) & (x0 | ((x5 | ~x6 | ~x3 | x4) & (x3 | ~x5 | (~x4 ^ x6))));
  assign n2127 = x4 ? ((x1 | (x0 ? (x2 | (x5 ^ x6)) : (x5 | ~x6))) & (x0 | ~x1 | ((~x5 | ~x6) & (~x2 | x5 | x6)))) : ((x0 | x1 | x2 | ~x5 | x6) & (~x0 | x5 | (x1 ? (x2 | x6) : ~x6)));
  assign z158 = ~n2133 | (~x4 & ~n2129) | (~x1 & ~n2132);
  assign n2129 = n2131 & (~x1 | n2130) & (x3 | n665 | ~n1192);
  assign n2130 = (~x5 | ((~x0 | ~x2 | x3 | ~x6 | ~x7) & (x0 | x7 | (x2 ? (~x3 | x6) : (x3 | ~x6))))) & (~x0 | x5 | ((~x6 | ~x7 | x2 | ~x3) & (x6 | x7 | ~x2 | x3)));
  assign n2131 = x5 | x7 | (x3 ? ~n317 : (x6 | ~n686));
  assign n2132 = (~x6 | (x0 ? (~x4 | ((~x5 | x7) & (~x2 | x5 | ~x7))) : (x4 | (~x5 ^ x7)))) & (x5 | x6 | ~x7 | (x0 ^ ~x4));
  assign n2133 = ~n2134 & ~n2136 & (~n369 | n2135) & (~x1 | n2137);
  assign n2134 = ~n425 & ((x5 & (~x1 | ~x2) & (~x0 ^ ~x4)) | (x4 & ~x5 & (x0 ? (~x1 & ~x2) : x1)));
  assign n2135 = ((x2 ? (x3 | x6) : (~x3 | ~x6)) | (x0 ? (x1 | x5) : (~x1 | ~x5))) & (~x3 | x5 | x6 | x0 | x1 | ~x2) & (x3 | ~x5 | ~x6 | ~x0 | ~x1 | x2);
  assign n2136 = ~n434 & ((x1 & (x0 ? (~x2 & x4) : ~x4)) | (~x0 & x2 & ~x4) | (~x1 & ((~x3 & x4 & ~x0 & ~x2) | (x0 & (~x2 ^ x4)))));
  assign n2137 = (~x0 | x2 | x4 | x5 | x6) & (x0 | ((x5 | x6 | ~x7 | x2 | ~x4) & (~x2 | ((~x4 | ~x5 | ~x6) & (x6 | ~x7 | x4 | x5)))));
  assign z159 = n2139 | n2143 | n2146 | n2147 | (~n425 & ~n2145);
  assign n2139 = ~x6 & (n2141 | ~n2142 | (x0 & ~n2140));
  assign n2140 = (x1 | ~x2 | x3 | x4 | ~x5 | ~x7) & (x5 | ((x1 | x2 | ~x3 | x4 | ~x7) & (x7 | ((~x3 | ~x4 | x1 | ~x2) & (~x1 | x3 | (~x2 ^ ~x4))))));
  assign n2141 = ~x5 & ((~x1 & ~x2 & ~x3 & x7) | (~x0 & x2 & (x1 ? x7 : (x3 & ~x7))));
  assign n2142 = ~x3 | ~x5 | ((x7 | ~n992) & (~x4 | ~x7 | ~n317));
  assign n2143 = x6 & ((x5 & ~n2144) | (n870 & n361 & n992));
  assign n2144 = (x0 | ~x1 | ~x2 | x7) & (x1 | ((~x0 | ((~x4 | ~x7 | ~x2 | ~x3) & (x2 | x3 | x7))) & (x4 | ((x2 | x3 | x7) & (~x3 | ~x7 | x0 | ~x2)))));
  assign n2145 = (x2 & ((x0 & ~x5 & (x3 | x4)) | (x3 & (x4 | (~x0 & x5))))) | (x1 & x5) | (~x5 & (~x1 | (~x3 & ~x4 & x0 & ~x2)));
  assign n2146 = ~n437 & ~n847 & ((x0 & x2 & ~x3 & ~x4) | (~x2 & x3 & (~x0 | x4)));
  assign n2147 = ~n434 & (x1 ? (~x2 & (~x3 | (x0 & ~x4))) : (x2 & (~x0 | x3 | x4)));
  assign z160 = ~n2151 | (~n617 & ~n2149) | (x3 & ~n2150);
  assign n2149 = (x0 | ((~x1 | x3 | x7) & (x1 | ~x3 | ~x4 | ~x5 | ~x7))) & (~x0 | ((x1 | x7 | (x3 & (x4 | x5))) & (x3 | x4 | (~x1 & x5)))) & (x3 | x7 | ((x4 | ~x5) & (x1 | ~x4 | x5)));
  assign n2150 = x0 ? (x7 | ((~x4 | x6 | x1 | ~x2) & (x2 | ((~x4 | ~x6) & (~x1 | x4 | x6))))) : ((x1 | x2 | x4 | ~x6 | ~x7) & (~x1 | ~x2 | ~x4 | x6 | x7));
  assign n2151 = n2158 & ~n2157 & ~n2156 & ~n2152 & ~n2155;
  assign n2152 = ~x4 & ((n531 & n532 & ~n2154) | (x2 & ~n2153));
  assign n2153 = (~x5 | x6 | ~x7 | ~x0 | x1 | x3) & (x0 | x7 | ((~x1 | ~x3 | ~x5 | x6) & (x1 | x3 | x5 | ~x6)));
  assign n2154 = x1 ? (x3 | ~x7) : (~x3 | x7);
  assign n2155 = (x2 ^ x6) & ((~x1 & x3 & (x0 ^ ~x7)) | (~x0 & x7 & (x1 | ~x3)));
  assign n2156 = x4 & n865 & (x1 ? (~x2 & ~n425) : (x2 & n292));
  assign n2157 = ~x2 & x6 & ((x0 & x7 & (x1 ^ ~x3)) | (x3 & ~x7 & ~x0 & x1));
  assign n2158 = ~n2159 & (x2 | ~x4 | ~x6 | ~n783 | n1367);
  assign n2159 = x7 & ~x6 & x3 & x2 & ~x0 & ~x1;
  assign z161 = (~x4 & ~n2161) | (x4 & ~n2163) | ~n2166 | (~x0 & ~n2165);
  assign n2161 = (~x0 | n2162) & (~n400 | (x3 ? n437 : ~n372));
  assign n2162 = (x3 | ((~x1 | x2 | ~x5 | ~x6 | ~x7) & (x1 | ((~x6 | ~x7 | x2 | x5) & (x6 | x7 | ~x2 | ~x5))))) & (x1 | ~x2 | ~x3 | ~x5 | (~x6 ^ x7));
  assign n2163 = (x3 | x5 | ~n372 | ~n524) & (~x5 | ~n783 | n2164);
  assign n2164 = (~x3 | (x2 ? (~x6 | ~x7) : (x6 | x7))) & (~x2 | x3 | (~x6 ^ x7));
  assign n2165 = (~x1 | ~x2 | ~x3 | x4 | ~x5 | x7) & (x1 | ~x4 | ((x3 | x5 | ~x7) & (x2 | (x3 ? (x5 ^ x7) : (~x5 | x7)))));
  assign n2166 = ~n2167 & ~n2168 & ~n2169 & (x4 | n392 | ~n1924);
  assign n2167 = x2 & ((x0 & x1 & ~x3 & ~x4 & ~x7) | (~x0 & ((x4 & ~x7 & ~x1 & x3) | (~x4 & x7 & x1 & ~x3))));
  assign n2168 = (~x0 | (x4 & (~x1 | ~x2))) & (~x3 | ~x7) & (x3 | x7) & (~x1 | ~x2 | x4) & (x0 | x1 | ~x4);
  assign n2169 = ~x4 & n321 & (x3 ? ((~x5 & x7) | (~x2 & x5 & ~x7)) : (~x5 ^ x7));
  assign z162 = x4 ? (n2173 | ~n2174) : (x3 ? ~n2172 : ~n2171);
  assign n2171 = ((x2 & ~x6) | (x0 ? (x1 | ~x5) : ~x1)) & (~x1 | ((~x0 | ~x2 | x5 | x6 | x7) & (~x6 | ~x7 | x2 | ~x5))) & (~x2 | x6 | ((x0 | (x1 & ~x5)) & (x1 | ~x5 | ~x7))) & (x5 | ((x1 | x2 | ~x6 | ~x7) & (x0 | (~x6 & ~x7))));
  assign n2172 = (x1 & (x0 | (x2 & ~x5 & ~x6))) | (x0 & (~x5 | (x2 & ~x6))) | (~x0 & ~x1 & x5 & ((x6 & x7) | (~x2 & (x6 | x7))));
  assign n2173 = x3 & ~n617 & ((x0 & ~x1 & x5 & ~x7) | (~x0 & (x1 ? (~x5 & ~x7) : (x5 & x7))));
  assign n2174 = x1 ? ((~x0 | x2) & (x5 | x6 | x0 | ~x2)) : (x0 ? (x5 & (~x2 | x6)) : (~x5 | ((x3 | ~x6) & (x2 | (x3 & ~x6)))));
  assign z163 = n2176 | n2179 | n2182 | ~n2184 | (~x0 & ~n2178);
  assign n2176 = ~x6 & ((~x1 & ~n2177) | (n664 & n361 & n1336));
  assign n2177 = (~x0 | ((~x2 | x3 | x4 | ~x5 | ~x7) & (~x4 | x5 | x7 | x2 | ~x3))) & (x2 | ~x3 | ~x5 | ~x7 | (x0 & ~x4));
  assign n2178 = (~x3 | ((~x1 | ~x2 | ~x5 | x6) & (x4 | ((x5 | (~x1 ^ (x2 & ~x6))) & (x1 | x2 | ~x5 | ~x6))))) & (~x1 | ~x2 | ~x4 | ((~x5 | x6) & (x3 | x5 | ~x6)));
  assign n2179 = x6 & (x0 ? ~n2180 : ~n2181);
  assign n2180 = (x4 | x5 | ~x7 | x1 | x2 | x3) & (((~x1 | x2 | x3 | x4) & (~x3 | ~x4 | x1 | ~x2)) | (x5 ^ x7));
  assign n2181 = (x1 | ~x2 | ~x3 | ~x5 | ~x7) & (~x1 | x4 | x7 | (x2 ? (~x3 | ~x5) : (x3 | x5)));
  assign n2182 = ~n2183 & (x1 ? (~x5 ^ ~x7) : (~x5 & ~x7));
  assign n2183 = (x4 | x6 | ~x2 | x3) & (x0 | ~x3 | ~x4 | (~x2 ^ ~x6));
  assign n2184 = ~n2186 & ~n2187 & (~n1336 | ~n552) & (n2185 | n2188);
  assign n2185 = (x3 | ~x4) & (~x0 | ~x3 | x4);
  assign n2186 = (x1 ^ x5) & ((~x2 & (x3 ? (x4 & x6) : (~x4 & ~x6))) | (~x4 & x6 & x2 & ~x3));
  assign n2187 = ~x1 & ((~x2 & ~x3 & ~x4 & x5 & x6) | (x2 & x3 & x4 & ~x5 & ~x6));
  assign n2188 = (x1 | ((~x5 | ~x6) & (~x2 | x5 | x6))) & (x2 | (x1 ^ ~x5));
  assign z164 = n2190 | ~n2193 | n2199 | (x0 & ~n2200);
  assign n2190 = ~x2 & ((~x5 & ~n2191) | (n2192 & (~x1 | x7)));
  assign n2191 = x0 ? ((x1 | x3 | x4 | ~x6 | ~x7) & (~x1 | ~x3 | ~x4 | x6 | x7)) : (x4 | ((~x6 | ~x7 | ~x1 | x3) & (~x3 | x6 | (x1 & ~x7))));
  assign n2192 = ~x6 & x5 & ~x4 & ~x0 & ~x3;
  assign n2193 = n2196 & (n437 | n2194) & (x4 | ~n487 | n2195);
  assign n2194 = x2 ? (x3 | x4 | (~x0 & ~x1 & x5)) : (~x3 | (~x4 & (x0 | ~x5)));
  assign n2195 = (~x3 | x5 | ~x6 | x7) & (~x5 | ((x3 | ~x6 | ~x7) & (x1 | (x3 ? (x6 | x7) : ~x6))));
  assign n2196 = ~n2197 & ~n2198 & (~x4 | ~n374 | (~n342 & ~n459));
  assign n2197 = (x0 ? (~x2 & ~x6) : (x2 & x6)) & (x3 ? (~x4 & x7) : x4);
  assign n2198 = ~x7 & ~x6 & ~x4 & ~x2 & ~x0 & x1;
  assign n2199 = ~x6 & ((x0 & ~x2 & ~x4 & ~x7) | (~x0 & x4 & (x2 ? (x3 & ~x7) : ~x3)));
  assign n2200 = (~x1 | x2 | x3 | x4 | ~x6 | ~x7) & (x1 | ~x2 | ((~x6 | x7 | x3 | ~x4) & (~x3 | (x4 ? (x6 | x7) : ~x6))));
  assign z165 = n2203 | ~n2204 | n2207 | (~x2 & ~n2202) | n2208;
  assign n2202 = (x3 | (x0 ? ((x5 | ~x7 | x1 | x4) & (~x5 | x7 | ~x1 | ~x4)) : (x4 | (x1 ? (x5 | ~x7) : (~x5 | x7))))) & (x0 | ~x3 | x4 | (x5 ^ x7));
  assign n2203 = (~x1 ^ ~x2) & ((x0 & ~x4 & (x3 ^ x7)) | (x4 & ((x3 & x7) | (~x0 & ~x3 & ~x7))));
  assign n2204 = ~n2206 & ~n2205 & (~n345 | ~n370 | n520 | n1054);
  assign n2205 = x0 & ((x1 & x2 & ~x3 & ~x4 & x7) | (~x1 & ((~x3 & x4 & ~x7) | (~x2 & x3 & (~x4 ^ x7)))));
  assign n2206 = ~x0 & x4 & (~x3 ^ x7) & (~x1 ^ x2);
  assign n2207 = ~x4 & n487 & ((~x5 & ~n406) | (~x1 & x5 & ~n392));
  assign n2208 = x1 & (n2209 | (x7 & n850 & n487 & ~n520));
  assign n2209 = ~x7 & ~n798 & ((n351 & n532) | (~x0 & n850));
  assign z166 = n1945 | n2212 | (x2 ? ~n2214 : ~n2211);
  assign n2211 = (x0 & ((x1 & ((x4 & x7) | (~x6 & ~x7 & ~x4 & ~x5))) | (x4 & (x7 ? (~x5 | ~x6) : x5)))) | (x4 & ((x1 & (x5 ? (~x6 & ~x7) : x7)) | (~x5 & (x7 ? ~x6 : (~x0 | ~x1 | x6))))) | (~x4 & ((x6 & x7 & ~x1 & x5) | (~x0 & ((x5 & (x6 | x7)) | (~x1 & (~x6 ^ x7))))));
  assign n2212 = ~x4 & ((~x5 & ~n2213) | (x2 & n294 & n595));
  assign n2213 = (x0 | x1 | x2 | ~x3 | x6 | x7) & (~x0 | ~x1 | x3 | (~x2 ^ (~x6 & ~x7)));
  assign n2214 = (x1 | (x0 ? x4 : (~x4 | ~x5))) & (x0 | (x4 ? (~x5 | ~x6) : (x5 & (~x1 | x6))));
  assign z167 = n2218 | ~n2219 | (~x3 & (n2217 | (~x5 & ~n2216)));
  assign n2216 = (x6 | ((x0 | ((x1 | x2 | ~x4 | x7) & (~x1 | ~x2 | x4 | ~x7))) & (~x0 | ~x1 | x2 | ~x4 | x7))) & (~x0 | x1 | x4 | ~x6 | (~x2 ^ ~x7));
  assign n2217 = n850 & n595 & (x2 ^ (~x6 & ~x7));
  assign n2218 = ~n1826 & ((~x1 & ((~x6 & x7 & ~x0 & ~x5) | (x0 & x5 & (~x6 | ~x7)))) | (~x0 & ((~x5 & x6 & ~x7) | (x1 & (x5 ? (~x6 & ~x7) : x6)))));
  assign n2219 = ~n2221 & ~n2222 & n2223 & ((x2 & x3) | n2220 | (~x2 & ~x3));
  assign n2220 = x0 ? ((x6 | x7 | ~x1 | x5) & (x1 | ~x5 | (x6 & x7))) : ((~x1 | (x5 ? (x6 | x7) : ~x6)) & (x5 | (x6 ? x7 : x1)));
  assign n2221 = x7 & (((~x2 ^ x5) & (x0 ? (~x1 & x6) : (x1 & ~x6))) | (x0 & x1 & ~x2 & x5) | (~x0 & ~x1 & x2 & ~x5 & x6));
  assign n2222 = n783 & ((n358 & n612) | (n357 & n611));
  assign n2223 = (~n1336 | ~n781) & (~n509 | ~n850 | ~n783 | ~n374);
  assign z168 = n2227 | n2228 | n2230 | ~n2231 | (x5 & ~n2225);
  assign n2225 = (~n288 | ~n992 | x6 | ~x7) & (x1 | ~x6 | n2226);
  assign n2226 = (x0 | x2 | ~x3 | ~x4 | ~x7) & (~x0 | x3 | x4 | (~x2 ^ ~x7));
  assign n2227 = x2 & ((~x0 & ~x1 & x6) | ((x3 | x4) & ((~x1 & x6) | (~x0 & x1 & ~x6))));
  assign n2228 = ~n2229 & (x1 ? (~x6 ^ x7) : (~x6 ^ ~x7));
  assign n2229 = (x0 & ~x2 & ~x3 & ~x4) | (x2 & (~x0 | x3 | x4));
  assign n2230 = ~x7 & n312 & n865 & (x1 ? n1230 : n748);
  assign n2231 = x3 | x4 | (x6 ? ~n1336 : n2232);
  assign n2232 = (~x0 | x1 | x2 | ~x7) & (x0 | ~x1 | ~x2 | x7);
  assign z169 = n2234 | ~n2235 | n2239 | (~n425 & ~n2240);
  assign n2234 = n288 & ((~x0 & x1 & x2 & x5 & x7) | (~x1 & ((~x2 & x5 & ~x7) | (x0 & ~x5 & (x2 ^ x7)))));
  assign n2235 = ~n2236 & n2238 & (x7 | ~n784 | n2237);
  assign n2236 = x2 & ~x3 & ((x4 & x7 & ~x0 & x1) | (x0 & (x1 ? (~x4 & ~x7) : (x4 & x7))));
  assign n2237 = (x0 | x1 | x2 | x4 | ~x6) & (~x0 | ~x1 | ~x2 | ~x4 | x6);
  assign n2238 = (x0 | ((~x7 | ((~x2 | ~x3) & (x1 | (~x2 & ~n2054)))) & (x2 | x7 | (~x1 & ~n2054)))) & (~x3 | ((x1 | ~x2 | ~x7) & (~x0 | x2 | x7)));
  assign n2239 = ~x2 & ((~x0 & ~x1 & x3 & ~x4 & ~x7) | (~x3 & ((~x1 & x4 & ~x7) | (x0 & ((x4 & ~x7) | (x1 & ~x4 & x7))))));
  assign n2240 = (x0 | ((x1 | x2 | ~x3 | ~x4 | ~x5) & (~x1 | ~x2 | x3 | x4 | x5))) & (x3 | x4 | ~x5 | ~x0 | x1 | ~x2);
  assign z170 = n2242 | n2245 | (x0 ? ~n2243 : ~n2244);
  assign n2242 = n269 & n1415;
  assign n2243 = (x1 & (x2 | (~x3 & ~x4))) | (x2 & (x3 ? (x5 & x6) : (~x4 & ~x6))) | (~x3 & ~x4 & ~x5) | (x3 & (x4 | (~x1 & ~x2 & x5)));
  assign n2244 = (x1 | ((~x2 | x3 | x6) & (x2 | ~x3 | ~x4 | ~x5 | ~x6))) & (~x2 | x6 | ((x3 | ~x5) & (x4 | x5 | ~x1 | ~x3))) & (x3 | ((~x1 | (x2 & ~x6)) & (x4 | ~x5) & (x5 | (~x4 & ~x6))));
  assign n2245 = ~x7 & ((n1336 & n552) | (~n617 & ~n2246));
  assign n2246 = (~x0 | x1 | ~x3 | x4 | ~x5) & (x0 | ((~x1 | ~x3 | x4 | x5) & (~x4 | ~x5 | x1 | x3)));
  assign z171 = ~n2249 | ~n2253 | ((x0 | ~x7) & ~n2248 & (~x0 | x7));
  assign n2248 = (x1 | x4 | ~x5 | (~x2 ^ ~x6)) & (~x1 | x2 | ~x4 | x5 | x6);
  assign n2249 = n2250 & ~n2251 & (~n870 | ~n1602 | n2252);
  assign n2250 = x4 ? ((~x1 | ((~x0 | x2 | ~x5) & (x5 | x6 | x0 | ~x2))) & (~x0 | x1 | (x5 & (~x2 | x6)))) : ((x0 | ((~x1 | (~x5 & (x2 | ~x6))) & (~x2 | (x5 ? x6 : x1)))) & (~x0 | x1 | x2 | ~x5 | ~x6));
  assign n2251 = ~x2 & x6 & ((x0 & x1 & x4 & ~x5) | (~x0 & ~x1 & (~x4 ^ x5)));
  assign n2252 = (x2 | x6) & (~x1 | ~x2 | ~x6);
  assign n2253 = (n617 | n2254) & (~n616 | n2255);
  assign n2254 = (x0 | ~x1 | x3 | x4 | x5 | x7) & (x1 | ~x5 | (x0 ? (x7 | (x3 ^ x4)) : (~x7 | (~x3 ^ x4))));
  assign n2255 = (x0 | x1 | x2 | ~x3 | x4 | x6) & (~x1 | ((x0 | ~x2 | ~x3 | ~x4 | ~x6) & (~x0 | x3 | x6 | (~x2 ^ x4))));
  assign z172 = ~n2262 | (x1 ? ~n2257 : (n2260 | (~x4 & ~n2261)));
  assign n2257 = (~n1050 | n2259) & (~n1029 | ~n1018) & (n665 | n2258);
  assign n2258 = (x0 | ~x2 | ~x3 | x4 | ~x6) & (x6 | (x0 ? (x2 ? (x3 | x4) : (~x3 | ~x4)) : (x2 | (~x3 ^ x4))));
  assign n2259 = (x2 | ~x3 | x5 | x6 | ~x7) & (~x2 | ~x6 | (x3 ? (x5 | ~x7) : (~x5 | x7)));
  assign n2260 = ~n440 & (x0 ? (x3 & (x2 ? (x4 & x6) : ~x6)) : (~x3 & x4 & (x2 ^ ~x6)));
  assign n2261 = (~x2 | (x0 ? ((~x6 | ~x7 | ~x3 | ~x5) & (x6 | x7 | x3 | x5)) : (~x6 | (x3 ? (x5 | x7) : (~x5 | ~x7))))) & (x0 | x2 | x6 | (x3 ? (x5 | x7) : (~x5 | ~x7)));
  assign n2262 = ~n2264 & ~n2265 & ~n2266 & (~x4 | n2263);
  assign n2263 = (x5 | (x0 ? (x3 | (x1 ? (x2 | ~x6) : (~x2 | x6))) : (x1 | ~x3 | (~x2 ^ ~x6)))) & (x0 | ~x1 | ~x3 | ~x5 | (~x2 ^ ~x6));
  assign n2264 = x2 & ((~x0 & (x1 ? ((~x3 & ~x5 & x6) | (x5 & ~x6)) : (~x5 & ~x6))) | (~x1 & ((x3 & ~x5 & ~x6) | (x5 & x6 & x0 & ~x3))));
  assign n2265 = ~x2 & ((x0 & ~x3 & (x1 ? (~x5 & ~x6) : x5)) | (x6 & (x1 ? (~x5 & (~x0 | x3)) : x5)));
  assign n2266 = ~x5 & n452 & ((~x0 & ~x2 & ~x3 & ~x6) | (x0 & (x2 ? (~x3 & x6) : (x3 & ~x6))));
  assign z173 = ~n2272 | (x6 & ~n2271) | (~x0 & (n2268 | n2269));
  assign n2268 = ~n505 & ((x3 & ~x5 & n374) | (x2 & (x3 ? n372 : (x5 & n374))));
  assign n2269 = x2 & ((~n425 & ~n2270) | (x1 & n313 & n1048));
  assign n2270 = x1 ? (~x3 | x4) : (x3 | ~x4);
  assign n2271 = (x1 | x4 | ((x0 | x2 | ~x3 | ~x5) & (~x2 | (x0 ? (~x3 ^ x5) : (x3 | x5))))) & (x0 | ~x1 | ~x4 | (x2 ? (x3 | x5) : (~x3 | ~x5)));
  assign n2272 = n2276 & (n437 | n2273) & (~x0 | (~n2274 & ~n2275));
  assign n2273 = (~x0 | (x2 ? (x3 | x4 | (~x1 & x5)) : (~x3 | (x1 & ~x4)))) & (x2 | ((~x3 | (x1 ? (x4 ? x5 : x0) : (x4 | x5))) & (x0 | x3 | (x1 & ~x4))));
  assign n2274 = ~n425 & ((~x3 & ~x4 & ~x5 & n542) | (x3 & n354 & (x4 | x5)));
  assign n2275 = n288 & ((n542 & n1048) | (~x5 & n354 & n374));
  assign n2276 = x3 ? ((x0 | x1 | ~x4 | (~x2 ^ x6)) & (~x0 | ~x1 | x2 | x4 | x6)) : (x0 ? ((x2 | ~x4 | x6) & (x1 | (x2 ? (~x4 | ~x6) : x6))) : (~x1 | x4 | (~x2 ^ ~x6)));
  assign z174 = ~n2284 | n2283 | n2281 | n2280 | n2278 | n2279;
  assign n2278 = n783 & n548 & ((~x2 & x3 & ~x5 & x7) | (x2 & x5 & (x3 ^ ~x7)));
  assign n2279 = ~x0 & ((x4 & x7 & ~x2 & ~x3) | (~x1 & ((~x2 & ~x3 & x7) | (x4 & ~x7 & x2 & x3))));
  assign n2280 = ~x0 & ~n505 & ((x2 & ~x3 & (~x5 ^ x7)) | (x3 & (x2 ? (~x5 & x7) : (x5 & ~x7))));
  assign n2281 = ~n437 & ~n2282;
  assign n2282 = x0 ? (x3 | x4 | (x1 ? (x2 | ~x5) : (~x2 | x5))) : (~x1 | ~x3 | ~x4 | (~x2 ^ ~x5));
  assign n2283 = n1167 & ((~x3 & ~x5 & x7 & n542) | (n354 & (x3 ? (~x5 ^ x7) : (x5 & ~x7))));
  assign n2284 = ((x2 ? (x3 | ~x7) : (~x3 | x7)) | (x0 ? (~x1 | x4) : (x1 | ~x4))) & ((x3 ^ x7) | (x0 ? ((x2 | ~x4) & (x1 | (x2 & ~x4))) : (~x1 | x4)));
  assign z175 = ~n2287 | ~n2291 | ~n2294 | (x0 & ~n2286);
  assign n2286 = x1 ? (x3 | x4 | (x2 ? (x5 | ~x6) : (~x5 | x6))) : (~x3 | ~x4 | ~x6 | (~x2 ^ ~x5));
  assign n2287 = ~n2288 & ~n2289 & (~n1906 | ~n2076) & (n2270 | ~n2290);
  assign n2288 = x0 & ~x1 & x2 & (x3 ? (~x4 & ~x5) : (x4 & x5));
  assign n2289 = ~x2 & (x1 ? (~x4 & (~x3 ^ x5)) : (x4 & x5));
  assign n2290 = ~x0 & x6 & (~x2 ^ x5);
  assign n2291 = ~n2292 & (~x3 | n559 | n2293);
  assign n2292 = ~x2 & ((~x3 & ~x4 & x5 & ~x0 & x1) | (x0 & ~x5 & (x1 ? (x3 & ~x4) : (~x3 & x4))));
  assign n2293 = (~x0 | x1 | ~x4 | x6 | ~x7) & (x0 | x4 | (x1 ? (x6 | ~x7) : (~x6 | x7)));
  assign n2294 = (n505 | n2295) & (~n929 | n2296);
  assign n2295 = (x0 | ((~x3 | x5 | x6) & (~x2 | (x5 & (~x3 | x6))))) & (x3 | ((x6 | x7 | ~x2 | x5) & (~x0 | x2 | ~x5 | ~x6 | ~x7)));
  assign n2296 = (x0 | x1 | x4 | ~x5 | x6 | x7) & (x5 | ~x7 | ((x0 | ~x1 | x4 | ~x6) & (~x0 | ((x4 | x6) & (x1 | ~x4 | ~x6)))));
  assign z176 = n2298 | n2301 | ~n2303 | (~n559 & ~n2302);
  assign n2298 = ~x4 & ((n2299 & ~n2300) | (n292 & n335 & n992));
  assign n2299 = x0 & x6;
  assign n2300 = (~x1 | ((~x2 | x3 | ~x5) & (x5 | ~x7 | x2 | ~x3))) & (x3 | ((~x2 | ~x5 | x7) & (x1 | x2 | x5 | ~x7)));
  assign n2301 = ~n520 & ((x0 & ((~x2 & x5) | (~x1 & x2 & ~x5))) | (x5 & x7 & x1 & ~x2) | (x2 & ((~x1 & ~x5 & x7) | (~x0 & (x1 ? ~x5 : (x5 & ~x7))))));
  assign n2302 = (~x4 | ~x6 | ~x7 | x0 | x1 | ~x3) & (x6 | (x0 ? ((~x4 | x7 | x1 | ~x3) & (x4 | ~x7 | ~x1 | x3)) : (~x4 | ~x7 | (x1 ^ x3))));
  assign n2303 = n2308 & ~n2307 & ~n2306 & ~n2304 & n2305;
  assign n2304 = ~x1 & ((~x0 & ~x2 & (x3 ? (~x5 & ~x6) : (x5 & x6))) | (x3 & ~x5 & ~x6 & x0 & x2));
  assign n2305 = (x0 | ~x1 | x2 | x3 | ~x5 | ~x6) & ((x3 ? (~x5 | x6) : (x5 | ~x6)) | (x0 ? (~x1 | x2) : (x1 | ~x2)));
  assign n2306 = ~n539 & ((n321 & n615) | (n349 & n616));
  assign n2307 = n351 & n544 & ((n1906 & n374) | (n345 & n372));
  assign n2308 = (x7 | n2309) & (n2310 | ((~x1 | x2 | ~x5 | x7) & (x1 | (x2 ? (x5 | x7) : (~x5 | ~x7)))));
  assign n2309 = x0 ? (x3 | ((x1 | x2 | ~x5 | ~x6) & (~x1 | ~x2 | x5 | x6))) : (~x3 | ((~x1 | ~x2 | ~x5 | x6) & (x5 | ~x6 | x1 | x2)));
  assign n2310 = (x0 | x4 | (~x3 ^ ~x6)) & (~x0 | x3 | ~x4 | ~x6);
  assign z177 = ~n2317 | (x3 ? ~n2314 : (x1 ? ~n2313 : ~n2312));
  assign n2312 = (x2 | x4 | (x0 ? ((~x6 | x7) & (~x5 | x6 | ~x7)) : (x5 ? (x6 | x7) : (~x6 | ~x7)))) & (~x0 | ~x4 | ((x5 | x6 | ~x7) & (~x2 | (~x6 ^ x7))));
  assign n2313 = (~x4 | (x0 ? (x7 | (x2 ? (x5 | x6) : (~x5 | ~x6))) : (~x6 | ~x7 | (~x2 ^ ~x5)))) & (x0 | ~x2 | x4 | x5 | (~x6 ^ x7));
  assign n2314 = x1 ? (x2 | n2316) : n2315;
  assign n2315 = (~x4 | (x0 ? ((x6 | x7 | x2 | ~x5) & (~x6 | ~x7 | ~x2 | x5)) : (~x2 | ((x6 | ~x7) & (x5 | ~x6 | x7))))) & (x0 | x4 | ((~x5 | ~x6 | x7) & (x2 | (~x6 ^ x7))));
  assign n2316 = (x4 | ((x6 | x7 | x0 | x5) & (~x0 | ((x6 | ~x7) & (x5 | ~x6 | x7))))) & (x0 | ~x4 | ~x5 | (~x6 ^ x7));
  assign n2317 = ~n2319 & n2320 & ~n2321 & (n425 | n2318) & ~n2322;
  assign n2318 = x1 ? ((x0 | ~x2 | ~x3 | x4) & (x3 | ((~x0 | x4 | (~x2 & x5)) & (~x4 | ~x5 | x0 | x2)))) : ((~x0 | ~x2 | ~x3 | ~x4 | ~x5) & ((~x4 ^ x5) | (x0 ? (x2 | ~x3) : (~x2 | x3))));
  assign n2319 = ~x0 & (x1 ? (~n950 & ~n539) : (n1190 & n929));
  assign n2320 = (~x0 | x1 | x2 | x3 | ~x4 | ~x6) & ((x3 ^ x6) | ((x0 | x1 | x2 | ~x4) & (~x0 | (x1 ? (x2 | ~x4) : (~x2 | x4)))));
  assign n2321 = ~x0 & ((x3 & ~x4 & ~x6 & ~x1 & x2) | (x1 & ((~x4 & x6 & ~x2 & ~x3) | (x4 & ~x6 & x2 & x3))));
  assign n2322 = ~n520 & ((~x0 & ~x1 & x2 & x4 & x5) | (x0 & ~x2 & ~x4 & (x1 ^ ~x5)));
  assign z178 = ~n2328 | (x0 ? ~n2326 : (n2325 | (~x4 & ~n2324)));
  assign n2324 = (x7 | ((x6 | ((~x1 | (x2 ? (x3 | ~x5) : (~x3 | x5))) & (x1 | x2 | x3 | ~x5))) & (x1 | ~x6 | (x2 ? (~x3 | ~x5) : (x3 | x5))))) & (x1 | ~x5 | ~x7 | (x2 ? (~x3 | x6) : (x3 | ~x6)));
  assign n2325 = x5 & n1230 & (x1 ? (~x3 & ~n437) : (x3 & n374));
  assign n2326 = x1 ? (~n929 | ~n339) : n2327;
  assign n2327 = (x2 | ~x3 | ~x4 | ~x5 | ~x6 | ~x7) & (x5 | (((~x4 ^ ~x7) | (x2 ? (~x3 | x6) : (x3 | ~x6))) & (~x2 | ~x3 | ~x4 | ~x6 | x7)));
  assign n2328 = n2330 & (n1054 | n2329) & (x1 ? n2332 : n2331);
  assign n2329 = (x4 | x6 | ~x7 | x1 | ~x2 | x3) & (x2 | ((~x4 | x6 | x7 | x1 | ~x3) & (~x1 | ~x6 | (x3 ? (x4 | ~x7) : (~x4 | x7)))));
  assign n2330 = x2 ? ((x7 | (x1 ^ ~x4) | (x0 ^ ~x3)) & (~x3 | ~x7 | (x0 ? (x1 | x4) : (~x1 | ~x4)))) : ((~x1 | ((x4 | ~x7 | x0 | x3) & (~x0 | ~x3 | (x4 ^ x7)))) & (x0 | x1 | ((~x4 | ~x7) & (~x3 | x4 | x7))));
  assign n2331 = x0 ? (x2 ? ((x5 | ~x7 | x3 | x4) & (~x5 | x7 | ~x3 | ~x4)) : (x4 ? ((x5 | x7) & (x3 | ~x5 | ~x7)) : ((~x5 | x7) & (~x3 | x5 | ~x7)))) : (~x2 | ((x5 | ~x7 | ~x3 | x4) & (x3 | (x4 ? (x5 ^ x7) : (~x5 | x7)))));
  assign n2332 = x7 ? ((~x4 ^ x5) | (x0 ? (x2 | x3) : (x2 ^ ~x3))) : ((~x0 | x2 | x3 | x4 | x5) & (x0 | ((x2 | ~x4 | ~x5) & (x4 | x5 | ~x2 | x3))));
  assign z179 = ~n2343 | ~n2342 | n2341 | n2340 | n2334 | n2337;
  assign n2334 = x0 & (x2 ? ~n2336 : ~n2335);
  assign n2335 = (~x7 | (x1 ? (~x5 | (x3 ? (x4 | ~x6) : (~x4 | x6))) : (x3 | x5 | (x4 ^ x6)))) & (~x3 | ~x4 | x5 | x7 | (~x1 ^ ~x6));
  assign n2336 = (~x5 | x6 | x7 | ~x1 | x3 | x4) & (x1 | ((~x3 | ~x4 | ~x5 | ~x6 | x7) & (x4 | (x3 ? (x6 | (~x5 ^ x7)) : (~x6 | (x5 ^ x7))))));
  assign n2337 = ~x0 & (x5 ? ~n2339 : ~n2338);
  assign n2338 = x1 ? ((x2 | x3 | ~x4 | x6 | ~x7) & (~x2 | ~x3 | x4 | ~x6 | x7)) : ((x2 | ~x4 | (x3 ? (x6 | ~x7) : (~x6 | x7))) & (x4 | ((x6 | ~x7 | x2 | x3) & (~x2 | (x3 ? (x6 | x7) : (~x6 | ~x7))))));
  assign n2339 = x2 ? (x1 ? (x6 | (x3 ? (~x4 | x7) : (x4 | ~x7))) : (~x6 | (x3 ? (~x4 | ~x7) : (x4 | x7)))) : (x7 | ((~x1 | (x3 ? (x4 | ~x6) : (~x4 | x6))) & (x4 | x6 | x1 | ~x3)));
  assign n2340 = x1 & ((~x0 & x2 & ~x3 & x5 & x6) | (~x2 & ((~x5 & x6 & ~x0 & ~x3) | (x0 & (x3 ? (~x5 & ~x6) : (x5 & x6))))));
  assign n2341 = x5 & n1100 & ((x1 & ~x2 & x4 & x6) | (~x1 & (x2 ? (~x4 & x6) : (x4 & ~x6))));
  assign n2342 = ((~x2 ^ x5) | ((~x3 | x6 | x0 | ~x1) & (~x0 | x1 | (x3 ^ x6)))) & (x0 | x1 | ((x5 | ~x6 | x2 | ~x3) & (~x5 | x6 | ~x2 | x3)));
  assign n2343 = (x3 | n2345) & (n2344 | (~x2 ^ ~x4));
  assign n2344 = (x0 | ~x1 | x5 | (x3 ^ x6)) & (x1 | (x0 ? (x3 ? (~x5 | x6) : (x5 | ~x6)) : (x3 ? (x5 | x6) : (~x5 | ~x6))));
  assign n2345 = (x0 | x1 | x2 | ~x4 | x5 | x6) & (~x0 | ((x1 | x2 | ~x4 | ~x5 | ~x6) & (~x1 | x4 | (x2 ? x5 : (~x5 | x6)))));
  assign z180 = ~n2354 | n2347 | ~n2349;
  assign n2347 = x1 & ((~x2 & ~n2348) | (~x0 & n929 & n1197));
  assign n2348 = (x0 | ~x4 | ((~x6 | ~x7 | x3 | ~x5) & (x6 | x7 | ~x3 | x5))) & (~x3 | x4 | ~x5 | ~x6 | ~x7) & (x3 | x5 | x6 | x7 | (~x0 & x4));
  assign n2349 = ~n2352 & n2353 & (n425 | n2350) & (~x2 | n2351);
  assign n2350 = (x5 | ((~x0 | ~x1 | x2 | ~x3 | ~x4) & (x0 | ((~x1 | ~x2 | ~x3 | x4) & (x1 | x2 | x3 | ~x4))))) & (x1 | ~x2 | ~x5 | (x3 ^ x4));
  assign n2351 = (x6 | (x0 ? (x3 | (x1 ? (x4 | x5) : (~x4 | ~x5))) : (~x1 | ~x3 | (~x4 ^ x5)))) & (x0 | ~x6 | ((~x1 | x3 | ~x4) & (x4 | ~x5 | x1 | ~x3)));
  assign n2352 = ~x1 & ((x4 & ((x2 & ~x5 & (x3 ^ ~x6)) | (x5 & x6 & ~x2 & x3))) | (~x2 & ~x4 & (x3 ? (~x5 & ~x6) : (x5 & x6))));
  assign n2353 = (~n542 | ((x3 | x4 | ~x5 | x6) & (~x3 | (x4 ? (~x5 | x6) : (x5 | ~x6))))) & (x3 | x4 | x5 | ~x6 | ~n317);
  assign n2354 = (n437 | n2355) & (x1 | (x0 ? n2356 : n2357));
  assign n2355 = x1 ? (x2 ? ((x3 | x4 | ~x5) & (x0 | (x3 ? (~x4 | ~x5) : x4))) : (x3 | ~x4)) : (x4 ? ((x2 | ~x3 | x5) & (x3 | ~x5 | x0 | ~x2)) : ((~x0 | ((~x3 | ~x5) & (x2 | x3 | x5))) & (~x3 | (~x2 ^ x5))));
  assign n2356 = (x4 | ((~x6 | ~x7 | x3 | x5) & (~x3 | ~x5 | (x2 ? (~x6 | ~x7) : (x6 | x7))))) & (x2 | x3 | ((x5 | ~x6 | ~x7) & (~x4 | ~x5 | x6 | x7)));
  assign n2357 = (x5 | ~x6 | ~x7 | x2 | ~x3 | ~x4) & (x3 | ((~x4 | ~x5 | x6 | x7) & (~x2 | x4 | x5 | ~x6 | ~x7)));
  assign z181 = n2359 | n2361 | ~n2365 | (~n617 & ~n2364);
  assign n2359 = x2 & ((n1585 & n1197) | (~x1 & ~n2360));
  assign n2360 = (x3 | x4 | x5 | x6 | x7) & (~x5 | ((x0 | x7 | (x3 ? (x4 | ~x6) : (~x4 | x6))) & (~x0 | ~x3 | x4 | x6 | ~x7)));
  assign n2361 = ~x2 & (x7 ? ~n2363 : ~n2362);
  assign n2362 = (x3 | ((~x6 | ((x1 | x4 | x5) & (x0 | (x4 ^ x5)))) & (~x0 | ~x1 | ~x4 | x5 | x6))) & (~x0 | ~x1 | ~x3 | ~x5 | (x4 ^ x6));
  assign n2363 = (x0 | ((x1 | x3 | x4 | ~x5 | ~x6) & (~x1 | ~x3 | ~x4 | x5 | x6))) & (x4 | ~x5 | ~x6 | ~x0 | ~x3);
  assign n2364 = x4 ? ((~x7 | ((x1 | x3 | ~x5) & (x0 | ((x3 | ~x5) & (x1 | ~x3 | x5))))) & (~x0 | x1 | x3 | x5 | x7)) : ((~x0 | ((x3 | x5 | ~x7) & (~x5 | x7 | x1 | ~x3))) & (~x1 | ((x3 | x5 | ~x7) & (~x5 | x7 | x0 | ~x3))));
  assign n2365 = ~n2367 & ~n2368 & n2370 & (~x2 | n2366);
  assign n2366 = (x4 | x5 | ~x7 | ~x0 | x1 | ~x3) & (x3 | ((x0 | ~x1 | ~x4 | ~x5 | x7) & (x1 | ((x5 | ~x7 | x0 | x4) & (~x0 | ~x5 | (~x4 ^ x7))))));
  assign n2367 = ~x0 & (x3 ? ((x5 & ~x7 & ~x2 & x4) | (~x5 & x7 & x2 & ~x4)) : (x2 ? (x4 ? (~x5 & ~x7) : (x5 & x7)) : (x4 ? (~x5 & x7) : (x5 & ~x7))));
  assign n2368 = ~n440 & ((x2 & n2369) | (~x0 & (x2 ? n361 : n373)));
  assign n2369 = x0 & (x1 ? (~x3 & ~x4) : (x3 & x4));
  assign n2370 = ~n532 | ((x7 | (x3 ? ((x4 | x5) & (x1 | ~x4 | ~x5)) : (x4 | ~x5))) & (~x4 | ~x7 | (x5 & (~x1 | x3))));
  assign z182 = ~n2374 | (x1 & (x5 ? ~n2373 : ~n2372));
  assign n2372 = (x2 | ((x0 | x3 | ~x4 | ~x6 | ~x7) & (~x3 | ((~x6 | x7 | x0 | ~x4) & (~x0 | ~x7 | (~x4 ^ x6)))))) & (~x0 | x3 | x7 | (~x4 ^ x6));
  assign n2373 = (~x4 | x6 | x7 | ~x0 | x2 | ~x3) & (x0 | (x3 ? (x4 ? (~x6 | ~x7) : (x6 | x7)) : ((x4 | x6 | ~x7) & (~x6 | x7 | ~x2 | ~x4))));
  assign n2374 = ~n2377 & n2378 & (x1 | (x3 & n2375) | (~x3 & n2376));
  assign n2375 = x4 ? ((~x6 | x7 | x0 | x5) & (~x0 | ~x7 | ((x5 | x6) & (x2 | ~x5 | ~x6)))) : ((~x0 | ~x2 | x5 | ~x6 | ~x7) & (x0 | x6 | ((x5 | ~x7) & (~x2 | ~x5 | x7))));
  assign n2376 = x0 ? ((x2 | x4 | ~x5 | x6 | ~x7) & (~x4 | x7 | (x5 ^ x6))) : ((~x6 | ~x7 | ~x4 | x5) & (x4 | ((~x6 | x7 | x2 | ~x5) & (~x2 | x6 | (x5 ^ x7)))));
  assign n2377 = n310 & ((~x1 & ~x2 & ~x3 & ~x4 & x5) | (x1 & x4 & ((x3 & ~x5) | (x2 & ~x3 & x5))));
  assign n2378 = ~n2380 & (~x6 | n2381) & (n2379 | (x1 & x2));
  assign n2379 = (~x5 | x6 | x3 | ~x4) & (~x3 | ((x5 | ~x6 | x0 | x4) & (~x0 | (x4 ? (x5 | ~x6) : (~x5 | x6)))));
  assign n2380 = (~x5 ^ x6) & ((~x0 & ~x1 & x3 & x4) | (~x3 & ~x4 & (x0 | x1)));
  assign n2381 = x0 ? (x2 | ((x4 | x5 | x1 | ~x3) & (~x4 | ~x5 | ~x1 | x3))) : (~x2 | ((x4 | ~x5 | x1 | x3) & (~x1 | ~x3 | x5)));
  assign z183 = ~n2389 | (x1 ? ~n2385 : (x3 ? ~n2383 : ~n2384));
  assign n2383 = x5 ? ((~x0 | x4 | (x6 ^ x7)) & (~x2 | ((x0 | (x4 ? (x6 | ~x7) : (~x6 | x7))) & (~x6 | x7 | ~x0 | ~x4)))) : ((~x6 | x7 | x0 | ~x4) & (x2 | ((x0 | x4 | x6 | x7) & (~x0 | ~x4 | (x6 ^ x7)))));
  assign n2384 = x5 ? ((x0 | ~x2 | x4 | ~x6 | x7) & (~x0 | ((x4 | x6 | x7) & (~x2 | ~x6 | (~x4 ^ x7))))) : (((~x0 ^ x6) | ((~x4 | x7) & (x2 | x4 | ~x7))) & (~x6 | ~x7 | ~x0 | ~x4));
  assign n2385 = ~n2386 & (n585 | n2388) & (n1015 | n2387);
  assign n2386 = x6 & n544 & ((x2 & x4 & ~x5 & x7) | (~x2 & ~x7 & (~x4 ^ ~x5)));
  assign n2387 = (~x0 | x2 | ~x3 | ~x6 | x7) & (x0 | x6 | ~x7 | (x2 & x3));
  assign n2388 = (~x0 | x2 | x3 | ~x5 | x7) & (x0 | ~x2 | ~x3 | x5 | ~x7);
  assign n2389 = ~n2391 & ~n2392 & ~n2393 & (n589 | n2390) & ~n2395;
  assign n2390 = (~x5 | ((x0 | ((x1 | x2 | x7) & (~x1 | ~x2 | ~x3 | ~x7))) & (~x0 | x1 | x2 | x3 | ~x7))) & (~x0 | x5 | x7 | (x1 ? x3 : (~x2 | ~x3)));
  assign n2391 = ~x1 & (x0 ? ((x6 & ~x7 & ~x2 & x4) | (~x6 & x7 & x2 & ~x4)) : ((~x6 & x7 & ~x2 & x4) | (x2 & ~x4 & (~x6 ^ x7))));
  assign n2392 = x1 & ((~x2 & x7 & (x0 ? (~x4 ^ x6) : (~x4 & x6))) | (~x0 & ~x7 & ((~x4 & ~x6) | (x2 & x4 & x6))));
  assign n2393 = ~n368 & ((x3 & n345 & n370) | (x1 & ~n2394));
  assign n2394 = (~x2 | x3 | x4 | ~x7) & (x2 | ~x3 | ~x4 | x7);
  assign n2395 = x4 & x7 & n354 & (x0 ? (x3 & x6) : (~x3 & ~x6));
  assign z184 = ~n2399 | (x5 ? (x7 ? ~n2398 : ~n2397) : (x7 ? ~n2397 : ~n2398));
  assign n2397 = (~x6 | (x0 ? (x1 | (x2 & (x3 | x4))) : (~x1 | ~x2 | (~x3 & ~x4)))) & (x0 | x6 | ((~x3 | ~x4 | x1 | ~x2) & (~x1 | (x2 & x3 & x4))));
  assign n2398 = (x1 | ((x2 | ((~x3 | x6) & (x0 | ~x4))) & (~x6 | ((x0 | (~x2 & ~x3)) & (~x2 | ~x3 | ~x4))) & (~x2 | x6 | (~x0 & (x3 | x4))))) & (x3 | ~x6 | ~x1 | x2) & (~x0 | ((x4 | x6 | x2 | ~x3) & (~x1 | ((x3 | x4 | ~x6) & (x2 | (x3 & ~x6))))));
  assign n2399 = ~n2401 & (~n544 | n2404) & (x0 ? n2400 : n2403);
  assign n2400 = (x6 | ((x1 | x2 | x3 | x5) & (~x1 | ~x5 | (x2 ? (x3 | x4) : (~x3 | ~x4))))) & (x1 | ~x2 | x5 | ~x6 | (~x3 ^ x4));
  assign n2401 = x3 & ((x0 & ~n2402) | (n292 & n351 & n992));
  assign n2402 = (~x5 | x6 | x7 | ~x1 | x2 | x4) & (x5 | ~x6 | ~x7 | x1 | ~x2 | ~x4);
  assign n2403 = (~x1 | x2 | ~x3 | ~x5 | ~x6) & (x1 | ((~x2 | ~x5 | x6 | (~x3 ^ x4)) & (x4 | x5 | ~x6 | x2 | x3)));
  assign n2404 = (x5 | ~x6 | ~x7 | x1 | x2 | ~x4) & (x4 | ~x5 | ((~x1 | ~x2 | ~x6 | x7) & (x1 | x6 | (x2 ^ ~x7))));
  assign z185 = ~n2406 | (~n437 & ~n2411) | (~n425 & ~n2410);
  assign n2406 = ~n2408 & ~n2409 & (~n958 | ~n339) & (~x6 | n2407);
  assign n2407 = (~x3 | ((~x2 | ~x4 | x5 | x0 | ~x1) & (~x0 | ((~x4 | ~x5 | x1 | ~x2) & (x4 | x5 | ~x1 | x2))))) & (x0 | x3 | ((x1 | (x2 ? (x4 | x5) : (~x4 | ~x5))) & (~x1 | ~x2 | x4 | ~x5)));
  assign n2408 = ~x0 & ((x3 & ((x1 & x2 & ~x4 & x6) | (~x1 & (x2 ? (x4 & ~x6) : x6)))) | (x1 & ~x3 & (x2 ? (x4 & x6) : ~x6)));
  assign n2409 = x0 & ((~x3 & x6 & x1 & ~x2) | (~x1 & ~x6 & (x2 ? (~x3 & ~x4) : x3)));
  assign n2410 = x0 ? (x1 ? (x2 ? (x3 | x4) : (~x3 | (~x4 & ~x5))) : (x2 | x3)) : (~x2 | ((~x3 | (x1 ? (~x4 | ~x5) : x4)) & (x1 | (x4 ? x3 : ~x5))));
  assign n2411 = x0 ? (x1 | ~x2 | (x4 ? (x3 & x5) : ~x3)) : (x1 ? ((x2 | ~x3) & (x4 | x5 | ~x2 | x3)) : (x2 | x3 | (x4 & x5)));
  assign z186 = ~n2415 | ~n2418 | (~x6 & (n2413 | (x2 & ~n2414)));
  assign n2413 = ~n1355 & ((~x0 & x4 & (x2 ? (x3 & ~x5) : (~x3 & x5))) | (x0 & ~x2 & x3 & ~x4 & ~x5));
  assign n2414 = (~x4 | ~x5 | x7 | ~x0 | x1 | ~x3) & (x3 | (x0 ? ((~x5 | ~x7 | x1 | x4) & (x5 | x7 | ~x1 | ~x4)) : (x4 | (x1 ? (~x5 | x7) : (x5 | ~x7)))));
  assign n2415 = ~n2417 & (~n1415 | ~n1018) & (~x4 | ~n349 | n2416);
  assign n2416 = (~x2 | ~x3 | ~x5 | x7) & (x2 | x3 | x5 | ~x7);
  assign n2417 = x2 & (((x3 ^ x4) & ((~x1 & ~x7) | (~x0 & x1 & x7))) | (~x0 & ~x1 & x3 & x4 & x7) | (x0 & x1 & ~x3 & ~x4 & ~x7));
  assign n2418 = ~n2421 & (n440 | n2419) & (x4 | n2420);
  assign n2419 = (x0 | x3 | (x1 ? (~x2 | x4) : (x2 | ~x4))) & (~x0 | x1 | ~x2 | ~x3 | ~x4);
  assign n2420 = (x0 | x1 | x3 | ~x5 | x7) & (~x0 | ((x3 | x5 | ~x7 | x1 | ~x2) & (~x3 | ~x5 | x7 | ~x1 | x2)));
  assign n2421 = ~x2 & (x3 ? (x1 ? (~x7 & (~x0 | x4)) : x7) : ((x1 & ~x4 & x7) | (x0 & (~x1 ^ x7))));
  assign z187 = n2423 | n2427 | ~n2428 | (~x3 & ~n2426);
  assign n2423 = x7 & (x1 ? ~n2425 : ~n2424);
  assign n2424 = x2 ? ((x3 ? (~x4 | x6) : (x4 | ~x6)) | (~x0 ^ ~x5)) : (x6 | ((x4 | x5 | ~x0 | ~x3) & (x0 | x3 | (x4 ^ x5))));
  assign n2425 = (x4 | x5 | ~x6 | ~x0 | x2 | ~x3) & (x0 | ((x2 | x3 | ~x4 | ~x5 | ~x6) & (~x2 | ((x5 | ~x6 | ~x3 | ~x4) & (~x5 | x6 | x3 | x4)))));
  assign n2426 = (~x0 | x1 | ~x2 | ~x4) & (x0 | (x1 ? ((~x5 | ~x6 | ~x2 | ~x4) & (x5 | x6 | x2 | x4)) : (~x5 | (x2 ? (x4 | x6) : (~x4 | ~x6)))));
  assign n2427 = ~n1054 & ((n542 & ~n447) | (x3 & n354 & n547));
  assign n2428 = n2430 & ~n2429 & (x5 | ~n321 | ~n373 | n1042);
  assign n2429 = ~x3 & x5 & ((x0 & ~x2 & ~x4 & ~x6) | (~x0 & x2 & (x4 ^ x6)));
  assign n2430 = (x0 | ~x2 | ~x4 | (x3 ^ x5)) & (x2 | ((~x3 | x4 | (x0 & ~x5)) & (~x0 | x5 | (x3 ^ x4))));
  assign z188 = n2432 | ~n2433 | n2442 | (x1 & ~n2441);
  assign n2432 = ~x2 & ((~x0 & x1 & x3 & x4 & x5) | (~x1 & ((~x4 & x5 & ~x0 & ~x3) | (x4 & (x0 ? (~x3 ^ x5) : (x3 & ~x5))))));
  assign n2433 = ~n2434 & ~n2435 & n2436 & n2440 & (x1 | n2439);
  assign n2434 = ~n1015 & ((x0 & ~n1232) | (~x2 & n783 & ~n798));
  assign n2435 = ~n390 & ((x0 & ~n402) | (x2 & n783 & n784));
  assign n2436 = x1 ? (~x6 | n2437) : ((x6 | n2437) & (~x0 | ~x3 | n2438));
  assign n2437 = (~x0 | x2 | x3 | x4 | x5 | x7) & (x0 | ~x4 | ~x7 | (x2 ? (~x3 | x5) : (x3 | ~x5)));
  assign n2438 = (x2 | x4 | (x5 ? (~x6 | x7) : (x6 | ~x7))) & (~x2 | ~x4 | ~x5 | x6 | ~x7);
  assign n2439 = ((x0 ? (x2 | x4) : (~x2 | ~x4)) | (x3 ? (~x5 ^ x6) : (~x5 | ~x6))) & (x4 | x5 | x6 | ~x0 | ~x2 | x3);
  assign n2440 = ((x1 ^ ~x2) | ((~x0 | (x3 ? (x4 | ~x5) : (~x4 | x5))) & (x4 | ~x5 | x0 | x3))) & (~x0 | ~x1 | ~x2 | x3 | x4 | x5) & (x0 | ~x3 | ((~x2 | x4 | x5) & (~x1 | ((x4 | x5) & (~x2 | ~x4 | ~x5)))));
  assign n2441 = (~x0 | x2 | ~x3 | ~x4 | ~x5 | ~x6) & (x0 | ((~x2 | x4 | ~x5 | (~x3 ^ x6)) & (~x4 | x5 | ((x3 | x6) & (x2 | ~x3 | ~x6)))));
  assign n2442 = ~x0 & ((n1252 & n786) | (~x7 & ~n2443));
  assign n2443 = x1 ? ((x4 | ~x5 | x6 | x2 | ~x3) & (~x4 | x5 | ~x6 | ~x2 | x3)) : (~x3 | ~x6 | (x2 ? (~x4 | ~x5) : (x4 | x5)));
  assign z189 = ~n2449 | ~n2452 | (~x2 & (~n2445 | ~n2448));
  assign n2445 = (~x5 | n2446) & (~x0 | x5 | n2447);
  assign n2446 = (~x4 | ~x6 | x7 | ~x0 | x1 | ~x3) & (x0 | (x1 ? (~x6 | (x3 ? (x4 | x7) : (~x4 | ~x7))) : (x6 | ((x4 | x7) & (x3 | ~x4 | ~x7)))));
  assign n2447 = (x1 | x3 | x4 | x6 | ~x7) & (~x1 | ~x3 | (x4 ? (x6 | ~x7) : (x6 ^ x7)));
  assign n2448 = (x5 | ((~x0 | ((x1 | x4 | ~x6) & (~x4 | x6 | ~x1 | x3))) & (x4 | ((x1 | x3 | ~x6) & (x0 | ~x1 | ~x3 | x6))) & (~x4 | (x1 ^ x6) | (x0 & ~x3)))) & (x4 | ((~x5 | x6 | ~x1 | x3) & (~x0 | (x1 ? (~x5 | x6) : (x3 | ~x6))))) & (~x4 | ~x5 | (x0 ? (x1 ^ x6) : (x1 | ~x6)));
  assign n2449 = (~x2 | n2450) & (n416 | n2451);
  assign n2450 = x5 ? ((~x0 | ((x4 | x6 | ~x1 | x3) & (x1 | ~x4 | ~x6))) & (x1 | x3 | ~x4 | ~x6) & (x0 | (x1 ? (~x4 ^ x6) : (x4 | x6)))) : ((x1 | ((~x0 | (~x4 ^ x6)) & (~x4 | ~x6 | x0 | ~x3))) & (x0 | ~x1 | x4 | x6));
  assign n2451 = x0 ? ((~x1 | ~x2 | x3 | x4 | x7) & (x1 | x2 | (x3 ? (x4 | ~x7) : (~x4 | x7)))) : ((x1 | ~x2 | ~x3 | ~x4 | ~x7) & (~x1 | x2 | x3 | x4 | x7));
  assign n2452 = (n699 | n2453) & (~x2 | (~n2454 & ~n2456 & n2457));
  assign n2453 = (x3 | x5 | ~x6 | x0 | x1 | ~x2) & (x2 | ((x0 | ~x3 | (x1 ? (~x5 | x6) : (x5 | ~x6))) & (x3 | x5 | ~x6 | ~x0 | ~x1)));
  assign n2454 = ~n2455 & ~x1 & ~x6;
  assign n2455 = (~x5 | ~x7 | ~x0 | ~x4) & (x0 | x5 | (x3 ? (x4 | x7) : (~x4 | ~x7)));
  assign n2456 = ~n425 & (x3 ? (n351 & n349) : (n850 & n321));
  assign n2457 = (~x0 | x1 | ~x3 | x7 | n420) & (x0 | ~x1 | (x3 ? ~n1018 : (~x7 | n420)));
  assign z190 = ~n1613 | (x2 ? ~n2459 : (x5 ? ~n1611 : ~n1612));
  assign n2459 = (~x6 | n1609) & (x0 | x6 | n2460);
  assign n2460 = (x1 | x3 | x5 | ~x7) & (~x3 | ((x4 | x5 | ~x7) & (~x1 | ((x5 | ~x7) & (~x4 | ~x5 | x7)))));
  assign z191 = ~n2463 | ~n1618 | (~x3 & ~x7 & ~n2462);
  assign n2462 = (~x4 | (x0 ? (x5 | (x1 ? x6 : (~x2 | ~x6))) : (~x5 | (x1 ? (x2 | x6) : (~x2 | ~x6))))) & (x1 | x4 | (~x2 ^ x6) | (~x0 ^ x5));
  assign n2463 = (~x6 | (x7 ? n2464 : n2465)) & (~n647 | ~n1631) & (x6 | (x7 ? n2465 : n2464));
  assign n2464 = (x2 | ((x3 | ~x4 | x5 | x0 | ~x1) & ((~x0 & ~x5) | (x1 ? (x3 | x4) : (~x3 | ~x4))))) & (x0 | ~x2 | ((x4 | x5 | x1 | x3) & (~x1 | (x3 ? x4 : (~x4 | ~x5)))));
  assign n2465 = x1 ? ((x0 | ~x2 | x3 | x4 | x5) & (x2 | ~x3 | (~x4 & (~x0 | ~x5)))) : ((x3 | ((~x0 | ~x5 | (x2 ^ x4)) & (x2 | ~x4 | (x0 & x5)))) & (~x2 | ~x3 | x4 | (x0 & x5)));
  assign z192 = ~n2471 | (x3 ? (n2468 | (n1883 & ~n2467)) : ~n2469);
  assign n2467 = (x1 | ~x2 | x4 | (x6 ^ x7)) & (x2 | ((~x1 | ~x6 | (x4 ^ x7)) & (x6 | ~x7 | x1 | x4)));
  assign n2468 = ~x5 & n1050 & ((x1 & ~x2 & x6 & ~x7) | (~x1 & (x2 ? (~x6 ^ x7) : (~x6 & x7))));
  assign n2469 = x5 ? ((x0 | n1638) & (~x4 | x7 | ~n2470)) : ((~x0 | n1638) & (x4 | ~x7 | ~n2470));
  assign n2470 = x6 & x2 & ~x0 & x1;
  assign n2471 = ~n1642 & ~n2473 & ~n2474 & n2475 & (x7 | n2472);
  assign n2472 = (~x3 | x4 | x5 | ~x0 | x1 | ~x2) & (x3 | ((~x0 | x1 | ~x2 | ~x4 | ~x5) & (x2 | (~x4 ^ x5) | (x0 ^ ~x1))));
  assign n2473 = ~x0 & ((~x1 & ~x2 & ~x3 & x4 & ~x7) | (x3 & (x2 ? ((~x4 & ~x7) | (x1 & x4 & x7)) : (~x4 & x7))));
  assign n2474 = x0 & (x2 ? (x7 & ((~x3 & ~x4) | (~x1 & x3 & x4))) : (~x7 & ((x3 & x4) | (x1 & ~x3 & ~x4))));
  assign n2475 = x0 | ((x7 | n948) & (~x5 | ~x7 | ~n354 | ~n361));
  assign z193 = n2477 | ~n2478 | ~n2481 | n2485 | (~x0 & ~n2484);
  assign n2477 = x1 & ((~x3 & x4 & ~x5 & ~x0 & x2) | (~x4 & (x0 ? (x2 ? (~x3 & x5) : (x3 & ~x5)) : ((x3 & x5) | (~x2 & ~x3 & ~x5)))));
  assign n2478 = ~n2479 & (n585 | n2480);
  assign n2479 = ~x1 & ((~x0 & x2 & ~x3 & ~x4 & ~x5) | (x4 & ((~x3 & x5 & ~x0 & ~x2) | (x0 & ((x3 & x5) | (~x2 & ~x3 & ~x5))))));
  assign n2480 = (x2 | ((~x0 | ~x1 | ~x3 | ~x5 | x7) & (x0 | x1 | x3 | x5 | ~x7))) & (x1 | ~x2 | (x3 ^ x7) | (~x0 ^ x5));
  assign n2481 = (~x0 | n2482) & (~n345 | n2483);
  assign n2482 = x3 ? ((~x5 ^ x6) | (x1 ? (x2 | ~x4) : x4)) : (((x1 ^ ~x2) | (x4 ? (x5 | x6) : (~x5 | ~x6))) & (x1 | x2 | x4 | x5 | x6));
  assign n2483 = (x5 | ~x6 | x7 | x0 | ~x3 | ~x4) & (x4 | ~x5 | ((x6 | ~x7 | x0 | ~x3) & (~x0 | ~x6 | (x3 ^ ~x7))));
  assign n2484 = x3 ? ((~x5 | ~x6 | ~x1 | ~x4) & (x1 | (x4 ? (x5 | x6) : (~x5 | ~x6)))) : ((~x1 | ~x2 | x4 | x5 | x6) & ((~x5 ^ x6) | (x1 ? (x2 | ~x4) : (~x2 ^ ~x4))));
  assign n2485 = x1 & ((~x6 & ~n2486) | (x6 & n1354 & n487 & ~n392));
  assign n2486 = (x3 | (x0 ? ((~x5 | ~x7 | x2 | x4) & (x5 | x7 | ~x2 | ~x4)) : (~x4 | (x2 ? (~x5 | x7) : (x5 | ~x7))))) & (x0 | ~x3 | ~x4 | (x2 ? (~x5 | ~x7) : (x5 | x7)));
  assign z194 = ~n2494 | (x5 ? ~n2490 : (x1 ? ~n2489 : ~n2488));
  assign n2488 = x0 ? ((x2 | x7 | ((~x4 | ~x6) & (x3 | x4 | x6))) & (x6 | ~x7 | ~x3 | ~x4) & (~x2 | ((~x4 | x6 | ~x7) & (~x3 | (x4 ? x6 : (~x6 | ~x7)))))) : ((((x4 | ~x6) & (x3 | ~x4 | x6)) | (x2 ^ ~x7)) & (~x4 | x6 | x7 | x2 | ~x3) & (~x6 | ~x7 | x3 | x4));
  assign n2489 = ((x2 ^ ~x7) | ((x4 | ~x6 | ~x0 | x3) & (x0 | ((x4 | x6) & (~x3 | ~x4 | ~x6))))) & (x3 | ((~x4 | ((~x6 | ~x7 | x0 | ~x2) & (~x0 | x6 | x7))) & (x0 | x4 | ((x6 | ~x7) & (x2 | ~x6 | x7))))) & (~x0 | x2 | x7 | ((~x4 | x6) & (~x3 | x4 | ~x6)));
  assign n2490 = ~n2492 & ~n2493 & (x2 ? (~n349 | n390) : n2491);
  assign n2491 = (~x0 | x1 | x4 | ~x6 | x7) & (x0 | x6 | (x1 ? (~x4 | ~x7) : (x4 | x7)));
  assign n2492 = ~n585 & (x0 ? (x1 ? (~x2 & ~x7) : (x2 & x7)) : (~x1 & (x2 ? ~x7 : (~x3 & x7))));
  assign n2493 = ~x2 & x4 & n374 & (x0 ? n1671 : n647);
  assign n2494 = (x0 | n2498) & (~x0 | n2495) & (n2496 | n2497);
  assign n2495 = (~x7 | ((x1 | x2 | x4 | x6) & (~x1 | ((x4 | ~x6 | ~x2 | x3) & (x2 | ~x4 | x6))))) & (x1 | x7 | ((~x3 | x4 | x6) & (~x2 | (x4 ^ x6))));
  assign n2496 = (~x0 | x2 | ~x6 | ~x7) & (x0 | (x2 ? (x6 | ~x7) : (~x6 | x7)));
  assign n2497 = x1 ? (~x3 | x4) : ~x4;
  assign n2498 = ((x4 ? (x6 | x7) : (~x6 | ~x7)) | (x1 ? x2 : (~x2 | ~x3))) & (~x4 | x6 | ~x7 | x1 | x2 | ~x3) & (~x1 | ~x2 | ~x6 | ((~x3 | ~x4 | ~x7) & (x4 | x7)));
  assign z195 = n2500 | ~n2504 | (~x0 & ~n2503) | (~n665 & ~n2502);
  assign n2500 = ~x7 & ((~x5 & ~n2501) | (n451 & n313 & n992));
  assign n2501 = x6 ? ((~x3 | (x0 ? (x1 | ~x2) : (x2 | ~x4))) & (~x0 | ((x1 | ~x2 | ~x4) & (x3 | x4 | ~x1 | x2))) & (x0 | (x1 ? (~x2 | (x3 & x4)) : x2))) : (x0 ? (~x2 | (x4 ? x3 : x1)) : (x2 | (~x1 & (x3 | ~x4))));
  assign n2502 = x0 ? ((~x1 | ((x2 | x6) & (x4 | ~x6 | ~x2 | x3))) & (x2 | ((x3 | x4 | x6) & (~x6 | (x1 & (~x3 | ~x4)))))) : ((~x1 | ((~x2 | ~x3 | x6) & (x4 | ~x6 | x2 | x3))) & (~x2 | ~x3 | x4 | x6) & (x1 | ((~x3 | (x2 ? ~x6 : (~x4 | x6))) & (~x2 | (x6 ? ~x4 : x3)))));
  assign n2503 = x2 ? ((~x4 | x5 | x6 | x1 | ~x3) & (x4 | ~x5 | (x1 ? (~x3 ^ ~x6) : (x3 | ~x6)))) : ((~x1 | x5 | ~x6 | (~x3 ^ x4)) & (x1 | x3 | ~x4 | ~x5 | x6));
  assign n2504 = (n406 | n2507) & (~n615 | n2505) & (~x0 | n2506);
  assign n2505 = x0 ? (x1 | ((~x3 | (~x2 ^ ~x6)) & (~x2 | (x6 ? ~x4 : x3)))) : ((~x1 | ((x2 | x6) & (x4 | ~x6 | ~x2 | x3))) & (x2 | ~x6 | (x1 & ~x3)));
  assign n2506 = (x3 | ((x4 | x5 | ~x6 | x1 | ~x2) & (~x1 | ((~x5 | ~x6 | x2 | ~x4) & (x5 | x6 | ~x2 | x4))))) & (x1 | ~x3 | x6 | (x2 ? ~x5 : (x4 | x5)));
  assign n2507 = (x0 | ~x1 | ~x2 | ~x4 | ~x5 | ~x6) & (x2 | ((x0 | x1 | x4 | ~x5 | x6) & (~x0 | ((x5 | x6 | x1 | ~x4) & (~x5 | ~x6 | ~x1 | x4)))));
  assign z196 = n2509 | ~n2511 | n2518 | (~x1 & ~n2519);
  assign n2509 = x2 & ((n1585 & n996) | (x3 & ~n2510));
  assign n2510 = x0 ? (x1 | ((~x6 | ~x7 | ~x4 | ~x5) & (x6 | x7 | x4 | x5))) : (~x1 | x5 | ~x6 | (~x4 ^ ~x7));
  assign n2511 = n2513 & ~n2517 & (n437 | n2512) & (x4 | n2516);
  assign n2512 = (~x2 | (x1 ? (x3 | (x4 & (x0 | x5))) : (~x3 | (~x4 & ~x5)))) & (x1 | x2 | (x3 ? (x4 | x5) : ~x4));
  assign n2513 = ~n2515 & (~n464 | ~n1415) & (~x2 | ~n349 | ~n2514);
  assign n2514 = x4 & (x3 ? (~x6 & ~x7) : (x6 & x7));
  assign n2515 = ~x2 & x3 & (x1 ? (~x6 & (x4 | ~x7)) : (x4 & x6));
  assign n2516 = (~x0 | x1 | x2 | x3 | x6 | x7) & (x0 | ~x2 | ~x3 | (x1 ? (~x6 | ~x7) : (x6 | x7)));
  assign n2517 = n542 & ((n313 & n1048) | (x7 & n373 & ~n1085));
  assign n2518 = ~x3 & ((~x2 & ((~x6 & x7 & ~x1 & ~x4) | (x1 & x6 & (~x4 | x7)))) | (~x1 & x2 & ((~x6 & ~x7) | (~x4 & x6 & x7))));
  assign n2519 = (x2 | ~x3 | x4 | ~x5 | ~x6) & (x6 | ((~x2 | ~x7 | (x3 ? (x4 | x5) : (~x4 | ~x5))) & (x2 | x3 | ~x4 | x5 | x7)));
  assign z197 = (~x2 & (~n2521 | (x6 & ~n2524))) | ~n2525 | (x2 & ~x6 & ~n2524);
  assign n2521 = (~x0 | n2523) & (~n2522 | ((~x4 | x6) & (x1 | x4 | ~x6)));
  assign n2522 = ~x7 & ~x5 & ~x0 & ~x3;
  assign n2523 = (~x5 | ~x6 | x7 | x1 | ~x3 | x4) & (~x4 | ((x6 | x7 | x3 | x5) & (~x1 | ~x6 | ~x7 | (~x3 ^ ~x5))));
  assign n2524 = (x4 | ~x5 | x7 | x0 | ~x3) & (~x4 | ~x7 | ((x0 | ((~x1 | ~x3 | ~x5) & (x3 | x5))) & (x1 | ((x3 | x5) & (~x0 | ~x3 | ~x5)))));
  assign n2525 = ~n2527 & n2528 & ~n2530 & (n1367 | n2526) & n2531;
  assign n2526 = x4 ? (~x2 | (x0 & x1)) : x2;
  assign n2527 = ~x4 & n545 & ((n542 & n664) | (n354 & ~n440));
  assign n2528 = x0 | (n2529 & (~x2 | ~x3 | x4 | n440));
  assign n2529 = (~x1 | x2 | x3 | x4 | x5 | x7) & (x1 | ~x2 | ~x3 | ~x4 | ~x5 | ~x7);
  assign n2530 = ~x2 & ~x3 & ((x4 & x5 & x7) | (~x5 & ~x7 & x0 & ~x4));
  assign n2531 = n2394 & ((x0 & ~n321) | ~n929 | ~n2058);
  assign z198 = ~n2535 | (x0 & ~n2533) | (x5 & ~n406 & ~n2534);
  assign n2533 = (x6 | ((x1 | ~x2 | x3 | x4 | ~x5) & (~x1 | x2 | ~x4 | (x3 ^ x5)))) & (~x1 | x2 | ~x3 | x5 | (x4 & ~x6));
  assign n2534 = (x0 | ((x4 | x6) & (~x1 | ~x4 | ~x6))) & (~x4 | ~x6 | ~x1 | x2) & (x1 | ((x2 | x4 | x6) & (~x0 | ~x4 | ~x6)));
  assign n2535 = ~n2536 & ~n2537 & ~n2538 & ~n2539 & (~n958 | ~n339);
  assign n2536 = x5 & x4 & x3 & ~x0 & ~x1;
  assign n2537 = (~x0 | ~x1) & ((~x5 & x6 & x3 & x4) | (~x3 & (x4 ? (~x5 & ~x6) : (x5 & x6))));
  assign n2538 = ~x4 & ((x0 & x1 & ~x3 & x5) | (x3 & ~x5 & (~x0 | ~x1)));
  assign n2539 = x3 & x4 & x5 & ~x6 & (~x0 ^ ~x1);
  assign z199 = n2541 | ~n2544 | (x5 & ~n2543);
  assign n2541 = x0 & ((~x7 & ~n2542) | (~x3 & n1906 & n1637));
  assign n2542 = (~x4 | ~x5 | x6 | x1 | x2 | ~x3) & (~x1 | ~x2 | x3 | x5 | (~x4 ^ x6));
  assign n2543 = (x0 & ((x2 & ~x6) | (x1 & (x2 | ~x6)))) | (x4 & (~x6 ^ x7)) | (~x4 & (x6 ^ x7)) | (~x0 & ~x1 & x6);
  assign n2544 = (x0 & ((x1 & x2) | (x5 & x6))) | (~x4 & (x5 | ~x6)) | (x6 & (x5 ? x1 : x4)) | (x5 & ~x6 & (~x0 | (~x1 & ~x2)));
  assign z200 = (~x7 & ((n1671 & ~n2547) | (x5 & ~n2546))) | ~n2548 | (~x5 & x7 & ~n2546);
  assign n2546 = x0 ? ((x3 & ((x1 & x2) | (x4 & ~x6))) | (x2 & ~x6) | (x1 & (~x6 | (x2 & x4)))) : (x6 & (~x1 | (~x2 & ~x3 & ~x4)));
  assign n2547 = (~x0 | ~x2 | ~x4 | x5 | x6) & (x0 | x2 | x4 | ~x5 | ~x6);
  assign n2548 = (x0 | x1 | ~x5 | ~x6) & (~x0 | x5 | x6 | (n864 & n1884));
  assign z201 = ~n2551 | n2554 | n2555 | (~x2 & ~n2550);
  assign n2550 = (x1 | x7 | ((x0 | x3 | ~x4 | x6) & (~x0 | ~x3 | (x4 ^ x6)))) & (~x4 | x6 | ~x7 | x0 | ~x1 | x3);
  assign n2551 = ~n2553 & n2552 & (x3 | x4 | n437 | ~n1192);
  assign n2552 = (~x0 & (x6 | x7)) | (x1 & x2) | (x6 & x7) | (~x7 & ((~x1 & ~x2) | (x0 & ~x6)));
  assign n2553 = ~x2 & ~x6 & ((x0 & ~x1 & ~x3 & ~x7) | (~x0 & x3 & (~x1 ^ x7)));
  assign n2554 = ~x0 & (x1 ? (x2 & ~x6) : (x6 & x7));
  assign n2555 = n278 & n288 & ((~x1 & x5 & ~x6 & ~x7) | (x1 & x7 & (~x5 ^ ~x6)));
  assign z202 = ~n2560 | n2559 | ~n2557 | n2558;
  assign n2557 = (~n283 | ~n993) & (x7 | (x2 ? ~n349 : n1544));
  assign n2558 = x1 & ~x3 & ((x4 & ~x7 & ~x0 & ~x2) | (~x4 & x7 & x0 & x2));
  assign n2559 = n748 & n531 & (x3 ? (x7 & n321) : (~x7 & n349));
  assign n2560 = (~x0 | x2 | ((~x1 | ~x7) & (x4 | x7 | x1 | ~x3))) & (x1 | ~x7 | (x0 & ~x2 & (~x3 | ~x4)));
  assign z203 = n2563 | ~n2564 | (~x7 & (n2562 | (n283 & n1388)));
  assign n2562 = x0 & ((n1251 & n1728) | (x4 & n312 & n1252));
  assign n2563 = ~x2 & ((~x0 & ((x4 & x5 & ~x1 & x3) | (~x4 & ~x5 & x1 & ~x3))) | (x0 & ~x1 & x3 & ~x4 & ~x5));
  assign n2564 = ~n2565 & n2566 & (x1 ? (~x0 | (x2 & ~n288)) : (x0 | ~x2));
  assign n2565 = x5 & (x3 ? (n548 & n460) : (n547 & n992));
  assign n2566 = (~x0 | x1 | x2 | x3) & (~x2 | ~x3 | x0 | ~x1);
  assign z204 = n2568 | ~n2569 | ~n2571 | (x1 & ~x6 & ~n2570);
  assign n2568 = n345 & n1070 & ((~x0 & ~x3 & x5 & x7) | (x0 & (x3 ? (x5 & ~x7) : (~x5 & x7))));
  assign n2569 = ~n509 | ((~x1 | ~x5 | (x0 ? (x4 | ~x6) : ~x4)) & (x5 | ~x6 | x0 | ~x4) & (x1 | (x0 ? (x4 | (x5 & x6)) : (~x4 | x5))));
  assign n2570 = x0 ? ((x4 | ~x5 | ~x7 | x2 | ~x3) & (~x4 | x5 | x7 | ~x2 | x3)) : (x2 | ((x5 | ~x7 | ~x3 | ~x4) & (~x5 | x7 | x3 | x4)));
  assign n2571 = (~x1 | ((~x3 | ~x4 | ~x0 | x2) & (~x2 | x3 | x4))) & n2572 & (x1 | ((x2 | x3 | ~x4) & (~x3 | (~x2 & (x0 | x4)))));
  assign n2572 = x3 | ((x2 | x4 | n832) & (~x4 | ((~n451 | ~n992) & (~x2 | n832))));
  assign z205 = n2576 | ~n2579 | (~n858 & ~n2574) | (~x1 & ~n2575);
  assign n2574 = (x2 | ((~x1 | ((~x6 | ~x7 | ~x4 | ~x5) & (x4 | x6 | x7))) & (x4 | ((x5 | (~x6 & ~x7)) & (x6 | (x7 ? x1 : ~x5)))))) & (x1 | ((~x6 | x7 | x4 | ~x5) & (~x2 | (~x4 & (~x5 | ~x6)))));
  assign n2575 = (~x0 | x2 | x3 | ~x4 | ~x5 | ~x6) & (x5 | ((x0 | ~x2 | ~x3 | ~x4 | ~x6) & (x4 | ((x0 | x2 | ~x3 | ~x6) & (~x0 | x3 | (x2 ^ x6))))));
  assign n2576 = ~x5 & ((~x6 & ~n2578) | (n532 & n1215 & ~n2577));
  assign n2577 = x1 ? (~x4 | ~x7) : (x4 | x7);
  assign n2578 = (~x3 | x4 | x7 | ~x0 | x1 | x2) & ((x1 ? (~x4 | x7) : (x4 | ~x7)) | (x0 ? (~x2 | x3) : (x2 | ~x3)));
  assign n2579 = ~n2580 & ~n2581 & n2582 & (~n292 | ~n654 | ~n463);
  assign n2580 = x1 & (x0 ? (~x3 & (x2 ? ~x4 : (x4 & x5))) : (x3 & (~x2 ^ x4)));
  assign n2581 = (x4 ^ x5) & ((x0 & ~x1 & x2 & ~x3) | (~x0 & (x1 ? (x2 & ~x3) : (~x2 & x3))));
  assign n2582 = ~x4 | ~x5 | (x3 ? ~n686 : (x6 | ~n992));
  assign z206 = n2593 | n2592 | ~n2589 | ~n2587 | n2584 | ~n2586;
  assign n2584 = ~x3 & ((n1336 & n786) | (~x7 & ~n2585));
  assign n2585 = (x0 | x1 | x2 | x4 | ~x5 | ~x6) & (~x0 | x5 | ((x4 | x6 | x1 | ~x2) & (~x1 | ~x4 | (~x2 ^ x6))));
  assign n2586 = (n399 | n535) & (n1079 | n1117);
  assign n2587 = ~n2588 & (~n1100 | ~n531 | (x1 ? ~x4 : ~n748));
  assign n2588 = ~n585 & ~n858 & ((n542 & n664) | (n354 & n870));
  assign n2589 = ~n2590 & n2591 & ((~x0 & ~n359) | n1291 | (x0 & ~n452));
  assign n2590 = ~n980 & (x2 ? (n870 & n349) : (n664 & n321));
  assign n2591 = x3 | ~n345 | ((x0 | ~x4 | ~x5) & (x5 | x6 | ~x0 | x4));
  assign n2592 = ~n1085 & (x0 ? (x3 & (x1 ? (~x2 & x4) : ~x4)) : (~x3 & (x1 ^ ~x4)));
  assign n2593 = ~n1971 & ((x0 & ~x1 & ~x3 & ~x4 & x6) | (~x0 & x3 & ~x6 & (x1 ^ ~x4)));
  assign z207 = (~x1 & ~n2595) | (x1 & ~n2596) | n2597 | (x5 & ~n2602);
  assign n2595 = (x2 | (x4 ? (~x6 | (~x7 & (x0 | ~x3))) : ((~x0 | ((x6 | ~x7) & (x3 | ~x6 | x7))) & (x6 | ((x3 | ~x7) & (x0 | ~x3 | x7)))))) & (~x0 | x3 | ~x4 | ~x6 | ~x7) & (~x2 | ((~x4 | x6 | ~x7 | x0 | ~x3) & (x7 | (~x0 & x3) | (x4 ^ x6))));
  assign n2596 = (x2 | ((~x6 | ~x7 | ~x3 | x4) & (~x4 | ((~x0 | ((x6 | ~x7) & (x3 | ~x6 | x7))) & (x6 | (x7 ? x3 : x0)))))) & (x0 | x3 | ~x4 | x6 | x7) & (x4 | ~x6 | ((~x2 | x3 | ~x7) & (x0 | (x7 ? x3 : ~x2))));
  assign n2597 = ~x5 & (n2599 | ~n2600 | (~x0 & ~n2598));
  assign n2598 = (~x1 | x2 | x4 | ~x6 | x7) & (x1 | ~x4 | ((x6 | x7 | ~x2 | x3) & (x2 | (x3 ? (x6 | ~x7) : (~x6 | x7)))));
  assign n2599 = ~n589 & ((~x0 & ~x1 & x2 & ~x3 & x7) | (x0 & ((x3 & x7 & ~x1 & x2) | (x1 & ~x7 & (x2 ^ x3)))));
  assign n2600 = ~n2601 & (n390 | n1117) & (~n292 | ~n313 | ~n459);
  assign n2601 = (~x4 ^ x6) & ((x0 & ~x1 & ~x2 & ~x7) | (~x0 & x1 & x2 & x7));
  assign n2602 = ~n2605 & (n390 | n2566) & (x2 ? n2603 : n2604);
  assign n2603 = (~x4 | x6 | ~x7 | x0 | ~x1 | x3) & (x1 | ((x0 | ~x3 | ~x4 | ~x6 | ~x7) & (~x0 | x3 | x4 | (~x6 ^ x7))));
  assign n2604 = x1 ? ((~x4 | x6 | ~x7 | x0 | ~x3) & (~x0 | x3 | (x4 ? (~x6 | ~x7) : (x6 | x7)))) : (x4 | ((~x6 | x7 | ~x0 | ~x3) & (x0 | (x3 ? (x6 | ~x7) : x7))));
  assign n2605 = ~n585 & ((~x0 & ~x1 & x2 & x3 & ~x7) | ((x1 ? (~x2 & ~x7) : (x2 & x7)) & (x0 ^ ~x3)));
  assign z208 = ~n2609 | (~n505 & ~n2607) | (~n665 & ~n2608);
  assign n2607 = (x0 | ((~x7 | ((x2 | x5 | (x3 ^ x6)) & (~x5 | (~x2 ^ (x3 & ~x6))))) & (x5 | x7 | (x2 ? ~x6 : (~x3 | x6))))) & (x3 | x5 | x7 | ((~x2 | x6) & (~x0 | x2 | ~x6)));
  assign n2608 = x2 ? ((x4 | ~x6 | ~x0 | x3) & (x0 | x1 | ~x3 | x6)) : (x0 ? ((x1 | (x6 ? ~x3 : x4)) & (~x3 | (x4 ^ x6)) & (~x4 | x6 | (~x1 & x3))) : ((x3 | ~x6) & (~x1 | x4 | (x3 & ~x6))));
  assign n2609 = n2610 & ~n2615 & (n440 | n2614) & (~n531 | n2613);
  assign n2610 = x3 ? (n559 | n2612) : n2611;
  assign n2611 = x1 ? ((x4 | x5 | ~x6 | x0 | ~x2) & (~x0 | ((x5 | x6 | ~x2 | x4) & (~x5 | ~x6 | x2 | ~x4)))) : (x0 ? (~x6 | (x2 ? (~x4 | x5) : (x4 | ~x5))) : (~x4 | x6 | (x2 ^ x5)));
  assign n2612 = (~x0 | x1 | ~x4 | x6) & (x0 | (x1 ? (x4 | x6) : (~x4 | ~x6)));
  assign n2613 = (x3 | x4 | ~x7 | x0 | ~x1 | ~x2) & (x2 | ((x0 | x1 | ~x3 | ~x4 | ~x7) & (~x0 | x7 | (x1 ? (~x3 | x4) : (x3 | ~x4)))));
  assign n2614 = x2 ? (x0 ? (x1 | (~x3 ^ (x4 & ~x6))) : ((~x4 | ~x6 | x1 | x3) & (~x1 | x4 | (x3 ^ x6)))) : ((x3 | x4 | ~x6 | ~x0 | ~x1) & (x0 | x1 | ~x3 | ~x4 | x6));
  assign n2615 = ~x6 & (x2 ? ~n2616 : (x5 & ~n2617));
  assign n2616 = x0 ? (x1 | ((~x5 | ~x7 | x3 | x4) & (~x3 | ~x4 | x5 | x7))) : (~x1 | ~x3 | x7 | (x4 ^ x5));
  assign n2617 = (~x0 | ~x1 | x3 | x4 | x7) & (x0 | ~x7 | (x1 ? (~x3 | x4) : (x3 | ~x4)));
  assign z209 = n2619 | n2623 | ~n2627 | (~n437 & ~n2622);
  assign n2619 = ~x3 & (x2 ? ~n2621 : ~n2620);
  assign n2620 = x1 ? ((x0 | x4 | x5 | x6 | x7) & (~x0 | ~x4 | ~x5 | ~x6 | ~x7)) : ((~x4 | x5 | ((~x6 | ~x7) & (~x0 | x6 | x7))) & (~x0 | x4 | ~x5 | (x6 ^ x7)));
  assign n2621 = x0 ? (x1 | ~x4 | (x6 ^ x7)) : (x4 | ((~x5 | x6 | x7) & (~x1 | ((x6 | x7) & (x5 | ~x6 | ~x7)))));
  assign n2622 = x0 ? (x1 ? (x3 | x4 | (~x2 & x5)) : (~x3 | ((~x4 | ~x5) & (x2 | (~x4 & ~x5))))) : ((x3 | ((x2 | (x1 ? (~x4 | ~x5) : x5)) & (x1 | (x5 ? (~x2 & x4) : ~x4)))) & (~x1 | ~x3 | ((x4 | x5) & (~x2 | (x4 & x5)))));
  assign n2623 = x3 & (n2624 | ~n2625 | (~n425 & ~n950 & n837));
  assign n2624 = ~n750 & (x4 ? (n349 & n374) : (n372 & n321));
  assign n2625 = n2626 & (n1513 | ((x0 | ~x2 | x6 | x7) & (~x0 | x2 | ~x6 | ~x7)));
  assign n2626 = (~x4 | ~x6 | ~x7 | x0 | x1 | ~x2) & (x4 | x6 | x7 | ~x0 | ~x1 | x2);
  assign n2627 = ~n2629 & ~n2630 & n2631 & (x0 | n2628);
  assign n2628 = (~x2 | ((x1 | x3 | x4 | x5 | x6) & (~x1 | ~x3 | ~x4 | ~x5 | ~x6))) & (x1 | x2 | ((~x5 | ~x6 | x3 | ~x4) & (~x3 | (x4 ? (~x5 | x6) : (x5 | ~x6)))));
  assign n2629 = ~x2 & n321 & ((n312 & n373) | (~x3 & ~n1707));
  assign n2630 = ~n950 & (x0 ? ((~x3 & x6 & x1 & ~x2) | (x3 & ~x6 & ~x1 & x2)) : (x1 & ~x2 & (~x3 ^ x6)));
  assign n2631 = x0 ? ((x3 | x4 | ~x6 | x1 | ~x2) & (~x3 | ~x4 | x6 | ~x1 | x2)) : (~x2 | ((x4 | ~x6 | x1 | ~x3) & (~x4 | x6 | ~x1 | x3)));
  assign z210 = ~n2635 | n2636 | n2640 | (x0 ? ~n2634 : ~n2633);
  assign n2633 = x1 ? (x2 ? ((x5 | ~x7 | x3 | x4) & (~x5 | x7 | ~x3 | ~x4)) : ((x3 | ~x5 | (x4 ^ x7)) & (x5 | ((~x4 | x7) & (~x3 | x4 | ~x7))))) : ((x2 | ~x3 | ~x7 | (~x4 ^ x5)) & (x7 | ((x4 | x5 | ~x2 | x3) & (x2 | (x3 ? (x4 | x5) : (~x4 | ~x5))))));
  assign n2634 = x7 ? ((x4 | x5 | ~x1 | x2) & (x1 | ((~x2 | ~x3 | ~x4 | ~x5) & (x2 | ((~x4 | x5) & (x3 | x4 | ~x5)))))) : ((x1 | x2 | x4 | x5) & ((x1 ? (x2 | x3) : (~x2 | ~x3)) | (~x4 ^ x5)));
  assign n2635 = x2 ? (x4 ? ((x1 | x3 | ~x7) & (x0 | (x1 ? (x3 | x7) : ~x7))) : ((x1 ^ x7) | (x0 ^ ~x3))) : ((~x0 | ~x1 | ~x3 | ~x4 | x7) & (x0 | x1 | x3 | x4 | ~x7));
  assign n2636 = ~x5 & ((n992 & n2637) | n2639 | (~x1 & ~n2638));
  assign n2637 = ~x7 & ~x6 & x3 & ~x4;
  assign n2638 = (~x4 | x6 | x7 | x0 | ~x2 | ~x3) & (~x7 | ((x0 | x2 | x3 | ~x4 | x6) & (~x0 | ~x6 | (x2 ? (~x3 | ~x4) : (x3 | x4)))));
  assign n2639 = ~n437 & ((~x2 & ~x3 & ~x4 & n349) | (x2 & x3 & (x4 ? n349 : n321)));
  assign n2640 = x5 & (n2641 | n2643 | (~x3 & ~n2642));
  assign n2641 = ~n425 & ((~x0 & ~x1 & x2 & ~x3 & ~x4) | (~x2 & ((x3 & x4 & ~x0 & x1) | (x0 & (x1 ? (~x3 & x4) : (x3 & ~x4))))));
  assign n2642 = (x4 | x6 | ~x7 | x0 | ~x1 | ~x2) & (~x4 | ~x6 | x7 | ~x0 | x1 | x2);
  assign n2643 = n509 & ~n705 & (x0 ? n292 : n543);
  assign z211 = ~n2648 | ~n2651 | (~n307 & ~n2645) | (~x0 & ~n2646);
  assign n2645 = x2 ? ((x1 | ((x5 | ~x6 | x0 | x3) & (~x0 | (x3 ? (x5 | x6) : ~x5)))) & (x0 | ((~x5 | (x3 ^ x6)) & (~x1 | ((~x5 | ~x6) & (~x3 | x5 | x6)))))) : (x3 ? (x5 ? ((~x1 | x6) & (~x0 | (~x1 & x6))) : ((x1 | ~x6) & (x0 | (x1 & ~x6)))) : ((x5 | (~x0 & (~x1 | x6))) & (x0 | x1 | ~x5 | ~x6)));
  assign n2646 = ~n2647 & (~n1252 | ~n786) & (n406 | n585 | n811);
  assign n2647 = n305 & ((x2 & ~n478) | (x4 & n357 & n292));
  assign n2648 = x2 ? (n2650 & (~x1 | x5 | n2649)) : (~x5 | n2649);
  assign n2649 = (~x0 | x3 | ~x4 | x6 | x7) & (x0 | ((~x3 | ~x4 | x6 | x7) & (~x6 | ~x7 | x3 | x4)));
  assign n2650 = x0 ? ((~x4 | x5 | x7 | x1 | ~x3) & (~x5 | ~x7 | x3 | x4)) : (~x5 | (x3 ? (x4 | ~x7) : (~x4 | x7)));
  assign n2651 = (x2 | n2652) & (~x0 | (~n2653 & (x4 | n2654)));
  assign n2652 = (~x0 | ((x4 | x5 | ~x7 | ~x1 | x3) & (~x5 | x7 | ~x3 | ~x4))) & (x5 | ((x0 | x1 | ~x4 | x7) & ((x0 & x1) | (x3 ? (x4 | ~x7) : (~x4 | x7)))));
  assign n2653 = ~n1096 & ((n542 & ~n434) | (n354 & n781));
  assign n2654 = (~x6 | ((x1 | ~x2 | ~x3 | ~x5 | ~x7) & (~x1 | ((x5 | ~x7 | x2 | ~x3) & (~x5 | x7 | ~x2 | x3))))) & (x1 | x6 | ~x7 | (x2 ? (~x3 | x5) : (x3 ^ x5)));
  assign z212 = ~n2657 | ~n2664 | (x1 & ~n2656);
  assign n2656 = (x0 | x3 | x4 | x5 | x6) & (x2 | ((~x4 | ~x5 | x6 | x0 | ~x3) & (~x0 | x4 | x5 | (~x3 ^ x6))));
  assign n2657 = ~n2658 & ~n2659 & n2663 & (~x2 | (~n2661 & ~n2662));
  assign n2658 = ~n390 & ((~x0 & ~x1 & x2 & x3 & x5) | (x1 & ((x0 & ~x3 & (x2 ^ x5)) | (~x0 & ~x2 & x3 & ~x5))));
  assign n2659 = ~n425 & ~n2660;
  assign n2660 = x1 ? (x0 ? (x3 | (x2 ? (x4 | ~x5) : (~x4 | x5))) : (~x3 | x4 | (~x2 ^ x5))) : (~x4 | (x0 ? (x3 | ~x5) : (~x3 | (~x2 ^ x5))));
  assign n2661 = ~n529 & (x4 ? (x7 & n321) : (~x7 & n349));
  assign n2662 = x5 & n1050 & ((n543 & n367) | (~x1 & n292));
  assign n2663 = x3 ? (x0 ? ((~x4 | ~x6 | ~x1 | x2) & (x4 | x6 | x1 | ~x2)) : ((~x1 | ~x2 | ~x4 | x6) & (x4 | ~x6 | x1 | x2))) : ((~x0 | x1 | ~x2 | x4 | ~x6) & (x0 | ((~x1 | ~x4 | ~x6) & (x4 | x6 | x1 | ~x2))));
  assign n2664 = ~n2665 & (n437 | n2668) & (x1 | n2667);
  assign n2665 = ~x2 & ((x4 & ~n2666) | (x0 & n647 & n1197));
  assign n2666 = (~x0 | ((x5 | ~x6 | x7 | x1 | ~x3) & (~x5 | x6 | ~x7 | ~x1 | x3))) & (x5 | ((x0 | x1 | x3 | ~x6 | x7) & (~x7 | ((~x1 | ~x3 | x6) & (x0 | (x1 ? x6 : (~x3 | ~x6)))))));
  assign n2667 = (~x6 | ((~x0 | x2 | x3 | (~x4 ^ x5)) & (~x2 | ((~x4 | ~x5 | ~x0 | ~x3) & (x0 | (x3 ? (x4 | x5) : (~x4 | ~x5))))))) & (x2 | x6 | (~x4 ^ x5) | (~x0 ^ ~x3));
  assign n2668 = (~x5 | ((x3 | x4 | x0 | ~x1) & (x2 | ((x0 | x1 | x3 | ~x4) & (~x0 | ~x3 | (x1 ^ ~x4)))))) & (x1 | x5 | ((x3 | ~x4 | x0 | ~x2) & (~x0 | (x2 ? (~x3 | ~x4) : (x3 | x4)))));
  assign z213 = n2670 | n2674 | n2675 | ~n2677 | (~x3 & ~n2673);
  assign n2670 = ~x7 & ((n1671 & ~n2672) | (~x1 & ~n2671));
  assign n2671 = x3 ? (~x4 | ((~x2 | ~x5 | x6) & (x0 | x2 | x5 | ~x6))) : ((~x0 | ((~x5 | x6 | x2 | x4) & (x5 | ~x6 | ~x2 | ~x4))) & (x0 | x2 | x4 | x5 | ~x6));
  assign n2672 = (~x2 | x5 | ((x4 | ~x6) & (~x0 | ~x4 | x6))) & (~x0 | x2 | ~x5 | (~x4 ^ x6));
  assign n2673 = x4 ? (x5 ? ((x1 | x2 | x7) & (~x0 | (x1 ? (x2 | ~x7) : x7))) : ((~x1 | x2 | x7) & (x0 | ~x2 | (x1 ^ x7)))) : (x1 ? (x2 ? (~x5 | x7) : (x5 | ~x7)) : (~x7 | (x5 ? (~x0 & x2) : ~x2)));
  assign n2674 = ~n307 & ((x0 & ~x1 & ~x2 & ~x3 & ~x5) | (x1 & ((~x2 & x3 & x5) | (~x0 & (x2 ? (x3 & ~x5) : x5)))));
  assign n2675 = ~n2676 & (x2 ? (x5 & ~n585) : (~x5 & ~n589));
  assign n2676 = (~x0 | x1 | ~x3 | ~x7) & (x0 | (x1 ? (~x3 | x7) : (x3 | ~x7)));
  assign n2677 = (~x3 | n2678) & (n1355 | n2679);
  assign n2678 = ((~x4 ^ x7) | ((x1 | (~x2 ^ x5)) & (~x0 | ~x1 | x2 | x5))) & (~x4 | ~x5 | ~x7 | x0 | x1 | ~x2) & (x5 | ((x0 | ~x7 | (x1 ? (x2 | ~x4) : x4)) & (~x0 | x1 | x2 | x4 | x7)));
  assign n2679 = (x5 | (x0 ? ((~x4 | ~x6 | x2 | ~x3) & (x4 | x6 | ~x2 | x3)) : (x2 | (x3 ? (x4 | x6) : (~x4 | ~x6))))) & (x0 | ~x2 | ~x5 | (x3 ? (x4 | ~x6) : (~x4 | x6)));
  assign z214 = n2681 | n2685 | ~n2688 | (x3 ? ~n2684 : ~n2687);
  assign n2681 = ~x0 & (x2 ? ~n2682 : ~n2683);
  assign n2682 = x3 ? ((x5 | ~x6 | x7 | ~x1 | x4) & (x6 | ((~x4 | ~x5 | ~x7) & (x1 | ((~x5 | ~x7) & (~x4 | x5 | x7)))))) : ((~x7 | ((~x5 | ~x6 | x1 | x4) & (~x1 | (x4 ? (~x5 | ~x6) : (x5 | x6))))) & (x5 | ~x6 | x7 | (x1 & ~x4)));
  assign n2683 = (x1 & ~x4 & (~x6 | x7)) | (~x1 & x4 & (x6 | ~x7)) | (~x5 & ~x7) | (x3 & x6) | (~x3 & ~x6) | (x5 & x7);
  assign n2684 = (~x4 | x5 | ~x6 | x0 | ~x1 | x2) & (x1 | ((x0 | ~x2 | x4 | x5 | x6) & (~x0 | ~x5 | (x2 ? (~x4 | ~x6) : (x4 | x6)))));
  assign n2685 = x0 & (~n2686 | (~n852 & ~n1989));
  assign n2686 = (~n268 | ~n996) & (n1591 | (n564 & (~n345 | ~n850)));
  assign n2687 = ((~x4 ^ x6) | ((~x0 | x1 | x2 | ~x5) & (x0 | ~x1 | ~x2 | x5))) & (x4 | x5 | x6 | ~x0 | ~x1 | x2) & (x0 | x1 | ~x5 | (x2 ? (~x4 | ~x6) : (x4 | x6)));
  assign n2688 = n2689 & (~n1100 | ((x1 | x2 | x5 | ~x6) & (~x2 | ((~x5 | ~x6) & (~x1 | x5 | x6)))));
  assign n2689 = ~n2690 & (n1085 | (x0 ? n1884 : (x2 | n2270)));
  assign n2690 = (x1 ? (~x2 & x5) : (x2 & ~x5)) & (x0 ? (x3 ^ x6) : (~x3 & ~x6));
  assign z215 = n2692 | n2696 | ~n2699 | (x7 & ~n2695);
  assign n2692 = x5 & ((n460 & n1693) | n2694 | (~x0 & ~n2693));
  assign n2693 = (~x7 | ((x1 | ~x2 | ~x3 | x4 | x6) & (~x1 | ((~x2 | ~x3 | ~x4 | x6) & (x2 | x3 | x4 | ~x6))))) & (x1 | x7 | ((~x4 | ~x6 | ~x2 | x3) & (x2 | x6 | (x3 ^ x4))));
  assign n2694 = ~n520 & ((~x0 & x1 & x2 & ~x4 & ~x7) | (x0 & ((~x4 & x7 & x1 & ~x2) | (x4 & ~x7 & ~x1 & x2))));
  assign n2695 = (x6 | ((x0 | x1 | x2 | ~x3 | x4) & (x3 | ((x0 | ~x1 | ~x2 | x4) & (~x0 | ~x4 | (x1 ^ ~x2)))))) & (~x2 | ~x6 | ((x0 | (x1 ? (~x3 | x4) : (x3 | ~x4))) & (~x3 | ~x4 | ~x0 | x1)));
  assign n2696 = ~x5 & (n2697 | n2698 | (n543 & n288 & n460));
  assign n2697 = x2 & n349 & ((n292 & n313) | (x3 & ~n1088));
  assign n2698 = ~n699 & (x0 ? ((~x3 & x6 & x1 & ~x2) | (x3 & ~x6 & ~x1 & x2)) : (~x1 & x2 & (~x3 ^ x6)));
  assign n2699 = ~n2700 & ~n2702 & n2703 & n2704 & (n798 | n2701);
  assign n2700 = ~x2 & (((~x3 ^ x6) & (x0 ? (~x1 & x4) : (x1 & ~x4))) | (x0 & x1 & x3 & ~x4 & ~x6) | (~x0 & ~x1 & ~x3 & x4 & x6));
  assign n2701 = (~x0 | x1 | ~x2 | x4 | x7) & (x0 | ~x1 | x2 | ~x4 | ~x7);
  assign n2702 = ~n447 & ((x0 & x1 & ~x2 & ~x7) | (~x0 & ~x1 & x7));
  assign n2703 = (x0 | x1 | ~x3 | ~n1600) & (~x0 | ~x1 | ~x2 | x3 | ~n1070);
  assign n2704 = ~n2705 & (n1427 | ((x1 | x4 | x6 | x7) & (~x1 | ~x4 | ~x6 | ~x7)));
  assign n2705 = (~x3 ^ x6) & ((x4 & ~x7 & ~x0 & x1) | (x0 & ~x1 & ~x4 & x7));
  assign z216 = ~n2707 | n2712 | (x4 & (n2714 | (~x3 & ~n2713)));
  assign n2707 = n2711 & (x4 | n2710) & (x1 ? n2709 : n2708);
  assign n2708 = (~x0 | ((x4 | x5 | ~x7 | x2 | x3) & (~x5 | x7 | ~x2 | ~x4))) & (x0 | ((~x4 | ((~x2 | x5 | ~x7) & (~x5 | x7 | x2 | ~x3))) & (~x2 | x4 | (x5 ^ x7)))) & (~x2 | ((~x4 | (x3 ? (x5 | ~x7) : (~x5 | x7))) & (~x3 | x4 | (x5 ^ x7))));
  assign n2709 = ((x5 ^ x7) | ((~x0 | x2 | x3 | x4) & (x0 | ~x2 | ~x4))) & (~x4 | x5 | ~x7 | ~x0 | x2 | x3) & (x0 | ~x2 | x4 | ((~x5 | x7) & (~x3 | x5 | ~x7)));
  assign n2710 = (~x3 | x6 | x7 | n559 | ~n783) & (x3 | n448 | (x6 ^ ~x7));
  assign n2711 = (x0 & ~x3 & (x4 ? x7 : ~x2)) | (~x0 & (x2 | (x3 & x4 & ~x7))) | (x1 & (x4 ^ x7)) | (x2 & (x3 | x4)) | (~x1 & (~x4 ^ x7));
  assign n2712 = ~n564 & ((~x0 & ~x3 & ~x4 & n374) | (x0 & (x3 ? (~x4 & n374) : ~n555)));
  assign n2713 = (~x0 | ((x1 | x2 | ~x5 | ~x6 | ~x7) & (~x1 | ~x2 | x5 | x6 | x7))) & (x5 | ~x6 | ~x7 | x0 | ~x1 | ~x2);
  assign n2714 = n1100 & ~n559 & (x1 ? (~x6 & ~x7) : (~x6 ^ ~x7));
  assign z217 = n2716 | n2720 | ~n2721 | (~n440 & ~n911) | ~n2723;
  assign n2716 = ~x1 & ((n2717 & n996) | n2719 | (~x4 & ~n2718));
  assign n2717 = x3 & ~x0 & ~x2;
  assign n2718 = (~x5 | x6 | x7 | x0 | x2 | ~x3) & (x5 | ((x0 | x2 | x3 | ~x6 | x7) & (~x7 | ((x0 | x2 | x3 | x6) & (~x0 | ~x2 | (x3 ^ x6))))));
  assign n2719 = ~n539 & ((n664 & n432) | (n870 & n1602));
  assign n2720 = ~x5 & ((x0 & x1 & x2 & ~x3 & ~x4) | (~x2 & ((~x0 & ~x3 & x4) | (x3 & (x0 ^ (x1 & ~x4))))));
  assign n2721 = ~n2722 & (~n588 | ((x1 | (~x0 ^ ~x3)) & (x0 | ((x3 | ~x4) & (~x1 | ~x3 | x4)))));
  assign n2722 = ~n416 & ((~x0 & ~x1 & x2 & x3 & x4) | (x0 & ~x2 & ~x3 & (x1 ^ ~x4)));
  assign n2723 = ~n2724 & ~n2726 & ~n2727 & (x0 | n2725);
  assign n2724 = ~n1085 & ((x0 & ~x1 & x2 & ~x3) | (~x0 & ((~x2 & x3 & x4) | (x1 & x2 & ~x3 & ~x4))));
  assign n2725 = x1 ? ((x2 | x3 | x4 | x5 | x6) & (~x2 | ~x3 | ~x4 | ~x5 | ~x6)) : (~x3 | x4 | ~x6 | (~x2 ^ ~x5));
  assign n2726 = n532 & ((~x1 & ~x3 & x4 & ~x5 & ~x6) | (x1 & ~x4 & (x3 ? (~x5 & ~x6) : (x5 & x6))));
  assign n2727 = x1 & (x0 ? (n929 & n464) : (~n443 & ~n539));
  assign z218 = ~n2730 | n2739 | (x6 ? (x7 ? ~n2738 : ~n2729) : (x7 ? ~n2729 : ~n2738));
  assign n2729 = (~x2 | ((x4 | x5 | ~x0 | x3) & (~x3 | ~x4 | x0 | ~x1))) & (~x1 | ((~x4 | x5 | x0 | ~x3) & (~x0 | x3 | x4))) & (x1 | ((x0 | x2 | x3 | ~x4 | ~x5) & (~x3 | (x0 ? (~x4 | (x2 & ~x5)) : x4)))) & (x0 | x2 | ~x3 | x4 | ~x5);
  assign n2730 = n2731 & ~n2734 & ~n2737 & (x1 ? n2733 : n2736);
  assign n2731 = ~n2732 & (~n509 | ~n783 | ~n611);
  assign n2732 = ~x1 & (x0 ? (~x2 & ~x4 & (x3 ^ x6)) : (x2 & x4 & (~x3 ^ x6)));
  assign n2733 = (x0 | ~x2 | ~x3 | x4 | x6) & (~x0 | x2 | ~x4 | (~x3 ^ x6));
  assign n2734 = ~n559 & ((x0 & ~x1 & x3 & n2735) | (~x0 & x1 & ~x3 & ~n390));
  assign n2735 = ~x7 & x4 & ~x6;
  assign n2736 = (~x4 | x5 | ~x6 | x0 | x2 | ~x3) & ((~x4 ^ x5) | ((~x0 | ~x2 | (~x3 ^ x6)) & (x0 | x2 | x3 | x6)));
  assign n2737 = n349 & ((x2 & ~x3 & ~x4 & ~x5 & x6) | (~x2 & ((x3 & (x4 ? (x5 & x6) : (~x5 & ~x6))) | (x5 & ~x6 & ~x3 & x4))));
  assign n2738 = x0 ? ((x1 | ((x3 | ~x4 | ~x5) & (~x2 | ~x3 | x4 | x5))) & (x2 | (x1 ? (~x3 | x4) : (x3 | ~x4)))) : (x3 | ((x4 | x5 | x1 | ~x2) & (~x1 | (x2 ? (~x4 | x5) : (x4 | ~x5)))));
  assign n2739 = ~x3 & ((n284 & n317) | (~x4 & ~n2740));
  assign n2740 = (x1 | ((x5 | ~x6 | ~x7 | ~x0 | ~x2) & (x0 | ((~x6 | ~x7 | x2 | x5) & (~x2 | ~x5 | x6 | x7))))) & (~x0 | ~x1 | ((x6 | x7 | ~x2 | x5) & (~x6 | ~x7 | x2 | ~x5)));
  assign z219 = n2743 | ~n2747 | ((x4 | (~x7 & ~n2746)) & (~x4 | x7 | ~n2742) & (~x7 | ~n2746));
  assign n2742 = (x3 | ~x5 | ~x6 | x0 | ~x1 | ~x2) & (x1 | ((~x5 | x6 | x0 | x2) & (~x3 | ((~x0 | x6 | (x2 ^ x5)) & (x5 | ~x6 | x0 | ~x2)))));
  assign n2743 = ~x4 & ((n1929 & ~n2745) | (x2 & ~n2744));
  assign n2744 = (~x5 | ((~x0 | x1 | ~x3 | ~x6 | x7) & (x0 | ~x7 | (x1 ? (~x3 | ~x6) : (x3 | x6))))) & (~x0 | x3 | x5 | x6 | (x1 ^ ~x7));
  assign n2745 = (~x0 | ~x1 | x3 | ~x5 | x6) & (x0 | ((~x1 | x5 | ~x6) & (~x5 | x6 | x1 | ~x3)));
  assign n2746 = (x3 | ~x5 | x6 | x0 | ~x1 | ~x2) & (x2 | ((x0 | ~x1 | x3 | x5 | x6) & (~x6 | ((~x0 | (x1 ? (x3 | ~x5) : (~x3 | x5))) & (~x3 | ~x5 | x0 | x1)))));
  assign n2747 = ~n2749 & ~n2750 & n2751 & (x1 | n2748);
  assign n2748 = (~x0 | ~x2 | ~x3 | ~x4 | ~x5 | ~x7) & (x5 | ((x4 | ~x7 | x0 | x3) & ((~x4 ^ x7) | (x0 ? (~x2 | ~x3) : x2))));
  assign n2749 = x5 & n349 & ((~x2 & n369) | (~x3 & n370));
  assign n2750 = ~n307 & (x2 ? (~x3 & ~n832) : ((n783 & n294) | (x3 & ~n832)));
  assign n2751 = ~n2753 & n2754 & (n2752 | (x0 ? (x3 | x5) : (~x3 | ~x5)));
  assign n2752 = (~x1 | x2 | x4 | ~x7) & (x1 | ~x2 | ~x4 | x7);
  assign n2753 = x0 & x1 & ((x4 & ~x7 & ~x2 & x3) | (~x4 & x7 & x2 & ~x3));
  assign n2754 = (((~x0 | x1 | x2 | x3) & (~x2 | ~x3 | x0 | ~x1)) | (x4 ^ x7)) & ((x3 ? (x4 | ~x7) : (~x4 | x7)) | (x0 ? (~x1 | x2) : (x1 | ~x2)));
  assign z220 = n2757 | ~n2758 | ~n2764 | (~x0 & ~n2756);
  assign n2756 = (x5 | ((x1 | x2 | x3 | x6 | ~x7) & (~x1 | ((~x6 | x7 | x2 | ~x3) & (~x2 | ~x7 | (x3 ^ x6)))))) & (~x2 | ~x5 | ((x1 | (x3 ? (x6 | ~x7) : (~x6 | x7))) & (~x6 | x7 | ~x1 | ~x3)));
  assign n2757 = n321 & ((~x2 & x5 & (x3 ? (x6 & ~x7) : (~x6 & x7))) | (~x5 & ((x2 & (x3 ? (~x6 & x7) : (x6 & ~x7))) | (~x6 & ~x7 & ~x2 & x3))));
  assign n2758 = ~n2759 & ~n2760 & n2761 & (~x2 | ~n349 | n529);
  assign n2759 = ~x2 & ((~x0 & ~x5 & (~x1 ^ ~x6)) | (x5 & ((~x0 & ~x1 & x3 & ~x6) | (x0 & (x1 ? (x3 & ~x6) : (~x3 & x6))))));
  assign n2760 = ~n836 & ((~x0 & x1 & ~x3 & x5) | (x0 & (x1 ? (~x3 & ~x5) : (x3 & x5))));
  assign n2761 = ~n2762 & (n2763 | (x0 ? (x1 | x6) : (~x1 | ~x6)));
  assign n2762 = (~x3 ^ x6) & ((~x0 & ~x1 & x2 & x5) | (x0 & (x1 ? (~x2 & x5) : (x2 & ~x5))));
  assign n2763 = (~x2 | ~x3 | x4 | x5 | x7) & (x2 | ((x3 | x4 | ~x5 | x7) & (~x3 | ~x4 | x5 | ~x7)));
  assign n2764 = x6 ? (~n2766 & (~x1 | n2765)) : n2767;
  assign n2765 = (~x4 | ((x0 | ((~x2 | ~x3 | ~x5 | ~x7) & (x2 | x3 | x5 | x7))) & (~x0 | x2 | x3 | ~x5 | x7))) & (~x0 | x4 | (x2 ? (x3 | ~x5) : (x5 | (~x3 ^ ~x7))));
  assign n2766 = ~x3 & x7 & n354 & (x0 ? (x4 ^ x5) : (~x4 ^ x5));
  assign n2767 = (x3 | n2768) & (~x3 | x5 | ~n783 | n936);
  assign n2768 = (~x0 | ~x1 | ~x2 | x4 | ~x5 | ~x7) & (x0 | ~x4 | ((~x1 | ~x2 | ~x5 | ~x7) & (x1 | x2 | x7)));
  assign z221 = n2771 | ~n2773 | ~n2775 | (x4 & (~n2770 | ~n2772));
  assign n2770 = x1 ? ((~x5 | ~x6 | x0 | ~x3) & (x2 | (x3 ? ~x6 : (x5 | x6)))) : ((x2 | ~x3 | x6) & (x5 | ~x6 | ~x2 | x3));
  assign n2771 = ~n425 & ((x1 & x2 & ~x3 & ~x4) | (~x1 & ((x4 & x5 & ~x2 & ~x3) | (x3 & (x2 ? (x4 ^ x5) : (~x4 & ~x5))))));
  assign n2772 = (~x5 | x6 | x7 | x1 | ~x2 | ~x3) & (x3 | x5 | (x2 ^ ~x6) | (x1 ^ ~x7));
  assign n2773 = ~n2774 & ((~x7 & (~x6 | (x4 & x5))) | (~x4 & ~x5) | ~n462 | (x6 & x7));
  assign n2774 = (x2 ? ~n946 : n288) & ((~x0 & x1 & ~x6) | (~x1 & x6));
  assign n2775 = ~n2776 & (n437 | (x1 ? (x2 | n946) : (~x2 | ~n288)));
  assign n2776 = n748 & (x3 ? (x5 & (x1 ^ ~x6)) : (~x6 & n595));
  assign z222 = ~n2778 | n2782 | (x4 & (n2783 | (~x3 & n1626)));
  assign n2778 = ~n2779 & ~n2780 & n2781 & (x7 | ~n279 | n315);
  assign n2779 = x2 & n321 & ((x3 & ~x4 & x5 & ~x7) | (~x3 & (x4 ? (x5 & x7) : (~x5 & ~x7))));
  assign n2780 = ~n1367 & (x2 ? (~x4 & (~x0 | ~x1)) : x4);
  assign n2781 = (x2 | x3 | x4 | ~x7) & (x0 | ~x2 | ~x4 | (x3 ? x7 : (~x5 | ~x7)));
  assign n2782 = ~x4 & ((x5 & x7 & ~x2 & x3) | (~x7 & ((~x2 & x3 & ~x5) | (~x0 & x2 & (~x3 ^ x5)))));
  assign n2783 = x7 & ~n399 & ((x0 & x1 & n1280) | (~n617 & (~x0 | ~x1)));
  assign z223 = n2788 | n2787 | n2786 | n2785 | n2242 | n1926;
  assign n2785 = n1924 & (x3 ? (x4 ? (~x5 & ~x6) : x5) : (x4 & (x5 ^ x6)));
  assign n2786 = ~n1168 & ~n392 & x6 & n654;
  assign n2787 = x4 & (~x0 | ~x1) & (x3 ? (~x5 & ~x6) : (x5 ^ x6));
  assign n2788 = n312 & n686 & n288;
  assign z224 = n2791 | ~n2792 | ~n2794 | (~x4 & ~n2790);
  assign n2790 = (~x5 | x7 | ~n958) & (x6 | (~n958 & (~x3 | x5 | x7 | ~n317)));
  assign n2791 = n1924 & (x6 ? (x5 ? ~n307 : x4) : ~x4);
  assign n2792 = ~n2793 & (~n686 | ~n1197) & (x0 | ~n780 | ~n384);
  assign n2793 = (~x0 ^ ~x1) & (x4 ? (~x5 & x6) : ~x6);
  assign n2794 = (x0 | x1 | ~x4 | x5 | ~x6) & (~x5 | ((x0 | x1 | x4 | x6) & (~x6 | (x0 & x1) | (~x4 ^ ~x7))));
  assign z225 = ~n2796 & (~x0 | ~x1 | ~x2 | (~x3 & ~x4));
  assign n2796 = ~x5 ^ (x6 & ~x7);
  assign z226 = (~n425 & ~n2798) | (n784 & ~n2799);
  assign n2798 = (~x0 & ~x1 & ~x2 & ~x3 & ~x4 & ~x5) | (x0 & x1 & x2 & (x3 | x4));
  assign n2799 = (x0 | x1 | x2 | x4 | ~x6 | ~x7) & (~x0 | ~x1 | ~x2 | ~x4 | x6 | x7);
  assign z227 = ~x7 & (~n2798 | (n784 & ~n2237));
  assign z228 = (~x3 | (~x4 & (~x5 | (~x6 & ~x7)))) & n837 & (x3 | x4 | x5 | x6 | x7);
  assign z229 = ~x0 & (~n2804 | (x3 & x5 & ~n2803));
  assign n2803 = (x1 | x2 | x4 | x6 | ~x7) & (~x1 | ~x2 | ~x4 | ~x6 | x7);
  assign n2804 = (x1 & x2 & x3 & x4 & x5 & x6) | (~x1 & ~x2 & (~x3 | (~x4 & (~x5 | ~x6))));
  assign z230 = n2807 | n2808 | ~n2809 | (n278 & ~n2806);
  assign n2806 = (~x1 | x3 | ~x4 | x5 | x6) & (x1 | ~x3 | x4 | ~x5 | ~x6);
  assign n2807 = ~x1 & (x2 ? (~x0 | ~x3) : (x0 | (x3 & x4)));
  assign n2808 = n1100 & n615 & ((n1906 & n547) | (n345 & n548));
  assign n2809 = x4 | ((x0 | ~x1 | x2 | x3) & (~x0 | x1 | ~x2 | ~x3 | x5));
  assign z231 = ~n2812 | (x5 & (n2811 | (n292 & n373 & n317)));
  assign n2811 = n547 & ((~x0 & x2 & (x1 ? (x3 & x7) : (~x3 & ~x7))) | (x0 & x1 & ~x2 & ~x3 & ~x7));
  assign n2812 = ~n2814 & ~n2815 & ~n2816 & (x2 | n2813) & n2817;
  assign n2813 = (x4 | ~x5 | ~x6 | x0 | x1 | ~x3) & (~x4 | ((~x0 | x6 | (x1 ? (x3 | ~x5) : (~x3 | x5))) & (x3 | x5 | ~x6 | x0 | ~x1)));
  assign n2814 = ~x1 & (x0 ? (~x2 ^ (x3 & x4)) : (x2 ? (~x3 & ~x4) : (x3 & x4)));
  assign n2815 = ~x0 & ~x3 & ((x4 & ~x5 & ~x1 & x2) | (x1 & (x2 ? (~x4 & ~x5) : (x4 & x5))));
  assign n2816 = x0 & ((x3 & ~x4 & x5 & ~x1 & x2) | (~x3 & x4 & ~x5 & x1 & ~x2));
  assign n2817 = (~x0 | ~x1 | x2 | x3 | x4) & (x0 | ((~x1 | x2 | ~x3) & (x3 | ~x4 | ~n451 | x1 | ~x2)));
  assign z232 = ~n2821 | (x5 & ((x6 & ~n2820) | (~n936 & n2819)));
  assign n2819 = ~x6 & x3 & ~x0 & ~x1;
  assign n2820 = (x3 | (x0 ? ((~x4 | ~x7 | ~x1 | x2) & (x4 | x7 | x1 | ~x2)) : (x1 | (x2 ? (~x4 | ~x7) : (x4 | x7))))) & (x0 | ~x1 | ~x3 | (x2 ? (~x4 | ~x7) : (x4 | x7)));
  assign n2821 = ~n2823 & n2824 & ~n2825 & (x2 | n2822) & ~n2826;
  assign n2822 = (x5 | (x0 ? ((~x4 | ~x6 | x1 | ~x3) & (x4 | x6 | ~x1 | x3)) : (x3 | ~x6 | (~x1 ^ ~x4)))) & (x0 | x4 | ~x5 | (x1 ? (~x3 | x6) : (~x3 ^ ~x6)));
  assign n2823 = ~x0 & ((x2 & ((x4 & ~x5 & ~x1 & x3) | (~x4 & x5 & x1 & ~x3))) | (x1 & ~x2 & (x3 ? (~x4 & ~x5) : (x4 & x5))));
  assign n2824 = x1 ? ((x3 | ~x4 | x0 | ~x2) & (~x0 | x2 | ~x3 | x4)) : ((~x0 | (x2 ? (~x3 | ~x4) : (x3 | x4))) & (x4 | ~n269 | x2 | x3) & (x0 | (x2 ? (~x3 | x4) : (~x4 | (~x3 & ~n269)))));
  assign n2825 = x0 & ((x3 & x4 & ~x5 & x1 & ~x2) | (~x1 & (~x3 ^ x5) & (x2 ^ x4)));
  assign n2826 = ~x6 & n1548 & ((x0 & ~x1 & ~x3 & x5) | (~x0 & ~x5 & (~x1 ^ x3)));
  assign z233 = n2828 | ~n2833 | (n2299 & ~n2832) | (x3 & ~n2831);
  assign n2828 = ~x0 & ((x1 & n509 & n1197) | n2830 | (~x1 & ~n2829));
  assign n2829 = (~x2 | x3 | ~x4 | ~x5 | ~x6 | ~x7) & (x2 | ((x3 | x4 | ~x5 | ~x6 | ~x7) & (~x3 | ((x6 | ~x7 | x4 | ~x5) & (~x6 | x7 | ~x4 | x5)))));
  assign n2830 = ~n1277 & ((~x1 & x2 & x4 & ~x6) | (x1 & x6 & (~x2 ^ x4)));
  assign n2831 = (x4 | ~x5 | x6 | ~x0 | x1 | ~x2) & (x5 | (x0 ? (x1 | (x2 ? (~x4 | x6) : (x4 ^ x6))) : ((x1 | x2 | ~x4 | x6) & (~x1 | ~x2 | x4 | ~x6))));
  assign n2832 = (x1 | ~x3 | x5 | x7 | (~x2 ^ ~x4)) & (x3 | ((x1 | ~x2 | x4 | ~x5 | ~x7) & (~x1 | ((~x5 | ~x7 | x2 | ~x4) & (x5 | x7 | ~x2 | x4)))));
  assign n2833 = ~n2835 & n2837 & (x5 ? n2834 : n2836);
  assign n2834 = x0 ? (x2 | ((~x1 | x3 | x4) & (~x4 | (x1 & ~x3)))) : ((~x2 | x3 | x4) & (~x1 | (x2 ? x4 : (x3 | ~x4))));
  assign n2835 = ~n529 & ((x0 & x1 & ~x2 & ~x4) | (~x0 & (x1 ? (~x2 & x4) : (x2 & ~x4))));
  assign n2836 = (x2 | (~x1 ^ ~x3) | (~x0 ^ x4)) & (x1 | ~x2 | (x0 ? (x3 | ~x4) : (~x3 | x4)));
  assign n2837 = ((~x0 ^ ~x2) | (x4 ? (~n273 | ~n451) : n2838)) & (~x0 | x2 | x4 | ~n273 | ~n451) & (x0 | ~x2 | ~x4 | n2838);
  assign n2838 = (~x1 | x3 | x5 | x6) & (~x5 | ~x6 | x1 | ~x3);
  assign z234 = ~n2845 | (~x2 & ~n2840) | (~x0 & (~n2844 | (x2 & ~n2843)));
  assign n2840 = (x5 | n2841) & (x0 | ~x5 | n2842);
  assign n2841 = (x1 | (x0 ? ((x6 | x7 | x3 | ~x4) & (~x6 | ~x7 | ~x3 | x4)) : ((x3 | (x4 ? (~x6 | x7) : (x6 | ~x7))) & (~x6 | ~x7 | ~x3 | ~x4)))) & (x0 | ~x1 | ((~x6 | ~x7 | x3 | x4) & (~x3 | (x4 ? (~x6 | x7) : (x6 | ~x7)))));
  assign n2842 = (x1 | ~x3 | ~x4 | ~x6 | x7) & (x4 | ((x1 | ~x3 | x6 | ~x7) & (~x1 | ~x6 | (~x3 ^ ~x7))));
  assign n2843 = x3 ? ((x5 | ~x6 | x7 | x1 | x4) & (~x5 | ((x6 | ~x7 | x1 | ~x4) & (~x1 | (x4 ? (~x6 | ~x7) : (x6 | x7)))))) : (x6 | ((~x1 | x4 | x5 | x7) & (x1 | (x4 ? (x5 | ~x7) : (~x5 | x7)))));
  assign n2844 = (x4 | (x1 ? ((~x3 | x5 | ~x6) & (x2 | x3 | ~x5 | x6)) : (~x6 | ((x3 | x5) & (x2 | ~x3 | ~x5))))) & (x1 | ((~x4 | ~x5 | x6 | x2 | ~x3) & (~x2 | ~x6 | (x3 ? (~x4 | ~x5) : x5))));
  assign n2845 = ~n2846 & ~n2847 & n2848 & n2849 & (~n460 | ~n848);
  assign n2846 = x1 & ((~x3 & ~x4 & x5 & ~x0 & x2) | (x4 & ((x3 & ~x5 & ~x0 & x2) | (x0 & ~x2 & (~x3 ^ x5)))));
  assign n2847 = x0 & ~x1 & ((x4 & x5 & ~x2 & ~x3) | (x2 & ~x4 & (~x3 ^ x5)));
  assign n2848 = x5 ? ((~x6 | n2836) & (~x2 | x6 | n1011)) : ((x6 | n2836) & (x2 | ~x6 | n1011));
  assign n2849 = (n454 | n661) & (n1011 | n2850);
  assign n2850 = (x2 | ~x5 | x6 | x7) & (~x2 | x5 | ~x6 | ~x7);
  assign z235 = ~n2864 | ~n2861 | ~n2858 | n2856 | n2852 | n2854;
  assign n2852 = ~x0 & ((n268 & n697) | (~x7 & ~n2853));
  assign n2853 = (~x6 | ((~x1 | ~x2 | x3 | ~x4 | ~x5) & (x1 | x2 | (x3 ? (x4 | x5) : (~x4 | ~x5))))) & (~x1 | ~x2 | x6 | (x3 ? (~x4 | x5) : (x4 | ~x5)));
  assign n2854 = ~n425 & ~n2855;
  assign n2855 = x0 ? ((x3 | ((~x2 | x4 | ~x5) & (~x1 | (x2 ? x4 : (~x4 | ~x5))))) & (x4 | x5 | x2 | ~x3) & (x1 | (~x3 & x5) | (x2 ^ x4))) : (x2 ? ((x4 | x5 | x1 | ~x3) & (~x4 | ((x3 | ~x5) & (~x1 | (x3 & ~x5))))) : (x4 ? ((~x3 | x5) & (x1 | (~x3 & x5))) : ((x3 | ~x5) & (~x1 | (x3 & ~x5)))));
  assign n2856 = ~n2857 & ((n288 & n312) | (n531 & n361));
  assign n2857 = (x0 | ~x1 | x2 | ~x7) & (~x0 | x1 | ~x2 | x7);
  assign n2858 = ~n2859 & (n2860 | ((x2 | ~x4 | x5 | x6) & (~x2 | x4 | ~x5 | ~x6)));
  assign n2859 = ~n948 & ((n543 & n349) | (n292 & n321));
  assign n2860 = (~x0 | ~x1 | x3 | x7) & (x0 | x1 | ~x3 | ~x7);
  assign n2861 = n2862 & n2863 & (n1630 | n1591);
  assign n2862 = (~n509 | ~n321 | ~n511) & (~n292 | ~n686 | ~n361);
  assign n2863 = x4 ? ((x6 | ~x7 | n455) & (x7 | n2079 | x3 | ~x6)) : ((~x6 | x7 | n455) & (~x3 | x6 | ~x7 | n2079));
  assign n2864 = (n950 | n2867) & (n1085 | n2865) & (~n748 | n2866);
  assign n2865 = (x3 | ~x4 | x7 | ~x0 | x1 | x2) & ((x1 ? (x2 | ~x4) : (~x2 | x4)) | (x0 ? (~x3 | x7) : (x3 | ~x7)));
  assign n2866 = (x0 | x1 | x6 | ~x7) & (~x0 | x3 | ~x6 | x7);
  assign n2867 = (x0 | ~x2 | ~x3 | (x1 ? (x6 | ~x7) : (~x6 | x7))) & (x3 | x6 | ~x7 | ~x0 | ~x1 | x2);
  assign z236 = n2869 | ~n2872 | (~n699 & ~n2876) | (~n440 & ~n2877);
  assign n2869 = x2 & (x3 ? ~n2871 : (n321 & n2870));
  assign n2870 = ~x4 & (x5 ? (x6 & x7) : (~x6 & ~x7));
  assign n2871 = (x0 | ~x1 | x4 | x5 | x6 | x7) & (x1 | ((x6 | ~x7 | ~x4 | x5) & (~x5 | ~x6 | x7 | ~x0 | x4)));
  assign n2872 = (n1085 | n2875) & (n665 | n2874) & (n2577 | n2873);
  assign n2873 = (~x5 | ~x6 | x2 | x3) & (x0 | ~x2 | (x3 ? (~x5 | ~x6) : (x5 | x6)));
  assign n2874 = x2 ? (x1 ? (x3 | ((x4 | ~x6) & (x0 | (x4 & ~x6)))) : (~x3 | (x4 ^ x6))) : ((~x3 | (x1 ? (~x4 | x6) : (x4 | ~x6))) & (x1 | x3 | (~x4 & x6)));
  assign n2875 = (~x3 | x4 | x7 | ~x1 | x2) & (x1 | ((~x0 | ~x2 | x3 | x4 | x7) & (~x4 | ~x7 | x2 | ~x3)));
  assign n2876 = x1 ? (x2 ? ((x5 | x6 | ~x0 | x3) & (x0 | ~x3 | (~x5 ^ x6))) : (~x6 | (x3 ^ x5))) : (x6 | (x2 ? (x3 | ~x5) : (~x3 | x5)));
  assign n2877 = (x0 | ((x4 | ~x6 | x1 | x3) & (~x1 | ~x2 | ((~x4 | x6) & (~x3 | x4 | ~x6))))) & (x3 | x6 | ~x1 | x2) & (x1 | ((~x4 | ~x6 | ~x2 | x3) & (x2 | (x3 ? (x4 ^ x6) : (x4 | ~x6)))));
  assign z237 = ~n2880 | n2884 | (x2 ? (n321 & ~n2885) : ~n2879);
  assign n2879 = (~x4 | ((~x3 | (x5 ? (x6 | x7) : (~x6 | ~x7))) & (x6 | x7 | x3 | x5))) & (x3 | x4 | ~x5 | ((~x6 | ~x7) & (~x0 | x6 | x7)));
  assign n2880 = ~n2881 & ~n2883 & (n437 | n2882);
  assign n2881 = ~x4 & (x2 ? (~x6 & ((~x0 & x3 & x5) | (~x3 & ~x5))) : (x6 & (~x3 ^ x5)));
  assign n2882 = (x4 | x5 | x2 | ~x3) & (~x2 | ((x3 | x4 | ~x5) & (~x4 | (x0 & x1) | (~x3 & x5))));
  assign n2883 = ~x3 & x4 & x5 & ((~x2 & ~x6) | (~x0 & x2 & x6));
  assign n2884 = n487 & (x3 ? ((x4 & x5 & n374) | (~x5 & (n372 | (~x4 & n374)))) : (x4 ? (~x5 & n374) : (x5 & n372)));
  assign n2885 = (~x6 | ((~x3 | x4 | x5 | ~x7) & (~x4 | ((~x5 | ~x7) & (x3 | (~x5 & ~x7)))))) & (~x3 | x6 | (x5 ? x4 : x7));
  assign z238 = n2887 | n2891 | ~n2892 | (~x4 & ~n2890);
  assign n2887 = ~x6 & ((~x7 & ~n2889) | (n595 & n1929 & ~n2888));
  assign n2888 = x3 ? (x4 ^ x5) : (~x4 | x5);
  assign n2889 = (x4 | ((~x0 | ~x1 | x2 | ~x3 | ~x5) & (x0 | ~x2 | (x1 ? (~x3 | ~x5) : (x3 | x5))))) & (~x0 | ~x1 | x2 | ~x4 | (~x3 ^ x5));
  assign n2890 = (~x1 | x3 | x5 | x6 | x7) & (~x0 | ((~x5 | x6 | x7 | x1 | ~x3) & (x3 | ((x5 | x6 | x7) & (~x5 | ~x6 | ~x7) & (~x1 | (x5 ^ x7))))));
  assign n2891 = n595 & n522 & (x3 ? ((~x5 & x7) | (~x4 & x5 & ~x7)) : (x4 & (x5 | ~x7)));
  assign n2892 = ~n2894 & ((x0 & ~n321) | (n2893 & (n399 | n389)));
  assign n2893 = (~x3 | x4 | x5 | ~x7) & (x3 | ((~x4 | ~x6 | x7) & (x6 | ~x7 | x4 | ~x5)));
  assign n2894 = ~n425 & ((x4 & n321 & ~n1231) | (~x0 & (n2076 | (x4 & ~n1231))));
  assign z239 = n2898 | ~n2899 | (~x7 & (x5 | ~n2896) & (~x5 | ~n2897));
  assign n2896 = (x1 & x2 & (x0 ? x3 : ~x6)) | (x4 & x6) | (~x6 & (~x4 | (x0 & (~x1 | ~x2))));
  assign n2897 = (x0 & ((x1 & x2) | ~x6)) | (~x4 & x6) | (~x6 & (x4 | (x1 & x2 & x3)));
  assign n2898 = (~x0 ^ ~x2) & (x4 ? (~x6 & (x1 | x7)) : (x6 & x7));
  assign n2899 = ~n2900 & (~n288 | ~n374 | ~n524) & (~n321 | ~n2735);
  assign n2900 = x7 & (x4 ^ x6) & (x0 ? (~x1 & x2) : ~x2);
  assign z240 = ~n2902 | (n542 & ((x5 & ~x7 & (x0 ^ ~x6)) | (x0 & ~x5 & (~x6 | x7))));
  assign n2902 = n2903 & n2904 & (x0 | (x1 & ~n870) | (~x1 & n665));
  assign n2903 = x5 | ((~x7 | ~n321) & (x6 | x7 | ~n1906 | n777));
  assign n2904 = (~x7 | ~n2905 | ~x0 | x5) & (x7 | ((~x0 | x1 | (x5 ^ x6)) & (~x5 | ((~x1 | ~x6 | ~n2905) & (x0 | (x6 ? ~x1 : ~n2905))))));
  assign n2905 = ~x4 & ~x3 & x1 & x2;
  assign z241 = ~n2908 | ~n2910 | (~x3 & ~n2907);
  assign n2907 = (x0 | x1 | x2 | ~x4 | x6 | x7) & (~x1 | ~x2 | ((~x6 | x7 | x0 | ~x4) & (x4 | (x0 ? (~x6 ^ x7) : (x6 | x7)))));
  assign n2908 = (x6 | ((x1 | ~x7) & (x0 | (~x7 & (x1 | ~x2))))) & ~n2909 & (~x0 | x1 | ~x6 | x7);
  assign n2909 = n544 & n372 & ((n345 & n850) | (n1906 & n351));
  assign n2910 = (x0 | x2 | ~x3 | x6 | x7) & (~x1 | ((~x3 | ~x6 | x7 | x0 | ~x2) & (x2 | (x0 ? (~x6 ^ x7) : (x6 | x7)))));
  assign z242 = n2913 | ~n2914 | n2915 | (n2522 & ~n2912);
  assign n2912 = (~x1 | ~x2 | ~x4 | x6) & (x1 | x2 | x4 | ~x6);
  assign n2913 = ~x3 & ((~x0 & ((~x1 & ~x2 & x4 & ~x7) | (x1 & x2 & (~x4 ^ x7)))) | (x0 & x1 & x2 & ~x4 & x7));
  assign n2914 = (~x7 & (x0 | (~x1 & ~x2 & (~x5 | ~n288)))) | (x1 & x2) | (~x0 & x7);
  assign n2915 = ~x0 & x3 & (x1 ? (x2 & x7) : (~x2 & ~x7));
  assign z243 = ~n2917 | (x4 & n312 & n929 & ~n891);
  assign n2917 = (x2 & ((~x5 & ~x6 & ~x3 & x4) | (x1 & (x3 | x4)))) | (~x1 & (~x2 | (~x3 & ~x4)));
  assign z244 = ~x2 ^ (~x3 & (~x4 | (~x5 & ~x6 & ~x7)));
  assign z245 = n2921 | ~n2922 | ~n2923 | (n312 & ~n2920);
  assign n2920 = (x3 | ~x4 | x7) & (~x7 | ((x0 | ((~x3 | ~x4) & (x3 | x4 | x1 | x2))) & (~x3 | ~x4 | (x1 & x2))));
  assign n2921 = ~x5 & x6 & ((~x1 & x3 & x4) | (~x0 & ((x3 & x4) | (~x1 & ~x3 & ~x4))));
  assign n2922 = ~n2788 & (x3 | x4 | (~x0 & ~x1 & ~x5));
  assign n2923 = n2924 & (~x4 | ~n509 | ~n595 | (~x5 & ~n450));
  assign n2924 = ~x3 | ~x4 | ~x5 | (x0 & x1);
  assign z246 = ~n2926 & (~x0 | ~x1 | ~x2 | ~x3);
  assign n2926 = (~x4 & ~x5 & ~x6 & ~x7) | (x4 & (x5 | x6 | x7));
  assign z247 = ~n2928 | n2932 | (~x3 & ((n317 & n339) | n2933));
  assign n2928 = ~n2929 & n2931 & (x7 | ~n312 | n2930);
  assign n2929 = (x5 | (~x6 & ~x7)) & (~x0 | ~x1) & (x0 | x1) & (~x5 | x6 | x7);
  assign n2930 = (~x0 | ~x1 | ~x2 | x3) & (x0 | x1 | x2 | ~x3);
  assign n2931 = ~x5 | ((~x0 | ~x1 | x2 | ~x6) & (x0 | x1 | (~x6 & ~x7)));
  assign n2932 = ~x6 & ((~x0 & ~x1 & x2 & ~x5 & ~x7) | (x0 & x1 & ~x2 & (~x5 ^ x7)));
  assign n2933 = x5 & n1548 & n595 & (x6 | x7);
  assign z040 = (~x3 & ~n743) | (~n425 & ~n746) | ~n751 | (x3 & ~n747);
  assign z248 = z226;
  assign z249 = z227;
  assign z251 = z250;
  assign z252 = z250;
  assign z253 = z250;
  assign z254 = z250;
  assign z255 = z250;
  assign z256 = z250;
  assign z257 = z250;
endmodule


