module x_300_mod_47_reg(
    input [300:1] X,
    output [6:1] R
    );


assign R = X % 47;

endmodule
