module x_200_mod_47_reg(
    input [200:1] X,
    output [6:1] R
    );


assign R = X % 47;

endmodule
