module x_200_mod_113(
    input [200:1] X,
    output [7:1] R
    );

wire [7:1] r1,r2,r3,r4,r5,r6,r7,r8,r9,r10,r11,r12,r13,r14,r15,r16,
	r17,r18,r19,r20,r21,r22,r23,r24,r25,r26,r27,r28,r29,r30,r31,r32,r33;   

X_2 label2 (.x0(X[12]),.x1(X[11]),.x2(X[10]),.x3(X[9]),.x4(X[8]),.x5(X[7]),
.z0(r1[7]),.z1(r1[6]),.z2(r1[5]),.z3(r1[4]),.z4(r1[3]),.z5(r1[2]),.z6(r1[1]));

X_3 label3 (.x0(X[18]),.x1(X[17]),.x2(X[16]),.x3(X[15]),.x4(X[14]),.x5(X[13]),
.z0(r2[7]),.z1(r2[6]),.z2(r2[5]),.z3(r2[4]),.z4(r2[3]),.z5(r2[2]),.z6(r2[1]));

X_4 label4 (.x0(X[24]),.x1(X[23]),.x2(X[22]),.x3(X[21]),.x4(X[20]),.x5(X[19]),
.z0(r3[7]),.z1(r3[6]),.z2(r3[5]),.z3(r3[4]),.z4(r3[3]),.z5(r3[2]),.z6(r3[1]));

X_5 label5 (.x0(X[30]),.x1(X[29]),.x2(X[28]),.x3(X[27]),.x4(X[26]),.x5(X[25]),
.z0(r4[7]),.z1(r4[6]),.z2(r4[5]),.z3(r4[4]),.z4(r4[3]),.z5(r4[2]),.z6(r4[1]));

X_6 label6 (.x0(X[36]),.x1(X[35]),.x2(X[34]),.x3(X[33]),.x4(X[32]),.x5(X[31]),
.z0(r5[7]),.z1(r5[6]),.z2(r5[5]),.z3(r5[4]),.z4(r5[3]),.z5(r5[2]),.z6(r5[1]));

X_7 label7 (.x0(X[42]),.x1(X[41]),.x2(X[40]),.x3(X[39]),.x4(X[38]),.x5(X[37]),
.z0(r6[7]),.z1(r6[6]),.z2(r6[5]),.z3(r6[4]),.z4(r6[3]),.z5(r6[2]),.z6(r6[1]));

X_8 label8 (.x0(X[48]),.x1(X[47]),.x2(X[46]),.x3(X[45]),.x4(X[44]),.x5(X[43]),
.z0(r7[7]),.z1(r7[6]),.z2(r7[5]),.z3(r7[4]),.z4(r7[3]),.z5(r7[2]),.z6(r7[1]));

X_9 label9 (.x0(X[54]),.x1(X[53]),.x2(X[52]),.x3(X[51]),.x4(X[50]),.x5(X[49]),
.z0(r8[7]),.z1(r8[6]),.z2(r8[5]),.z3(r8[4]),.z4(r8[3]),.z5(r8[2]),.z6(r8[1]));

X_10 label10 (.x0(X[60]),.x1(X[59]),.x2(X[58]),.x3(X[57]),.x4(X[56]),.x5(X[55]),
.z0(r9[7]),.z1(r9[6]),.z2(r9[5]),.z3(r9[4]),.z4(r9[3]),.z5(r9[2]),.z6(r9[1]));

X_11 label11 (.x0(X[66]),.x1(X[65]),.x2(X[64]),.x3(X[63]),.x4(X[62]),.x5(X[61]),
.z0(r10[7]),.z1(r10[6]),.z2(r10[5]),.z3(r10[4]),.z4(r10[3]),.z5(r10[2]),.z6(r10[1]));

X_12 label12 (.x0(X[72]),.x1(X[71]),.x2(X[70]),.x3(X[69]),.x4(X[68]),.x5(X[67]),
.z0(r11[7]),.z1(r11[6]),.z2(r11[5]),.z3(r11[4]),.z4(r11[3]),.z5(r11[2]),.z6(r11[1]));

X_13 label13 (.x0(X[78]),.x1(X[77]),.x2(X[76]),.x3(X[75]),.x4(X[74]),.x5(X[73]),
.z0(r12[7]),.z1(r12[6]),.z2(r12[5]),.z3(r12[4]),.z4(r12[3]),.z5(r12[2]),.z6(r12[1]));

X_14 label14 (.x0(X[84]),.x1(X[83]),.x2(X[82]),.x3(X[81]),.x4(X[80]),.x5(X[79]),
.z0(r13[7]),.z1(r13[6]),.z2(r13[5]),.z3(r13[4]),.z4(r13[3]),.z5(r13[2]),.z6(r13[1]));

X_15 label15 (.x0(X[90]),.x1(X[89]),.x2(X[88]),.x3(X[87]),.x4(X[86]),.x5(X[85]),
.z0(r14[7]),.z1(r14[6]),.z2(r14[5]),.z3(r14[4]),.z4(r14[3]),.z5(r14[2]),.z6(r14[1]));

X_16 label16 (.x0(X[96]),.x1(X[95]),.x2(X[94]),.x3(X[93]),.x4(X[92]),.x5(X[91]),
.z0(r15[7]),.z1(r15[6]),.z2(r15[5]),.z3(r15[4]),.z4(r15[3]),.z5(r15[2]),.z6(r15[1]));

X_17 label17 (.x0(X[102]),.x1(X[101]),.x2(X[100]),.x3(X[99]),.x4(X[98]),.x5(X[97]),
.z0(r16[7]),.z1(r16[6]),.z2(r16[5]),.z3(r16[4]),.z4(r16[3]),.z5(r16[2]),.z6(r16[1]));

X_18 label18 (.x0(X[108]),.x1(X[107]),.x2(X[106]),.x3(X[105]),.x4(X[104]),.x5(X[103]),
.z0(r17[7]),.z1(r17[6]),.z2(r17[5]),.z3(r17[4]),.z4(r17[3]),.z5(r17[2]),.z6(r17[1]));

X_19 label19 (.x0(X[114]),.x1(X[113]),.x2(X[112]),.x3(X[111]),.x4(X[110]),.x5(X[109]),
.z0(r18[7]),.z1(r18[6]),.z2(r18[5]),.z3(r18[4]),.z4(r18[3]),.z5(r18[2]),.z6(r18[1]));

X_20 label20 (.x0(X[120]),.x1(X[119]),.x2(X[118]),.x3(X[117]),.x4(X[116]),.x5(X[115]),
.z0(r19[7]),.z1(r19[6]),.z2(r19[5]),.z3(r19[4]),.z4(r19[3]),.z5(r19[2]),.z6(r19[1]));

X_21 label21 (.x0(X[126]),.x1(X[125]),.x2(X[124]),.x3(X[123]),.x4(X[122]),.x5(X[121]),
.z0(r20[7]),.z1(r20[6]),.z2(r20[5]),.z3(r20[4]),.z4(r20[3]),.z5(r20[2]),.z6(r20[1]));

X_22 label22 (.x0(X[132]),.x1(X[131]),.x2(X[130]),.x3(X[129]),.x4(X[128]),.x5(X[127]),
.z0(r21[7]),.z1(r21[6]),.z2(r21[5]),.z3(r21[4]),.z4(r21[3]),.z5(r21[2]),.z6(r21[1]));

X_23 label23 (.x0(X[138]),.x1(X[137]),.x2(X[136]),.x3(X[135]),.x4(X[134]),.x5(X[133]),
.z0(r22[7]),.z1(r22[6]),.z2(r22[5]),.z3(r22[4]),.z4(r22[3]),.z5(r22[2]),.z6(r22[1]));

X_24 label24 (.x0(X[144]),.x1(X[143]),.x2(X[142]),.x3(X[141]),.x4(X[140]),.x5(X[139]),
.z0(r23[7]),.z1(r23[6]),.z2(r23[5]),.z3(r23[4]),.z4(r23[3]),.z5(r23[2]),.z6(r23[1]));

X_25 label25 (.x0(X[150]),.x1(X[149]),.x2(X[148]),.x3(X[147]),.x4(X[146]),.x5(X[145]),
.z0(r24[7]),.z1(r24[6]),.z2(r24[5]),.z3(r24[4]),.z4(r24[3]),.z5(r24[2]),.z6(r24[1]));

X_26 label26 (.x0(X[156]),.x1(X[155]),.x2(X[154]),.x3(X[153]),.x4(X[152]),.x5(X[151]),
.z0(r25[7]),.z1(r25[6]),.z2(r25[5]),.z3(r25[4]),.z4(r25[3]),.z5(r25[2]),.z6(r25[1]));

X_27 label27 (.x0(X[162]),.x1(X[161]),.x2(X[160]),.x3(X[159]),.x4(X[158]),.x5(X[157]),
.z0(r26[7]),.z1(r26[6]),.z2(r26[5]),.z3(r26[4]),.z4(r26[3]),.z5(r26[2]),.z6(r26[1]));

X_28 label28 (.x0(X[168]),.x1(X[167]),.x2(X[166]),.x3(X[165]),.x4(X[164]),.x5(X[163]),
.z0(r27[7]),.z1(r27[6]),.z2(r27[5]),.z3(r27[4]),.z4(r27[3]),.z5(r27[2]),.z6(r27[1]));

X_29 label29 (.x0(X[174]),.x1(X[173]),.x2(X[172]),.x3(X[171]),.x4(X[170]),.x5(X[169]),
.z0(r28[7]),.z1(r28[6]),.z2(r28[5]),.z3(r28[4]),.z4(r28[3]),.z5(r28[2]),.z6(r28[1]));

X_30 label30 (.x0(X[180]),.x1(X[179]),.x2(X[178]),.x3(X[177]),.x4(X[176]),.x5(X[175]),
.z0(r29[7]),.z1(r29[6]),.z2(r29[5]),.z3(r29[4]),.z4(r29[3]),.z5(r29[2]),.z6(r29[1]));

X_31 label31 (.x0(X[186]),.x1(X[185]),.x2(X[184]),.x3(X[183]),.x4(X[182]),.x5(X[181]),
.z0(r30[7]),.z1(r30[6]),.z2(r30[5]),.z3(r30[4]),.z4(r30[3]),.z5(r30[2]),.z6(r30[1]));

X_32 label32 (.x0(X[192]),.x1(X[191]),.x2(X[190]),.x3(X[189]),.x4(X[188]),.x5(X[187]),
.z0(r31[7]),.z1(r31[6]),.z2(r31[5]),.z3(r31[4]),.z4(r31[3]),.z5(r31[2]),.z6(r31[1]));

X_33 label33 (.x0(X[198]),.x1(X[197]),.x2(X[196]),.x3(X[195]),.x4(X[194]),.x5(X[193]),
.z0(r32[7]),.z1(r32[6]),.z2(r32[5]),.z3(r32[4]),.z4(r32[3]),.z5(r32[2]),.z6(r32[1]));

X_34 label34 (.x0(X[200]),.x1(X[199]),
.z0(r33[7]),.z1(r33[6]),.z2(r33[5]),.z3(r33[4]),.z4(r33[3]),.z5(r33[2]),.z6(r33[1]));

wire [9:1] R_temp_1,R_temp_2,R_temp_3,R_temp_4,R_temp_5,R_temp_6,R_temp_7,R_temp_8,R_temp_9,R_temp_10,R_temp_11;

assign R_temp_1 = r1 + r2 + r3;
assign R_temp_2 = r4 + r5 + r6;
assign R_temp_3 = r7 + r8 + r9;
assign R_temp_4 = r10 + r11 + r12;
assign R_temp_5 = r13 + r14 + r15;
assign R_temp_6 = r16 + r17 + r18;
assign R_temp_7 = r19 + r20 + r21;
assign R_temp_8 = r22 + r23 + r24;
assign R_temp_9 = r25 + r26 + r27;
assign R_temp_10 = r28 + r29 + r30;
assign R_temp_11 = r31 + r32 + r33;

wire [10:1] R_temp_12,R_temp_13,R_temp_14,R_temp_15;

assign R_temp_12 = R_temp_1 + R_temp_2 + R_temp_3;
assign R_temp_13 = R_temp_4 + R_temp_5 + R_temp_6;
assign R_temp_14 = R_temp_7 + R_temp_8 + R_temp_9;
assign R_temp_15 = R_temp_10 + R_temp_11  + X[6:1];

wire [11:1] R_temp_16,R_temp_17;

assign R_temp_16 = R_temp_12 + R_temp_13;
assign R_temp_17 = R_temp_14 + R_temp_15;

wire [9:1] R_temp_18;

assign R_temp_18 = R_temp_16 [6:1] + 64 * R_temp_16 [7] + 15 * R_temp_16 [11:8] + 
            R_temp_17 [6:1] + 64* R_temp_17 [7] + 15* R_temp_17 [11:8];

wire [8:1] R_temp_19;

assign R_temp_19 = R_temp_18 [6:1] + 64 * R_temp_18 [7] + 15 * R_temp_18 [9:8];


reg [7:1]  R_temp;

always @(R_temp_19)
begin
  if (R_temp_19 >= 7'b1110001  )
    R_temp <= R_temp_19 - 7'b1110001;
  else
    R_temp <= R_temp_19;
end

assign R = R_temp;

endmodule