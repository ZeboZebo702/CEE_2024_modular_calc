module x_100_mod_503(
    input [100:1] X,
    output [9:1] R
    );

wire [9:1] r1,r2,r3,r4,r5,r6,r7,r8,r9,r10,r11,r12,r13,r14,r15,r16;

X_2 label2 (.x0(X[12]),.x1(X[11]),.x2(X[10]),.x3(X[9]),.x4(X[8]),.x5(X[7]),
.z0(r1[9]),.z1(r1[8]),.z2(r1[7]),.z3(r1[6]),.z4(r1[5]),.z5(r1[4]),.z6(r1[3]),.z7(r1[2]),.z8(r1[1]));

X_3 label3 (.x0(X[18]),.x1(X[17]),.x2(X[16]),.x3(X[15]),.x4(X[14]),.x5(X[13]),
.z0(r2[9]),.z1(r2[8]),.z2(r2[7]),.z3(r2[6]),.z4(r2[5]),.z5(r2[4]),.z6(r2[3]),.z7(r2[2]),.z8(r2[1]));

X_4 label4 (.x0(X[24]),.x1(X[23]),.x2(X[22]),.x3(X[21]),.x4(X[20]),.x5(X[19]),
.z0(r3[9]),.z1(r3[8]),.z2(r3[7]),.z3(r3[6]),.z4(r3[5]),.z5(r3[4]),.z6(r3[3]),.z7(r3[2]),.z8(r3[1]));

X_5 label5 (.x0(X[30]),.x1(X[29]),.x2(X[28]),.x3(X[27]),.x4(X[26]),.x5(X[25]),
.z0(r4[9]),.z1(r4[8]),.z2(r4[7]),.z3(r4[6]),.z4(r4[5]),.z5(r4[4]),.z6(r4[3]),.z7(r4[2]),.z8(r4[1]));

X_6 label6 (.x0(X[36]),.x1(X[35]),.x2(X[34]),.x3(X[33]),.x4(X[32]),.x5(X[31]),
.z0(r5[9]),.z1(r5[8]),.z2(r5[7]),.z3(r5[6]),.z4(r5[5]),.z5(r5[4]),.z6(r5[3]),.z7(r5[2]),.z8(r5[1]));

X_7 label7 (.x0(X[42]),.x1(X[41]),.x2(X[40]),.x3(X[39]),.x4(X[38]),.x5(X[37]),
.z0(r6[9]),.z1(r6[8]),.z2(r6[7]),.z3(r6[6]),.z4(r6[5]),.z5(r6[4]),.z6(r6[3]),.z7(r6[2]),.z8(r6[1]));

X_8 label8 (.x0(X[48]),.x1(X[47]),.x2(X[46]),.x3(X[45]),.x4(X[44]),.x5(X[43]),
.z0(r7[9]),.z1(r7[8]),.z2(r7[7]),.z3(r7[6]),.z4(r7[5]),.z5(r7[4]),.z6(r7[3]),.z7(r7[2]),.z8(r7[1]));

X_9 label9 (.x0(X[54]),.x1(X[53]),.x2(X[52]),.x3(X[51]),.x4(X[50]),.x5(X[49]),
.z0(r8[9]),.z1(r8[8]),.z2(r8[7]),.z3(r8[6]),.z4(r8[5]),.z5(r8[4]),.z6(r8[3]),.z7(r8[2]),.z8(r8[1]));

X_10 label10 (.x0(X[60]),.x1(X[59]),.x2(X[58]),.x3(X[57]),.x4(X[56]),.x5(X[55]),
.z0(r9[9]),.z1(r9[8]),.z2(r9[7]),.z3(r9[6]),.z4(r9[5]),.z5(r9[4]),.z6(r9[3]),.z7(r9[2]),.z8(r9[1]));

X_11 label11 (.x0(X[66]),.x1(X[65]),.x2(X[64]),.x3(X[63]),.x4(X[62]),.x5(X[61]),
.z0(r10[9]),.z1(r10[8]),.z2(r10[7]),.z3(r10[6]),.z4(r10[5]),.z5(r10[4]),.z6(r10[3]),.z7(r10[2]),.z8(r10[1]));

X_12 label12 (.x0(X[72]),.x1(X[71]),.x2(X[70]),.x3(X[69]),.x4(X[68]),.x5(X[67]),
.z0(r11[9]),.z1(r11[8]),.z2(r11[7]),.z3(r11[6]),.z4(r11[5]),.z5(r11[4]),.z6(r11[3]),.z7(r11[2]),.z8(r11[1]));

X_13 label13 (.x0(X[78]),.x1(X[77]),.x2(X[76]),.x3(X[75]),.x4(X[74]),.x5(X[73]),
.z0(r12[9]),.z1(r12[8]),.z2(r12[7]),.z3(r12[6]),.z4(r12[5]),.z5(r12[4]),.z6(r12[3]),.z7(r12[2]),.z8(r12[1]));

X_14 label14 (.x0(X[84]),.x1(X[83]),.x2(X[82]),.x3(X[81]),.x4(X[80]),.x5(X[79]),
.z0(r13[9]),.z1(r13[8]),.z2(r13[7]),.z3(r13[6]),.z4(r13[5]),.z5(r13[4]),.z6(r13[3]),.z7(r13[2]),.z8(r13[1]));

X_15 label15 (.x0(X[90]),.x1(X[89]),.x2(X[88]),.x3(X[87]),.x4(X[86]),.x5(X[85]),
.z0(r14[9]),.z1(r14[8]),.z2(r14[7]),.z3(r14[6]),.z4(r14[5]),.z5(r14[4]),.z6(r14[3]),.z7(r14[2]),.z8(r14[1]));

X_16 label16 (.x0(X[96]),.x1(X[95]),.x2(X[94]),.x3(X[93]),.x4(X[92]),.x5(X[91]),
.z0(r15[9]),.z1(r15[8]),.z2(r15[7]),.z3(r15[6]),.z4(r15[5]),.z5(r15[4]),.z6(r15[3]),.z7(r15[2]),.z8(r15[1]));

X_17 label17 (.x0(X[100]),.x1(X[99]),.x2(X[98]),.x3(X[97]),
.z0(r16[9]),.z1(r16[8]),.z2(r16[7]),.z3(r16[6]),.z4(r16[5]),.z5(r16[4]),.z6(r16[3]),.z7(r16[2]),.z8(r16[1]));

wire [11:1] R_temp_1,R_temp_2,R_temp_3,R_temp_4,R_temp_5;

assign R_temp_1 = r1 + r2 + r3;
assign R_temp_2 = r4 + r5 + r6;
assign R_temp_3 = r7 + r8 + r9;
assign R_temp_4 = r10 + r11 + r12;
assign R_temp_5 = r13 + r14 + r15;

wire [12:1] R_temp_6,R_temp_7;

assign R_temp_6 = R_temp_1 + R_temp_2 + R_temp_3;
assign R_temp_7 = R_temp_4 + R_temp_5 + r16;

wire [11:1] R_temp_8;

assign R_temp_8 = R_temp_6 [6:1] + 64 * R_temp_6 [9:7] + 9 * R_temp_6 [12:10] + 
            R_temp_7 [6:1] + 64* R_temp_7 [9:7] + 9 * R_temp_7 [12:10];

wire [10:1] R_temp_9;

assign R_temp_9 = R_temp_8 [6:1] + 64 * R_temp_8 [9:7] + 9 * R_temp_8 [11:10] + X[6:1];


reg [9:1]  R_temp;

always @(R_temp_9)
begin
  if (R_temp_9 >= 9'b111110111  )
    R_temp <= R_temp_9 - 9'b111110111;
  else
    R_temp <= R_temp_9;
end

assign R = R_temp;

endmodule